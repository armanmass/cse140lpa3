-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 20 2019 23:27:50

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23048\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23044\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23021\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22811\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22808\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22511\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22485\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22265\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22262\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22250\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22198\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22188\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21936\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21930\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21912\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21728\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21720\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21639\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21630\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21486\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21401\ : std_logic;
signal \N__21398\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21380\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21299\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21021\ : std_logic;
signal \N__21018\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20916\ : std_logic;
signal \N__20905\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20878\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20861\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20723\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20703\ : std_logic;
signal \N__20702\ : std_logic;
signal \N__20699\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20667\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20660\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20582\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20510\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20468\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20249\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20187\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20118\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20096\ : std_logic;
signal \N__20095\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20089\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20063\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19943\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19835\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19817\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19790\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19782\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19647\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19644\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19620\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19308\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19292\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19062\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18981\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18965\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18644\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18536\ : std_logic;
signal \N__18533\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18521\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18286\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18276\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18248\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17537\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17504\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17312\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17185\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16880\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16692\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16478\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15817\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15405\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15211\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14303\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13841\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13295\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12284\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \latticehx1k_pll_inst.clk\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un44_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un44_ci\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un220_ci\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un4_l_count_11\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.un4_l_count_16_cascade_\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu2.trig_rd_is_det_cascade_\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.un404_ci_cascade_\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.mem0.N_76_i\ : std_logic;
signal \uu2.mem0.N_73_i\ : std_logic;
signal \uu2.mem0.N_79_i\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu0.sec_clkDZ0\ : std_logic;
signal \oneSecStrb_cascade_\ : std_logic;
signal \uu2.N_118_cascade_\ : std_logic;
signal \uu2.N_117\ : std_logic;
signal \uu2.N_117_cascade_\ : std_logic;
signal \INVuu2.w_addr_user_nesr_7C_net\ : std_logic;
signal \uu2.mem0.N_75_i\ : std_logic;
signal \uu2.mem0.N_74_i\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.N_186\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_2_6\ : std_logic;
signal \uu2.N_150_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.N_115_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_0\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.mem0.N_78_i\ : std_logic;
signal \uu2.mem0.N_77_i\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmap_RNIAE522Z0Z_93_cascade_\ : std_logic;
signal \INVuu2.bitmap_215C_net\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.bitmap_RNIKL222Z0Z_212_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \Lab_UT.sec1_3\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmap_pmux_24_i_m2_am_1\ : std_logic;
signal \uu2.un51_w_data_displaying_cascade_\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.w_addr_displaying_4_1\ : std_logic;
signal \uu2.un51_w_data_displaying\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i5_mux_cascade_\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \uu2.bitmap_pmux_29_0_cascade_\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \INVuu2.bitmap_40C_net\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmap_RNI1PH82Z0Z_40_cascade_\ : std_logic;
signal \uu2.N_401_cascade_\ : std_logic;
signal \uu2.N_406\ : std_logic;
signal \uu2.un31_w_data_displaying_1\ : std_logic;
signal \uu2.un49_w_data_displaying_1\ : std_logic;
signal \uu2.mem0.N_81_i\ : std_logic;
signal \uu2.mem0.N_80_i\ : std_logic;
signal \uu2.mem0.N_72_i\ : std_logic;
signal \uu2.N_111_cascade_\ : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.w_data_i_a2_1_0_cascade_\ : std_logic;
signal \uu2.mem0.N_82_i\ : std_logic;
signal \uu2.mem0.N_110\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.N_225\ : std_logic;
signal \uu2.N_144_cascade_\ : std_logic;
signal \uu2.N_361\ : std_logic;
signal \uu2.mem0.w_data_0_a2_0_4_cascade_\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \uu2.N_109\ : std_logic;
signal \uu2.N_111\ : std_logic;
signal \uu2.N_109_cascade_\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \Lab_UT.dispString.N_61\ : std_logic;
signal \Lab_UT.dispString.un46_dOutP_i_m_3\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_3_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_6\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \Lab_UT.dispString.N_50\ : std_logic;
signal \Lab_UT.dispString.N_28_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_3\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.bitmap_pmux_25_bm_1\ : std_logic;
signal \Lab_UT.sec2_3\ : std_logic;
signal \Lab_UT.sec2_2\ : std_logic;
signal \Lab_UT.sec2_1\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \uu2.N_216_cascade_\ : std_logic;
signal \Lab_UT.sec1_1\ : std_logic;
signal \Lab_UT.sec1_2\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.bitmap_pmux_24_i_m2_bm_1_cascade_\ : std_logic;
signal \uu2.bitmap_RNI1UT12Z0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \Lab_UT.min2_2\ : std_logic;
signal \Lab_UT.min2_1\ : std_logic;
signal \Lab_UT.min2_3\ : std_logic;
signal \Lab_UT.min2_0\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.un437_ci_0_cascade_\ : std_logic;
signal \INVuu2.bitmap_69C_net\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \INVuu2.w_addr_displaying_8C_net\ : std_logic;
signal \uu2.un31_w_data_displaying_2\ : std_logic;
signal \uu2.un33_w_data_displaying\ : std_logic;
signal \uu2.w_addr_i_0_tzZ0Z_0\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_3C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_65\ : std_logic;
signal \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \uu2.un15_w_data_displaying_2\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.N_383_cascade_\ : std_logic;
signal \uu2.N_215\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_\ : std_logic;
signal \uu2.bitmap_RNIS4UH1Z0Z_314\ : std_logic;
signal \uu2.N_397\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux_cascade_\ : std_logic;
signal \uu2.bitmap_RNIELSJ2Z0Z_111\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.un21_w_addr_displaying_i\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.N_115\ : std_logic;
signal \uu2.N_144\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_2C_net\ : std_logic;
signal \Lab_UT.dispString.dOutP_1_iv_0_4\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_5\ : std_logic;
signal \Lab_UT.dispString.N_41_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_0Z0Z_0\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \Lab_UT.alarmchar_1\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_0Z0Z_2\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.N_32\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_0Z0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.didp.un2_did_alarmMatch_0_cascade_\ : std_logic;
signal \Lab_UT.sec2_0\ : std_logic;
signal \Lab_UT.loadalarm_0_0_cascade_\ : std_logic;
signal \Lab_UT.sec1_0\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_7\ : std_logic;
signal \uu2.un15_w_data_displaying_5\ : std_logic;
signal \uu2.o_adder_vbuf_w_addr_displaying_6_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_ness_6C_net\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.un15_w_data_displaying_6\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_36\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmap_pmux_25_am_1\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.bitmap_RNIV8902Z0Z_66\ : std_logic;
signal \Lab_UT.min1_2\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmap_pmux_26_bm_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \uu2.N_217\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_11\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_\ : std_logic;
signal \Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_0_sqmuxa_1\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_1_0_i_0\ : std_logic;
signal \Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_127_0_0\ : std_logic;
signal \Lab_UT.trig\ : std_logic;
signal \Lab_UT.dictrl.N_127_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.justentered_0\ : std_logic;
signal \Lab_UT.shifter_ret_3_RNIK5FS8_0\ : std_logic;
signal \Lab_UT.shifter_ret_3_RNIQBH29_0\ : std_logic;
signal \Lab_UT.armed\ : std_logic;
signal \Lab_UT.armed_cascade_\ : std_logic;
signal \Lab_UT.alarmMatch\ : std_logic;
signal \G_203\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8_2_reti\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8_10_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_6\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_7\ : std_logic;
signal bu_rx_data_i_4_fast_3 : std_logic;
signal \buart__rx_shifter_ret_5_fast\ : std_logic;
signal \Lab_UT.dictrl.g1_1Z0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_98_mux_1\ : std_logic;
signal \Lab_UT.dictrl.N_98_mux_0_0\ : std_logic;
signal \Lab_UT.dictrl.g0_3_1_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.un13_qPone\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_2\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_5\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.min1_0\ : std_logic;
signal \Lab_UT.min1_1\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_3\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_1\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_12\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.loadalarm_1\ : std_logic;
signal \Lab_UT.loadalarm_0_0\ : std_logic;
signal \Lab_UT.min1_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.dicRun_2\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.didp.countrce4.un13_qPone\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_0\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMtens_0\ : std_logic;
signal \Lab_UT.dictrl.N_116_mux_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_116_mux_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_1304_0_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1304_0\ : std_logic;
signal \Lab_UT.dictrl.N_1304_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_88_0_0\ : std_logic;
signal \Lab_UT.dictrl.g1_1_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0\ : std_logic;
signal \Lab_UT.dictrl.m25_xZ0Z1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_116_mux_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_4\ : std_logic;
signal \Lab_UT.dictrl.N_98_mux_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_1_1_0\ : std_logic;
signal bu_rx_data_fast_4 : std_logic;
signal \Lab_UT.dictrl.N_98_mux_0\ : std_logic;
signal \Lab_UT.dictrl.g0_3_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_4Z0Z_1\ : std_logic;
signal \buart__rx_shifter_ret_1_fast\ : std_logic;
signal \Lab_UT.dictrl.N_20_0\ : std_logic;
signal \Lab_UT.dictrl.g0_5_2\ : std_logic;
signal bu_rx_data_i_4_fast_7 : std_logic;
signal \buart__rx_sample_g\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_2\ : std_logic;
signal \Lab_UT.didp.di_Sones_1\ : std_logic;
signal \Lab_UT.didp.di_Sones_3\ : std_logic;
signal \Lab_UT.didp.di_Sones_2\ : std_logic;
signal \Lab_UT.didp.di_Mones_1\ : std_logic;
signal \Lab_UT.didp.di_Mones_0\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone\ : std_logic;
signal \Lab_UT.didp.di_Mones_2\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0\ : std_logic;
signal \Lab_UT.didp.di_Mones_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.ce_12_2_3\ : std_logic;
signal \Lab_UT.didp.un24_ce_2\ : std_logic;
signal \Lab_UT.didp.reset_12_1_3\ : std_logic;
signal \Lab_UT.didp.di_Mtens_1\ : std_logic;
signal \Lab_UT.didp.ce_12_3_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Mtens_3\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.un18_ce\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \resetGen.un241_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_count_2_0_4_cascade_\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \Lab_UT.dicRun_1\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.un252_ci\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \Lab_UT.dicLdASones_0\ : std_logic;
signal \Lab_UT.dictrl.g3_1\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_2000_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_2\ : std_logic;
signal \Lab_UT.dicLdAMones_2\ : std_logic;
signal \Lab_UT.dictrl.N_94_0\ : std_logic;
signal \Lab_UT.dictrl.N_2000_0\ : std_logic;
signal \Lab_UT.dictrl.g1\ : std_logic;
signal \Lab_UT.dictrl.g1_3_1\ : std_logic;
signal \Lab_UT.dictrl.N_88_0\ : std_logic;
signal \Lab_UT.dictrl.g1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_0_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_94_0_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_2000_0_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_96_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.m36_0\ : std_logic;
signal \Lab_UT.dictrl.g1_5_0\ : std_logic;
signal \Lab_UT.dictrl.m45_1\ : std_logic;
signal \Lab_UT.dictrl.m25Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_6_0\ : std_logic;
signal \Lab_UT.dictrl.N_5\ : std_logic;
signal \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.state_fast_0\ : std_logic;
signal bu_rx_data_i_4_0 : std_logic;
signal \Lab_UT.dictrl.g1_5\ : std_logic;
signal \Lab_UT.dictrl.g0_5_4\ : std_logic;
signal \Lab_UT.dicLdMones_1\ : std_logic;
signal \Lab_UT.dictrl.N_1300_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_2_0\ : std_logic;
signal \Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_\ : std_logic;
signal \buart__rx_shifter_0_fast_2\ : std_logic;
signal \Lab_UT.dictrl.g0_5_5\ : std_logic;
signal \Lab_UT.dictrl.N_7\ : std_logic;
signal \Lab_UT.dictrl.g0_4_a4_4\ : std_logic;
signal \Lab_UT.dictrl.N_5_2\ : std_logic;
signal \buart__rx_shifter_0_fast_3\ : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal bu_rx_data_4_rep1 : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal bu_rx_data_i_4_7_rep1 : std_logic;
signal \Lab_UT.dictrl.g0_28_1Z0Z_0\ : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal \Lab_UT.dictrl.m31_xZ0Z0\ : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal \Lab_UT.dictrl.g0_43_xZ0\ : std_logic;
signal \Lab_UT.dictrl.N_84_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstate8_2\ : std_logic;
signal \Lab_UT.dictrl.g1_0_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.g0_4_a4Z0Z_5\ : std_logic;
signal \Lab_UT.didp.countrce2.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_0\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.didp.countrce2.un13_qPone\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.di_Stens_1\ : std_logic;
signal \Lab_UT.LdStens\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.LdStens_i_4\ : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal \Lab_UT.didp.di_Sones_0\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.LdSones_i_4\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_1\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.dicLdStens_1\ : std_logic;
signal \Lab_UT.dictrl.N_101_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_fast_3\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep1\ : std_logic;
signal bu_rx_data_rdy_0_g : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.dictrl.g0_9Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.m25Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.N_116_mux_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_120_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1302_0\ : std_logic;
signal \Lab_UT.dictrl.N_119_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0\ : std_logic;
signal \Lab_UT.dictrl.N_120\ : std_logic;
signal \Lab_UT.dictrl.N_99\ : std_logic;
signal \Lab_UT.dictrl.N_96\ : std_logic;
signal \Lab_UT.dictrl.N_99_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_101\ : std_logic;
signal \Lab_UT.dictrl.N_100_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_104_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_99_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_96_0_0\ : std_logic;
signal \Lab_UT.dictrl.g2\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_5\ : std_logic;
signal \Lab_UT.dictrl.N_98_mux_2\ : std_logic;
signal bu_rx_data_i_4_5 : std_logic;
signal \resetGen.escKeyZ0Z_4\ : std_logic;
signal \resetGen.escKeyZ0Z_5_cascade_\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \Lab_UT.dictrl.g1_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_88_2\ : std_logic;
signal bu_rx_data_i_4_3 : std_logic;
signal \Lab_UT.dictrl.N_95_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_103_0\ : std_logic;
signal \Lab_UT.dictrl.g1_2_1_0\ : std_logic;
signal \Lab_UT.dictrl.g1_3\ : std_logic;
signal \Lab_UT.dictrl.N_88\ : std_logic;
signal \Lab_UT.dictrl.N_95\ : std_logic;
signal \Lab_UT.dictrl.N_103\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal \Lab_UT.dictrl.m63_0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_95_0_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_98_mux\ : std_logic;
signal \Lab_UT.dictrl.N_84\ : std_logic;
signal \Lab_UT.dictrl.N_89\ : std_logic;
signal \Lab_UT.dictrl.m68_1\ : std_logic;
signal \Lab_UT.dictrl.N_89_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_99_mux\ : std_logic;
signal \Lab_UT.dictrl.N_102\ : std_logic;
signal \Lab_UT.dictrl.g1_1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g1_2Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_102_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart__rx_ser_clk_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_83\ : std_logic;
signal \Lab_UT.dictrl.N_194_cascade_\ : std_logic;
signal \buart__rx_sample\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal m89_bm : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart__rx_N_27_0_i_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_107_mux_cascade_\ : std_logic;
signal m89_am : std_logic;
signal \buart__rx_hh_0\ : std_logic;
signal \buart__rx_hh_1\ : std_logic;
signal \Lab_UT.dictrl.N_102_mux\ : std_logic;
signal \buart__rx_N_27_0_i\ : std_logic;
signal \buart__rx_startbit_cascade_\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_94_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_2000_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.N_121_mux\ : std_logic;
signal \Lab_UT_dictrl_next_state_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12_RNOZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0_2\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12_RNOZ0Z_4\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12and_a0_1\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12and_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep2\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart__rx_valid_3\ : std_logic;
signal \Lab_UT_dictrl_next_state_3\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.dictrl.N_119_mux\ : std_logic;
signal \Lab_UT.dictrl.i9_mux_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_94\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_2\ : std_logic;
signal \Lab_UT.dictrl.N_90\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_119\ : std_logic;
signal \Lab_UT.dictrl.N_139_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_116_mux\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g2_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_5_1\ : std_logic;
signal \Lab_UT.dictrl.g2_0_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.N_103_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_1302_1_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_119_0_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.g1Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m46_i_0_a5_1\ : std_logic;
signal \Lab_UT.dictrl.N_86\ : std_logic;
signal \Lab_UT.dictrl.N_8\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0\ : std_logic;
signal \Lab_UT_dictrl_un1_next_state66_0\ : std_logic;
signal \Lab_UT.dictrl.m46_i_0_0_0\ : std_logic;
signal bu_rx_data_i_3_1 : std_logic;
signal bu_rx_data_i_4_7 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_i_4_4 : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_1\ : std_logic;
signal \g0_3_4_cascade_\ : std_logic;
signal g0_3_5 : std_logic;
signal \Lab_UT.dictrl.g1Z0Z_2\ : std_logic;
signal \N_12\ : std_logic;
signal \Lab_UT.dictrl.state_0_rep1\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.dictrl.N_13\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_i_4_3_rep1 : std_logic;
signal bu_rx_data_i_4_2 : std_logic;
signal m46_i_0_a3_2 : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_12_3_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart__rx_ser_clk\ : std_logic;
signal \buart__rx_startbit\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_3\ : std_logic;
signal clk_g : std_logic;
signal bu_rx_data_rdy : std_logic;
signal rst_g : std_logic;
signal bu_rx_data_rdy_0 : std_logic;
signal \resetGen.r_m3_i_a3_0_2\ : std_logic;
signal \N_6\ : std_logic;
signal \Lab_UT_dictrl_next_state_0_1_2\ : std_logic;
signal \Lab_UT_dictrl_next_state_0_0_0\ : std_logic;
signal \rst_RNIAL6V33\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__9186\&\N__9489\&\N__9465\&\N__9855\&\N__9942\&\N__9339\&\N__9438\&\N__9405\&\N__9375\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__9300\&\N__9624\&\N__9639\&\N__9309\&\N__9666\&\N__9684\&\N__9549\&\N__10467\&\N__10479\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__11514\&'0'&\N__10341\&'0'&\N__10815\&'0'&\N__10311\&'0'&\N__10452\&'0'&\N__10305\&'0'&\N__10608\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \latticehx1k_pll_inst.clk\,
            REFERENCECLK => \N__8217\,
            RESETB => \N__22914\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22829\,
            RE => \N__22907\,
            WCLKE => \N__10634\,
            WCLK => \N__22828\,
            WE => \N__10635\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23173\,
            DIN => \N__23172\,
            DOUT => \N__23171\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23173\,
            PADOUT => \N__23172\,
            PADIN => \N__23171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23164\,
            DIN => \N__23163\,
            DOUT => \N__23162\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23164\,
            PADOUT => \N__23163\,
            PADIN => \N__23162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23155\,
            DIN => \N__23154\,
            DOUT => \N__23153\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23155\,
            PADOUT => \N__23154\,
            PADIN => \N__23153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23146\,
            DIN => \N__23145\,
            DOUT => \N__23144\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23146\,
            PADOUT => \N__23145\,
            PADIN => \N__23144\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__22807\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23137\,
            DIN => \N__23136\,
            DOUT => \N__23135\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__23137\,
            PADOUT => \N__23136\,
            PADIN => \N__23135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23128\,
            DIN => \N__23127\,
            DOUT => \N__23126\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23128\,
            PADOUT => \N__23127\,
            PADIN => \N__23126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23119\,
            DIN => \N__23118\,
            DOUT => \N__23117\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23119\,
            PADOUT => \N__23118\,
            PADIN => \N__23117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23110\,
            DIN => \N__23109\,
            DOUT => \N__23108\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23110\,
            PADOUT => \N__23109\,
            PADIN => \N__23108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23101\,
            DIN => \N__23100\,
            DOUT => \N__23099\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23101\,
            PADOUT => \N__23100\,
            PADIN => \N__23099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10086\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23092\,
            DIN => \N__23091\,
            DOUT => \N__23090\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23092\,
            PADOUT => \N__23091\,
            PADIN => \N__23090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5648\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23070\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__23070\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__5646\ : InMux
    port map (
            O => \N__23067\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__5645\ : InMux
    port map (
            O => \N__23064\,
            I => \N__23060\
        );

    \I__5644\ : InMux
    port map (
            O => \N__23063\,
            I => \N__23057\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__23060\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__23057\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__5641\ : InMux
    port map (
            O => \N__23052\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__5640\ : InMux
    port map (
            O => \N__23049\,
            I => \N__23044\
        );

    \I__5639\ : InMux
    port map (
            O => \N__23048\,
            I => \N__23039\
        );

    \I__5638\ : InMux
    port map (
            O => \N__23047\,
            I => \N__23039\
        );

    \I__5637\ : LocalMux
    port map (
            O => \N__23044\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__23039\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__5634\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__23028\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__5632\ : InMux
    port map (
            O => \N__23025\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__5631\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23017\
        );

    \I__5630\ : InMux
    port map (
            O => \N__23021\,
            I => \N__23013\
        );

    \I__5629\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23010\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__23007\
        );

    \I__5627\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23004\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__23013\,
            I => \buart__rx_ser_clk\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__23010\,
            I => \buart__rx_ser_clk\
        );

    \I__5624\ : Odrv4
    port map (
            O => \N__23007\,
            I => \buart__rx_ser_clk\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__23004\,
            I => \buart__rx_ser_clk\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__22995\,
            I => \N__22991\
        );

    \I__5621\ : CascadeMux
    port map (
            O => \N__22994\,
            I => \N__22984\
        );

    \I__5620\ : InMux
    port map (
            O => \N__22991\,
            I => \N__22975\
        );

    \I__5619\ : InMux
    port map (
            O => \N__22990\,
            I => \N__22975\
        );

    \I__5618\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22970\
        );

    \I__5617\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22970\
        );

    \I__5616\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22961\
        );

    \I__5615\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22961\
        );

    \I__5614\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22961\
        );

    \I__5613\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22961\
        );

    \I__5612\ : InMux
    port map (
            O => \N__22981\,
            I => \N__22958\
        );

    \I__5611\ : InMux
    port map (
            O => \N__22980\,
            I => \N__22955\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__22975\,
            I => \N__22952\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__22970\,
            I => \N__22949\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__22961\,
            I => \N__22946\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__22958\,
            I => \N__22943\
        );

    \I__5606\ : LocalMux
    port map (
            O => \N__22955\,
            I => \buart__rx_startbit\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__22952\,
            I => \buart__rx_startbit\
        );

    \I__5604\ : Odrv4
    port map (
            O => \N__22949\,
            I => \buart__rx_startbit\
        );

    \I__5603\ : Odrv4
    port map (
            O => \N__22946\,
            I => \buart__rx_startbit\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__22943\,
            I => \buart__rx_startbit\
        );

    \I__5601\ : InMux
    port map (
            O => \N__22932\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__5600\ : CascadeMux
    port map (
            O => \N__22929\,
            I => \N__22925\
        );

    \I__5599\ : InMux
    port map (
            O => \N__22928\,
            I => \N__22922\
        );

    \I__5598\ : InMux
    port map (
            O => \N__22925\,
            I => \N__22919\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__22922\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__22919\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__5595\ : IoInMux
    port map (
            O => \N__22914\,
            I => \N__22911\
        );

    \I__5594\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22908\
        );

    \I__5593\ : IoSpan4Mux
    port map (
            O => \N__22908\,
            I => \N__22904\
        );

    \I__5592\ : SRMux
    port map (
            O => \N__22907\,
            I => \N__22901\
        );

    \I__5591\ : IoSpan4Mux
    port map (
            O => \N__22904\,
            I => \N__22896\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__22901\,
            I => \N__22893\
        );

    \I__5589\ : InMux
    port map (
            O => \N__22900\,
            I => \N__22890\
        );

    \I__5588\ : InMux
    port map (
            O => \N__22899\,
            I => \N__22887\
        );

    \I__5587\ : Span4Mux_s2_h
    port map (
            O => \N__22896\,
            I => \N__22882\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__22893\,
            I => \N__22882\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__22890\,
            I => \N__22877\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22877\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__22882\,
            I => \N__22872\
        );

    \I__5582\ : Span4Mux_s1_h
    port map (
            O => \N__22877\,
            I => \N__22872\
        );

    \I__5581\ : Odrv4
    port map (
            O => \N__22872\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5580\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22866\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__22863\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__5577\ : InMux
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__22857\,
            I => \N__22771\
        );

    \I__5575\ : ClkMux
    port map (
            O => \N__22856\,
            I => \N__22602\
        );

    \I__5574\ : ClkMux
    port map (
            O => \N__22855\,
            I => \N__22602\
        );

    \I__5573\ : ClkMux
    port map (
            O => \N__22854\,
            I => \N__22602\
        );

    \I__5572\ : ClkMux
    port map (
            O => \N__22853\,
            I => \N__22602\
        );

    \I__5571\ : ClkMux
    port map (
            O => \N__22852\,
            I => \N__22602\
        );

    \I__5570\ : ClkMux
    port map (
            O => \N__22851\,
            I => \N__22602\
        );

    \I__5569\ : ClkMux
    port map (
            O => \N__22850\,
            I => \N__22602\
        );

    \I__5568\ : ClkMux
    port map (
            O => \N__22849\,
            I => \N__22602\
        );

    \I__5567\ : ClkMux
    port map (
            O => \N__22848\,
            I => \N__22602\
        );

    \I__5566\ : ClkMux
    port map (
            O => \N__22847\,
            I => \N__22602\
        );

    \I__5565\ : ClkMux
    port map (
            O => \N__22846\,
            I => \N__22602\
        );

    \I__5564\ : ClkMux
    port map (
            O => \N__22845\,
            I => \N__22602\
        );

    \I__5563\ : ClkMux
    port map (
            O => \N__22844\,
            I => \N__22602\
        );

    \I__5562\ : ClkMux
    port map (
            O => \N__22843\,
            I => \N__22602\
        );

    \I__5561\ : ClkMux
    port map (
            O => \N__22842\,
            I => \N__22602\
        );

    \I__5560\ : ClkMux
    port map (
            O => \N__22841\,
            I => \N__22602\
        );

    \I__5559\ : ClkMux
    port map (
            O => \N__22840\,
            I => \N__22602\
        );

    \I__5558\ : ClkMux
    port map (
            O => \N__22839\,
            I => \N__22602\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__22838\,
            I => \N__22602\
        );

    \I__5556\ : ClkMux
    port map (
            O => \N__22837\,
            I => \N__22602\
        );

    \I__5555\ : ClkMux
    port map (
            O => \N__22836\,
            I => \N__22602\
        );

    \I__5554\ : ClkMux
    port map (
            O => \N__22835\,
            I => \N__22602\
        );

    \I__5553\ : ClkMux
    port map (
            O => \N__22834\,
            I => \N__22602\
        );

    \I__5552\ : ClkMux
    port map (
            O => \N__22833\,
            I => \N__22602\
        );

    \I__5551\ : ClkMux
    port map (
            O => \N__22832\,
            I => \N__22602\
        );

    \I__5550\ : ClkMux
    port map (
            O => \N__22831\,
            I => \N__22602\
        );

    \I__5549\ : ClkMux
    port map (
            O => \N__22830\,
            I => \N__22602\
        );

    \I__5548\ : ClkMux
    port map (
            O => \N__22829\,
            I => \N__22602\
        );

    \I__5547\ : ClkMux
    port map (
            O => \N__22828\,
            I => \N__22602\
        );

    \I__5546\ : ClkMux
    port map (
            O => \N__22827\,
            I => \N__22602\
        );

    \I__5545\ : ClkMux
    port map (
            O => \N__22826\,
            I => \N__22602\
        );

    \I__5544\ : ClkMux
    port map (
            O => \N__22825\,
            I => \N__22602\
        );

    \I__5543\ : ClkMux
    port map (
            O => \N__22824\,
            I => \N__22602\
        );

    \I__5542\ : ClkMux
    port map (
            O => \N__22823\,
            I => \N__22602\
        );

    \I__5541\ : ClkMux
    port map (
            O => \N__22822\,
            I => \N__22602\
        );

    \I__5540\ : ClkMux
    port map (
            O => \N__22821\,
            I => \N__22602\
        );

    \I__5539\ : ClkMux
    port map (
            O => \N__22820\,
            I => \N__22602\
        );

    \I__5538\ : ClkMux
    port map (
            O => \N__22819\,
            I => \N__22602\
        );

    \I__5537\ : ClkMux
    port map (
            O => \N__22818\,
            I => \N__22602\
        );

    \I__5536\ : ClkMux
    port map (
            O => \N__22817\,
            I => \N__22602\
        );

    \I__5535\ : ClkMux
    port map (
            O => \N__22816\,
            I => \N__22602\
        );

    \I__5534\ : ClkMux
    port map (
            O => \N__22815\,
            I => \N__22602\
        );

    \I__5533\ : ClkMux
    port map (
            O => \N__22814\,
            I => \N__22602\
        );

    \I__5532\ : ClkMux
    port map (
            O => \N__22813\,
            I => \N__22602\
        );

    \I__5531\ : ClkMux
    port map (
            O => \N__22812\,
            I => \N__22602\
        );

    \I__5530\ : ClkMux
    port map (
            O => \N__22811\,
            I => \N__22602\
        );

    \I__5529\ : ClkMux
    port map (
            O => \N__22810\,
            I => \N__22602\
        );

    \I__5528\ : ClkMux
    port map (
            O => \N__22809\,
            I => \N__22602\
        );

    \I__5527\ : ClkMux
    port map (
            O => \N__22808\,
            I => \N__22602\
        );

    \I__5526\ : ClkMux
    port map (
            O => \N__22807\,
            I => \N__22602\
        );

    \I__5525\ : ClkMux
    port map (
            O => \N__22806\,
            I => \N__22602\
        );

    \I__5524\ : ClkMux
    port map (
            O => \N__22805\,
            I => \N__22602\
        );

    \I__5523\ : ClkMux
    port map (
            O => \N__22804\,
            I => \N__22602\
        );

    \I__5522\ : ClkMux
    port map (
            O => \N__22803\,
            I => \N__22602\
        );

    \I__5521\ : ClkMux
    port map (
            O => \N__22802\,
            I => \N__22602\
        );

    \I__5520\ : ClkMux
    port map (
            O => \N__22801\,
            I => \N__22602\
        );

    \I__5519\ : ClkMux
    port map (
            O => \N__22800\,
            I => \N__22602\
        );

    \I__5518\ : ClkMux
    port map (
            O => \N__22799\,
            I => \N__22602\
        );

    \I__5517\ : ClkMux
    port map (
            O => \N__22798\,
            I => \N__22602\
        );

    \I__5516\ : ClkMux
    port map (
            O => \N__22797\,
            I => \N__22602\
        );

    \I__5515\ : ClkMux
    port map (
            O => \N__22796\,
            I => \N__22602\
        );

    \I__5514\ : ClkMux
    port map (
            O => \N__22795\,
            I => \N__22602\
        );

    \I__5513\ : ClkMux
    port map (
            O => \N__22794\,
            I => \N__22602\
        );

    \I__5512\ : ClkMux
    port map (
            O => \N__22793\,
            I => \N__22602\
        );

    \I__5511\ : ClkMux
    port map (
            O => \N__22792\,
            I => \N__22602\
        );

    \I__5510\ : ClkMux
    port map (
            O => \N__22791\,
            I => \N__22602\
        );

    \I__5509\ : ClkMux
    port map (
            O => \N__22790\,
            I => \N__22602\
        );

    \I__5508\ : ClkMux
    port map (
            O => \N__22789\,
            I => \N__22602\
        );

    \I__5507\ : ClkMux
    port map (
            O => \N__22788\,
            I => \N__22602\
        );

    \I__5506\ : ClkMux
    port map (
            O => \N__22787\,
            I => \N__22602\
        );

    \I__5505\ : ClkMux
    port map (
            O => \N__22786\,
            I => \N__22602\
        );

    \I__5504\ : ClkMux
    port map (
            O => \N__22785\,
            I => \N__22602\
        );

    \I__5503\ : ClkMux
    port map (
            O => \N__22784\,
            I => \N__22602\
        );

    \I__5502\ : ClkMux
    port map (
            O => \N__22783\,
            I => \N__22602\
        );

    \I__5501\ : ClkMux
    port map (
            O => \N__22782\,
            I => \N__22602\
        );

    \I__5500\ : ClkMux
    port map (
            O => \N__22781\,
            I => \N__22602\
        );

    \I__5499\ : ClkMux
    port map (
            O => \N__22780\,
            I => \N__22602\
        );

    \I__5498\ : ClkMux
    port map (
            O => \N__22779\,
            I => \N__22602\
        );

    \I__5497\ : ClkMux
    port map (
            O => \N__22778\,
            I => \N__22602\
        );

    \I__5496\ : ClkMux
    port map (
            O => \N__22777\,
            I => \N__22602\
        );

    \I__5495\ : ClkMux
    port map (
            O => \N__22776\,
            I => \N__22602\
        );

    \I__5494\ : ClkMux
    port map (
            O => \N__22775\,
            I => \N__22602\
        );

    \I__5493\ : ClkMux
    port map (
            O => \N__22774\,
            I => \N__22602\
        );

    \I__5492\ : Glb2LocalMux
    port map (
            O => \N__22771\,
            I => \N__22602\
        );

    \I__5491\ : GlobalMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__5490\ : gio2CtrlBuf
    port map (
            O => \N__22599\,
            I => clk_g
        );

    \I__5489\ : CascadeMux
    port map (
            O => \N__22596\,
            I => \N__22593\
        );

    \I__5488\ : InMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__5486\ : Span4Mux_v
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__5485\ : Span4Mux_h
    port map (
            O => \N__22584\,
            I => \N__22577\
        );

    \I__5484\ : InMux
    port map (
            O => \N__22583\,
            I => \N__22574\
        );

    \I__5483\ : InMux
    port map (
            O => \N__22582\,
            I => \N__22567\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22581\,
            I => \N__22567\
        );

    \I__5481\ : InMux
    port map (
            O => \N__22580\,
            I => \N__22567\
        );

    \I__5480\ : Odrv4
    port map (
            O => \N__22577\,
            I => bu_rx_data_rdy
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__22574\,
            I => bu_rx_data_rdy
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__22567\,
            I => bu_rx_data_rdy
        );

    \I__5477\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22551\
        );

    \I__5476\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22548\
        );

    \I__5475\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22545\
        );

    \I__5474\ : InMux
    port map (
            O => \N__22557\,
            I => \N__22542\
        );

    \I__5473\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22539\
        );

    \I__5472\ : SRMux
    port map (
            O => \N__22555\,
            I => \N__22534\
        );

    \I__5471\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22534\
        );

    \I__5470\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22492\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__22548\,
            I => \N__22489\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__22545\,
            I => \N__22486\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__22542\,
            I => \N__22469\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__22539\,
            I => \N__22466\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22463\
        );

    \I__5464\ : SRMux
    port map (
            O => \N__22533\,
            I => \N__22344\
        );

    \I__5463\ : SRMux
    port map (
            O => \N__22532\,
            I => \N__22344\
        );

    \I__5462\ : SRMux
    port map (
            O => \N__22531\,
            I => \N__22344\
        );

    \I__5461\ : SRMux
    port map (
            O => \N__22530\,
            I => \N__22344\
        );

    \I__5460\ : SRMux
    port map (
            O => \N__22529\,
            I => \N__22344\
        );

    \I__5459\ : SRMux
    port map (
            O => \N__22528\,
            I => \N__22344\
        );

    \I__5458\ : SRMux
    port map (
            O => \N__22527\,
            I => \N__22344\
        );

    \I__5457\ : SRMux
    port map (
            O => \N__22526\,
            I => \N__22344\
        );

    \I__5456\ : SRMux
    port map (
            O => \N__22525\,
            I => \N__22344\
        );

    \I__5455\ : SRMux
    port map (
            O => \N__22524\,
            I => \N__22344\
        );

    \I__5454\ : SRMux
    port map (
            O => \N__22523\,
            I => \N__22344\
        );

    \I__5453\ : SRMux
    port map (
            O => \N__22522\,
            I => \N__22344\
        );

    \I__5452\ : SRMux
    port map (
            O => \N__22521\,
            I => \N__22344\
        );

    \I__5451\ : SRMux
    port map (
            O => \N__22520\,
            I => \N__22344\
        );

    \I__5450\ : SRMux
    port map (
            O => \N__22519\,
            I => \N__22344\
        );

    \I__5449\ : SRMux
    port map (
            O => \N__22518\,
            I => \N__22344\
        );

    \I__5448\ : SRMux
    port map (
            O => \N__22517\,
            I => \N__22344\
        );

    \I__5447\ : SRMux
    port map (
            O => \N__22516\,
            I => \N__22344\
        );

    \I__5446\ : SRMux
    port map (
            O => \N__22515\,
            I => \N__22344\
        );

    \I__5445\ : SRMux
    port map (
            O => \N__22514\,
            I => \N__22344\
        );

    \I__5444\ : SRMux
    port map (
            O => \N__22513\,
            I => \N__22344\
        );

    \I__5443\ : SRMux
    port map (
            O => \N__22512\,
            I => \N__22344\
        );

    \I__5442\ : SRMux
    port map (
            O => \N__22511\,
            I => \N__22344\
        );

    \I__5441\ : SRMux
    port map (
            O => \N__22510\,
            I => \N__22344\
        );

    \I__5440\ : SRMux
    port map (
            O => \N__22509\,
            I => \N__22344\
        );

    \I__5439\ : SRMux
    port map (
            O => \N__22508\,
            I => \N__22344\
        );

    \I__5438\ : SRMux
    port map (
            O => \N__22507\,
            I => \N__22344\
        );

    \I__5437\ : SRMux
    port map (
            O => \N__22506\,
            I => \N__22344\
        );

    \I__5436\ : SRMux
    port map (
            O => \N__22505\,
            I => \N__22344\
        );

    \I__5435\ : SRMux
    port map (
            O => \N__22504\,
            I => \N__22344\
        );

    \I__5434\ : SRMux
    port map (
            O => \N__22503\,
            I => \N__22344\
        );

    \I__5433\ : SRMux
    port map (
            O => \N__22502\,
            I => \N__22344\
        );

    \I__5432\ : SRMux
    port map (
            O => \N__22501\,
            I => \N__22344\
        );

    \I__5431\ : SRMux
    port map (
            O => \N__22500\,
            I => \N__22344\
        );

    \I__5430\ : SRMux
    port map (
            O => \N__22499\,
            I => \N__22344\
        );

    \I__5429\ : SRMux
    port map (
            O => \N__22498\,
            I => \N__22344\
        );

    \I__5428\ : SRMux
    port map (
            O => \N__22497\,
            I => \N__22344\
        );

    \I__5427\ : SRMux
    port map (
            O => \N__22496\,
            I => \N__22344\
        );

    \I__5426\ : SRMux
    port map (
            O => \N__22495\,
            I => \N__22344\
        );

    \I__5425\ : Glb2LocalMux
    port map (
            O => \N__22492\,
            I => \N__22344\
        );

    \I__5424\ : Glb2LocalMux
    port map (
            O => \N__22489\,
            I => \N__22344\
        );

    \I__5423\ : Glb2LocalMux
    port map (
            O => \N__22486\,
            I => \N__22344\
        );

    \I__5422\ : SRMux
    port map (
            O => \N__22485\,
            I => \N__22344\
        );

    \I__5421\ : SRMux
    port map (
            O => \N__22484\,
            I => \N__22344\
        );

    \I__5420\ : SRMux
    port map (
            O => \N__22483\,
            I => \N__22344\
        );

    \I__5419\ : SRMux
    port map (
            O => \N__22482\,
            I => \N__22344\
        );

    \I__5418\ : SRMux
    port map (
            O => \N__22481\,
            I => \N__22344\
        );

    \I__5417\ : SRMux
    port map (
            O => \N__22480\,
            I => \N__22344\
        );

    \I__5416\ : SRMux
    port map (
            O => \N__22479\,
            I => \N__22344\
        );

    \I__5415\ : SRMux
    port map (
            O => \N__22478\,
            I => \N__22344\
        );

    \I__5414\ : SRMux
    port map (
            O => \N__22477\,
            I => \N__22344\
        );

    \I__5413\ : SRMux
    port map (
            O => \N__22476\,
            I => \N__22344\
        );

    \I__5412\ : SRMux
    port map (
            O => \N__22475\,
            I => \N__22344\
        );

    \I__5411\ : SRMux
    port map (
            O => \N__22474\,
            I => \N__22344\
        );

    \I__5410\ : SRMux
    port map (
            O => \N__22473\,
            I => \N__22344\
        );

    \I__5409\ : SRMux
    port map (
            O => \N__22472\,
            I => \N__22344\
        );

    \I__5408\ : Glb2LocalMux
    port map (
            O => \N__22469\,
            I => \N__22344\
        );

    \I__5407\ : Glb2LocalMux
    port map (
            O => \N__22466\,
            I => \N__22344\
        );

    \I__5406\ : Glb2LocalMux
    port map (
            O => \N__22463\,
            I => \N__22344\
        );

    \I__5405\ : GlobalMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__5404\ : gio2CtrlBuf
    port map (
            O => \N__22341\,
            I => rst_g
        );

    \I__5403\ : IoInMux
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__22335\,
            I => bu_rx_data_rdy_0
        );

    \I__5401\ : InMux
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22329\,
            I => \resetGen.r_m3_i_a3_0_2\
        );

    \I__5399\ : InMux
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N_6\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22317\
        );

    \I__5396\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22314\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__22314\,
            I => \N__22311\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__22311\,
            I => \N__22308\
        );

    \I__5393\ : Odrv4
    port map (
            O => \N__22308\,
            I => \Lab_UT_dictrl_next_state_0_1_2\
        );

    \I__5392\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22302\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__22302\,
            I => \Lab_UT_dictrl_next_state_0_0_0\
        );

    \I__5390\ : CEMux
    port map (
            O => \N__22299\,
            I => \N__22296\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22292\
        );

    \I__5388\ : CEMux
    port map (
            O => \N__22295\,
            I => \N__22289\
        );

    \I__5387\ : Span4Mux_s0_h
    port map (
            O => \N__22292\,
            I => \N__22286\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__22289\,
            I => \N__22283\
        );

    \I__5385\ : Span4Mux_v
    port map (
            O => \N__22286\,
            I => \N__22277\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__22283\,
            I => \N__22277\
        );

    \I__5383\ : CEMux
    port map (
            O => \N__22282\,
            I => \N__22274\
        );

    \I__5382\ : Odrv4
    port map (
            O => \N__22277\,
            I => \rst_RNIAL6V33\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__22274\,
            I => \rst_RNIAL6V33\
        );

    \I__5380\ : CascadeMux
    port map (
            O => \N__22269\,
            I => \N__22265\
        );

    \I__5379\ : CascadeMux
    port map (
            O => \N__22268\,
            I => \N__22259\
        );

    \I__5378\ : InMux
    port map (
            O => \N__22265\,
            I => \N__22256\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__22264\,
            I => \N__22253\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__22263\,
            I => \N__22244\
        );

    \I__5375\ : InMux
    port map (
            O => \N__22262\,
            I => \N__22237\
        );

    \I__5374\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22237\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__22256\,
            I => \N__22234\
        );

    \I__5372\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22227\
        );

    \I__5371\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22227\
        );

    \I__5370\ : InMux
    port map (
            O => \N__22251\,
            I => \N__22227\
        );

    \I__5369\ : InMux
    port map (
            O => \N__22250\,
            I => \N__22224\
        );

    \I__5368\ : CascadeMux
    port map (
            O => \N__22249\,
            I => \N__22221\
        );

    \I__5367\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22209\
        );

    \I__5366\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22209\
        );

    \I__5365\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22209\
        );

    \I__5364\ : InMux
    port map (
            O => \N__22243\,
            I => \N__22206\
        );

    \I__5363\ : InMux
    port map (
            O => \N__22242\,
            I => \N__22203\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22193\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__22234\,
            I => \N__22193\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22227\,
            I => \N__22188\
        );

    \I__5359\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22188\
        );

    \I__5358\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22185\
        );

    \I__5357\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22182\
        );

    \I__5356\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22173\
        );

    \I__5355\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22173\
        );

    \I__5354\ : InMux
    port map (
            O => \N__22217\,
            I => \N__22173\
        );

    \I__5353\ : InMux
    port map (
            O => \N__22216\,
            I => \N__22173\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__22209\,
            I => \N__22168\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__22206\,
            I => \N__22168\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22165\
        );

    \I__5349\ : InMux
    port map (
            O => \N__22202\,
            I => \N__22162\
        );

    \I__5348\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22159\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22154\
        );

    \I__5346\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22154\
        );

    \I__5345\ : InMux
    port map (
            O => \N__22198\,
            I => \N__22151\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__22193\,
            I => \N__22146\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__22188\,
            I => \N__22146\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22185\,
            I => \N__22137\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__22182\,
            I => \N__22137\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__22173\,
            I => \N__22137\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__22168\,
            I => \N__22137\
        );

    \I__5338\ : Span4Mux_h
    port map (
            O => \N__22165\,
            I => \N__22134\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__22162\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__22159\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22154\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__22151\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5333\ : Odrv4
    port map (
            O => \N__22146\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5332\ : Odrv4
    port map (
            O => \N__22137\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5331\ : Odrv4
    port map (
            O => \N__22134\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__22119\,
            I => \N__22116\
        );

    \I__5329\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22113\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22113\,
            I => \N__22110\
        );

    \I__5327\ : Odrv12
    port map (
            O => \N__22110\,
            I => \Lab_UT.dictrl.m46_i_0_a5_1\
        );

    \I__5326\ : InMux
    port map (
            O => \N__22107\,
            I => \N__22098\
        );

    \I__5325\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22098\
        );

    \I__5324\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22085\
        );

    \I__5323\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22082\
        );

    \I__5322\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22079\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__22098\,
            I => \N__22076\
        );

    \I__5320\ : InMux
    port map (
            O => \N__22097\,
            I => \N__22073\
        );

    \I__5319\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22068\
        );

    \I__5318\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22068\
        );

    \I__5317\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22065\
        );

    \I__5316\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22062\
        );

    \I__5315\ : InMux
    port map (
            O => \N__22092\,
            I => \N__22057\
        );

    \I__5314\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22057\
        );

    \I__5313\ : InMux
    port map (
            O => \N__22090\,
            I => \N__22049\
        );

    \I__5312\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22049\
        );

    \I__5311\ : InMux
    port map (
            O => \N__22088\,
            I => \N__22049\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__22044\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22044\
        );

    \I__5308\ : LocalMux
    port map (
            O => \N__22079\,
            I => \N__22041\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__22076\,
            I => \N__22033\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__22073\,
            I => \N__22033\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__22068\,
            I => \N__22024\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__22065\,
            I => \N__22024\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22024\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__22024\
        );

    \I__5301\ : InMux
    port map (
            O => \N__22056\,
            I => \N__22021\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__22049\,
            I => \N__22017\
        );

    \I__5299\ : Span4Mux_v
    port map (
            O => \N__22044\,
            I => \N__22012\
        );

    \I__5298\ : Span4Mux_s3_h
    port map (
            O => \N__22041\,
            I => \N__22012\
        );

    \I__5297\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22009\
        );

    \I__5296\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22004\
        );

    \I__5295\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22004\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__22033\,
            I => \N__21997\
        );

    \I__5293\ : Span4Mux_v
    port map (
            O => \N__22024\,
            I => \N__21997\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__21997\
        );

    \I__5291\ : InMux
    port map (
            O => \N__22020\,
            I => \N__21994\
        );

    \I__5290\ : Odrv4
    port map (
            O => \N__22017\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5289\ : Odrv4
    port map (
            O => \N__22012\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22009\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__22004\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5286\ : Odrv4
    port map (
            O => \N__21997\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__21994\,
            I => \Lab_UT.dictrl.N_86\
        );

    \I__5284\ : InMux
    port map (
            O => \N__21981\,
            I => \N__21978\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__21978\,
            I => \Lab_UT.dictrl.N_8\
        );

    \I__5282\ : CascadeMux
    port map (
            O => \N__21975\,
            I => \N__21972\
        );

    \I__5281\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21969\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__21969\,
            I => \N__21965\
        );

    \I__5279\ : InMux
    port map (
            O => \N__21968\,
            I => \N__21962\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__21965\,
            I => \N__21959\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__21962\,
            I => \N__21956\
        );

    \I__5276\ : Odrv4
    port map (
            O => \N__21959\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__5275\ : Odrv12
    port map (
            O => \N__21956\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__5274\ : CascadeMux
    port map (
            O => \N__21951\,
            I => \N__21938\
        );

    \I__5273\ : CascadeMux
    port map (
            O => \N__21950\,
            I => \N__21932\
        );

    \I__5272\ : InMux
    port map (
            O => \N__21949\,
            I => \N__21926\
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__21948\,
            I => \N__21923\
        );

    \I__5270\ : InMux
    port map (
            O => \N__21947\,
            I => \N__21920\
        );

    \I__5269\ : CascadeMux
    port map (
            O => \N__21946\,
            I => \N__21917\
        );

    \I__5268\ : InMux
    port map (
            O => \N__21945\,
            I => \N__21914\
        );

    \I__5267\ : CascadeMux
    port map (
            O => \N__21944\,
            I => \N__21907\
        );

    \I__5266\ : CascadeMux
    port map (
            O => \N__21943\,
            I => \N__21904\
        );

    \I__5265\ : CascadeMux
    port map (
            O => \N__21942\,
            I => \N__21900\
        );

    \I__5264\ : InMux
    port map (
            O => \N__21941\,
            I => \N__21890\
        );

    \I__5263\ : InMux
    port map (
            O => \N__21938\,
            I => \N__21890\
        );

    \I__5262\ : InMux
    port map (
            O => \N__21937\,
            I => \N__21890\
        );

    \I__5261\ : CascadeMux
    port map (
            O => \N__21936\,
            I => \N__21887\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__21935\,
            I => \N__21882\
        );

    \I__5259\ : InMux
    port map (
            O => \N__21932\,
            I => \N__21876\
        );

    \I__5258\ : InMux
    port map (
            O => \N__21931\,
            I => \N__21873\
        );

    \I__5257\ : InMux
    port map (
            O => \N__21930\,
            I => \N__21868\
        );

    \I__5256\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21868\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__21926\,
            I => \N__21865\
        );

    \I__5254\ : InMux
    port map (
            O => \N__21923\,
            I => \N__21862\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__21920\,
            I => \N__21859\
        );

    \I__5252\ : InMux
    port map (
            O => \N__21917\,
            I => \N__21856\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__21914\,
            I => \N__21853\
        );

    \I__5250\ : InMux
    port map (
            O => \N__21913\,
            I => \N__21840\
        );

    \I__5249\ : InMux
    port map (
            O => \N__21912\,
            I => \N__21840\
        );

    \I__5248\ : InMux
    port map (
            O => \N__21911\,
            I => \N__21840\
        );

    \I__5247\ : InMux
    port map (
            O => \N__21910\,
            I => \N__21840\
        );

    \I__5246\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21840\
        );

    \I__5245\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21840\
        );

    \I__5244\ : CascadeMux
    port map (
            O => \N__21903\,
            I => \N__21832\
        );

    \I__5243\ : InMux
    port map (
            O => \N__21900\,
            I => \N__21827\
        );

    \I__5242\ : InMux
    port map (
            O => \N__21899\,
            I => \N__21827\
        );

    \I__5241\ : InMux
    port map (
            O => \N__21898\,
            I => \N__21824\
        );

    \I__5240\ : InMux
    port map (
            O => \N__21897\,
            I => \N__21821\
        );

    \I__5239\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21817\
        );

    \I__5238\ : InMux
    port map (
            O => \N__21887\,
            I => \N__21802\
        );

    \I__5237\ : InMux
    port map (
            O => \N__21886\,
            I => \N__21802\
        );

    \I__5236\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21802\
        );

    \I__5235\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21802\
        );

    \I__5234\ : InMux
    port map (
            O => \N__21881\,
            I => \N__21802\
        );

    \I__5233\ : InMux
    port map (
            O => \N__21880\,
            I => \N__21802\
        );

    \I__5232\ : InMux
    port map (
            O => \N__21879\,
            I => \N__21802\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__21876\,
            I => \N__21787\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__21873\,
            I => \N__21787\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__21868\,
            I => \N__21787\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__21865\,
            I => \N__21787\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__21862\,
            I => \N__21787\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__21859\,
            I => \N__21787\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__21856\,
            I => \N__21787\
        );

    \I__5224\ : Span12Mux_s9_v
    port map (
            O => \N__21853\,
            I => \N__21782\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__21840\,
            I => \N__21782\
        );

    \I__5222\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21779\
        );

    \I__5221\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21774\
        );

    \I__5220\ : InMux
    port map (
            O => \N__21837\,
            I => \N__21774\
        );

    \I__5219\ : InMux
    port map (
            O => \N__21836\,
            I => \N__21767\
        );

    \I__5218\ : InMux
    port map (
            O => \N__21835\,
            I => \N__21767\
        );

    \I__5217\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21767\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__21827\,
            I => \N__21760\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21760\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__21821\,
            I => \N__21760\
        );

    \I__5213\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21757\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__21817\,
            I => \N__21750\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__21802\,
            I => \N__21750\
        );

    \I__5210\ : Span4Mux_v
    port map (
            O => \N__21787\,
            I => \N__21750\
        );

    \I__5209\ : Odrv12
    port map (
            O => \N__21782\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__21779\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__21774\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__21767\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5205\ : Odrv12
    port map (
            O => \N__21760\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__21757\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__21750\,
            I => \Lab_UT_dictrl_un1_next_state66_0\
        );

    \I__5202\ : InMux
    port map (
            O => \N__21735\,
            I => \N__21732\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__21732\,
            I => \Lab_UT.dictrl.m46_i_0_0_0\
        );

    \I__5200\ : InMux
    port map (
            O => \N__21729\,
            I => \N__21725\
        );

    \I__5199\ : InMux
    port map (
            O => \N__21728\,
            I => \N__21717\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__21725\,
            I => \N__21714\
        );

    \I__5197\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21709\
        );

    \I__5196\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21709\
        );

    \I__5195\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21706\
        );

    \I__5194\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21703\
        );

    \I__5193\ : InMux
    port map (
            O => \N__21720\,
            I => \N__21700\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__21717\,
            I => \N__21695\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__21714\,
            I => \N__21692\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__21709\,
            I => \N__21687\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21687\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__21703\,
            I => \N__21682\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__21700\,
            I => \N__21682\
        );

    \I__5186\ : InMux
    port map (
            O => \N__21699\,
            I => \N__21679\
        );

    \I__5185\ : InMux
    port map (
            O => \N__21698\,
            I => \N__21676\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__21695\,
            I => \N__21673\
        );

    \I__5183\ : Span4Mux_h
    port map (
            O => \N__21692\,
            I => \N__21664\
        );

    \I__5182\ : Span4Mux_v
    port map (
            O => \N__21687\,
            I => \N__21664\
        );

    \I__5181\ : Span4Mux_v
    port map (
            O => \N__21682\,
            I => \N__21664\
        );

    \I__5180\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21664\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__21676\,
            I => bu_rx_data_i_3_1
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__21673\,
            I => bu_rx_data_i_3_1
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__21664\,
            I => bu_rx_data_i_3_1
        );

    \I__5176\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21653\
        );

    \I__5175\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21645\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21642\
        );

    \I__5173\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21639\
        );

    \I__5172\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21632\
        );

    \I__5171\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21632\
        );

    \I__5170\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21632\
        );

    \I__5169\ : CascadeMux
    port map (
            O => \N__21648\,
            I => \N__21625\
        );

    \I__5168\ : LocalMux
    port map (
            O => \N__21645\,
            I => \N__21622\
        );

    \I__5167\ : Span4Mux_v
    port map (
            O => \N__21642\,
            I => \N__21614\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__21639\,
            I => \N__21614\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__21632\,
            I => \N__21614\
        );

    \I__5164\ : InMux
    port map (
            O => \N__21631\,
            I => \N__21607\
        );

    \I__5163\ : InMux
    port map (
            O => \N__21630\,
            I => \N__21607\
        );

    \I__5162\ : InMux
    port map (
            O => \N__21629\,
            I => \N__21607\
        );

    \I__5161\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21602\
        );

    \I__5160\ : InMux
    port map (
            O => \N__21625\,
            I => \N__21602\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__21622\,
            I => \N__21599\
        );

    \I__5158\ : InMux
    port map (
            O => \N__21621\,
            I => \N__21596\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__21614\,
            I => \N__21589\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__21607\,
            I => \N__21589\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__21602\,
            I => \N__21589\
        );

    \I__5154\ : Odrv4
    port map (
            O => \N__21599\,
            I => bu_rx_data_i_4_7
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21596\,
            I => bu_rx_data_i_4_7
        );

    \I__5152\ : Odrv4
    port map (
            O => \N__21589\,
            I => bu_rx_data_i_4_7
        );

    \I__5151\ : CascadeMux
    port map (
            O => \N__21582\,
            I => \N__21576\
        );

    \I__5150\ : CascadeMux
    port map (
            O => \N__21581\,
            I => \N__21573\
        );

    \I__5149\ : CascadeMux
    port map (
            O => \N__21580\,
            I => \N__21568\
        );

    \I__5148\ : CascadeMux
    port map (
            O => \N__21579\,
            I => \N__21565\
        );

    \I__5147\ : InMux
    port map (
            O => \N__21576\,
            I => \N__21562\
        );

    \I__5146\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21557\
        );

    \I__5145\ : CascadeMux
    port map (
            O => \N__21572\,
            I => \N__21553\
        );

    \I__5144\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21550\
        );

    \I__5143\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21547\
        );

    \I__5142\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21541\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21536\
        );

    \I__5140\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21533\
        );

    \I__5139\ : CascadeMux
    port map (
            O => \N__21560\,
            I => \N__21527\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__21557\,
            I => \N__21524\
        );

    \I__5137\ : InMux
    port map (
            O => \N__21556\,
            I => \N__21519\
        );

    \I__5136\ : InMux
    port map (
            O => \N__21553\,
            I => \N__21519\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__21550\,
            I => \N__21516\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21547\,
            I => \N__21513\
        );

    \I__5133\ : InMux
    port map (
            O => \N__21546\,
            I => \N__21506\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21545\,
            I => \N__21506\
        );

    \I__5131\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21506\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21503\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__21540\,
            I => \N__21499\
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__21539\,
            I => \N__21496\
        );

    \I__5127\ : Span4Mux_s2_h
    port map (
            O => \N__21536\,
            I => \N__21491\
        );

    \I__5126\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21491\
        );

    \I__5125\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21486\
        );

    \I__5124\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21486\
        );

    \I__5123\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21483\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21527\,
            I => \N__21480\
        );

    \I__5121\ : Span4Mux_s2_h
    port map (
            O => \N__21524\,
            I => \N__21475\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__21519\,
            I => \N__21475\
        );

    \I__5119\ : Span4Mux_s2_v
    port map (
            O => \N__21516\,
            I => \N__21466\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__21513\,
            I => \N__21466\
        );

    \I__5117\ : LocalMux
    port map (
            O => \N__21506\,
            I => \N__21466\
        );

    \I__5116\ : Span4Mux_h
    port map (
            O => \N__21503\,
            I => \N__21466\
        );

    \I__5115\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21459\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21459\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21459\
        );

    \I__5112\ : Span4Mux_h
    port map (
            O => \N__21491\,
            I => \N__21456\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21486\,
            I => bu_rx_data_6
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__21483\,
            I => bu_rx_data_6
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__21480\,
            I => bu_rx_data_6
        );

    \I__5108\ : Odrv4
    port map (
            O => \N__21475\,
            I => bu_rx_data_6
        );

    \I__5107\ : Odrv4
    port map (
            O => \N__21466\,
            I => bu_rx_data_6
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21459\,
            I => bu_rx_data_6
        );

    \I__5105\ : Odrv4
    port map (
            O => \N__21456\,
            I => bu_rx_data_6
        );

    \I__5104\ : InMux
    port map (
            O => \N__21441\,
            I => \N__21437\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21433\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__21437\,
            I => \N__21427\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21436\,
            I => \N__21424\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21433\,
            I => \N__21421\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21418\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__21431\,
            I => \N__21415\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21412\
        );

    \I__5096\ : Span12Mux_s6_h
    port map (
            O => \N__21427\,
            I => \N__21409\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21406\
        );

    \I__5094\ : Span4Mux_s3_h
    port map (
            O => \N__21421\,
            I => \N__21401\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21401\
        );

    \I__5092\ : InMux
    port map (
            O => \N__21415\,
            I => \N__21398\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__21412\,
            I => bu_rx_data_i_4_4
        );

    \I__5090\ : Odrv12
    port map (
            O => \N__21409\,
            I => bu_rx_data_i_4_4
        );

    \I__5089\ : Odrv4
    port map (
            O => \N__21406\,
            I => bu_rx_data_i_4_4
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__21401\,
            I => bu_rx_data_i_4_4
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__21398\,
            I => bu_rx_data_i_4_4
        );

    \I__5086\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21380\
        );

    \I__5085\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21377\
        );

    \I__5084\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21374\
        );

    \I__5083\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21371\
        );

    \I__5082\ : CascadeMux
    port map (
            O => \N__21383\,
            I => \N__21360\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21380\,
            I => \N__21349\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21377\,
            I => \N__21349\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21374\,
            I => \N__21346\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21337\
        );

    \I__5077\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21332\
        );

    \I__5076\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21332\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21368\,
            I => \N__21329\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21367\,
            I => \N__21326\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21366\,
            I => \N__21317\
        );

    \I__5072\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21317\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21317\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21317\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21308\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21359\,
            I => \N__21308\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21358\,
            I => \N__21308\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21357\,
            I => \N__21308\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21356\,
            I => \N__21303\
        );

    \I__5064\ : InMux
    port map (
            O => \N__21355\,
            I => \N__21303\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21300\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__21349\,
            I => \N__21289\
        );

    \I__5061\ : Span4Mux_v
    port map (
            O => \N__21346\,
            I => \N__21289\
        );

    \I__5060\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21284\
        );

    \I__5059\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21284\
        );

    \I__5058\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21281\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21274\
        );

    \I__5056\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21274\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21274\
        );

    \I__5054\ : Span4Mux_v
    port map (
            O => \N__21337\,
            I => \N__21271\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21264\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21264\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21264\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__21317\,
            I => \N__21255\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21255\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21255\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__21300\,
            I => \N__21255\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21299\,
            I => \N__21251\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21298\,
            I => \N__21248\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21297\,
            I => \N__21243\
        );

    \I__5043\ : InMux
    port map (
            O => \N__21296\,
            I => \N__21243\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21295\,
            I => \N__21240\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21237\
        );

    \I__5040\ : Span4Mux_h
    port map (
            O => \N__21289\,
            I => \N__21234\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21284\,
            I => \N__21227\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21281\,
            I => \N__21227\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21274\,
            I => \N__21227\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__21271\,
            I => \N__21220\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__21264\,
            I => \N__21220\
        );

    \I__5034\ : Span4Mux_v
    port map (
            O => \N__21255\,
            I => \N__21220\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21217\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21251\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__21248\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21243\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5029\ : LocalMux
    port map (
            O => \N__21240\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21237\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5027\ : Odrv4
    port map (
            O => \N__21234\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__21227\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5025\ : Odrv4
    port map (
            O => \N__21220\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5024\ : LocalMux
    port map (
            O => \N__21217\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \g0_3_4_cascade_\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21192\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21189\
        );

    \I__5020\ : Span4Mux_h
    port map (
            O => \N__21189\,
            I => \N__21186\
        );

    \I__5019\ : Odrv4
    port map (
            O => \N__21186\,
            I => g0_3_5
        );

    \I__5018\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21180\
        );

    \I__5017\ : LocalMux
    port map (
            O => \N__21180\,
            I => \Lab_UT.dictrl.g1Z0Z_2\
        );

    \I__5016\ : InMux
    port map (
            O => \N__21177\,
            I => \N__21174\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__21174\,
            I => \N__21171\
        );

    \I__5014\ : Odrv12
    port map (
            O => \N__21171\,
            I => \N_12\
        );

    \I__5013\ : CascadeMux
    port map (
            O => \N__21168\,
            I => \N__21164\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21159\
        );

    \I__5011\ : InMux
    port map (
            O => \N__21164\,
            I => \N__21159\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__21159\,
            I => \N__21154\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__21158\,
            I => \N__21150\
        );

    \I__5008\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21142\
        );

    \I__5007\ : Span4Mux_v
    port map (
            O => \N__21154\,
            I => \N__21139\
        );

    \I__5006\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21132\
        );

    \I__5005\ : InMux
    port map (
            O => \N__21150\,
            I => \N__21132\
        );

    \I__5004\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21132\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21148\,
            I => \N__21129\
        );

    \I__5002\ : CascadeMux
    port map (
            O => \N__21147\,
            I => \N__21126\
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__21146\,
            I => \N__21122\
        );

    \I__5000\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21117\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__21142\,
            I => \N__21108\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__21139\,
            I => \N__21108\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__21108\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__21129\,
            I => \N__21108\
        );

    \I__4995\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21103\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21103\
        );

    \I__4993\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21100\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21121\,
            I => \N__21095\
        );

    \I__4991\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21095\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__21117\,
            I => \N__21088\
        );

    \I__4989\ : Sp12to4
    port map (
            O => \N__21108\,
            I => \N__21088\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21103\,
            I => \N__21088\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21100\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__21095\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4985\ : Odrv12
    port map (
            O => \N__21088\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21078\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__21078\,
            I => \N__21074\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21077\,
            I => \N__21066\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__21074\,
            I => \N__21059\
        );

    \I__4980\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21048\
        );

    \I__4979\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21048\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21048\
        );

    \I__4977\ : InMux
    port map (
            O => \N__21070\,
            I => \N__21048\
        );

    \I__4976\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21048\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__21045\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21040\
        );

    \I__4973\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21040\
        );

    \I__4972\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21032\
        );

    \I__4971\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21029\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__21059\,
            I => \N__21026\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__21021\
        );

    \I__4968\ : Span4Mux_h
    port map (
            O => \N__21045\,
            I => \N__21021\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__21018\
        );

    \I__4966\ : InMux
    port map (
            O => \N__21039\,
            I => \N__21013\
        );

    \I__4965\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21013\
        );

    \I__4964\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21006\
        );

    \I__4963\ : InMux
    port map (
            O => \N__21036\,
            I => \N__21006\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21006\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__21032\,
            I => bu_rx_data_4
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21029\,
            I => bu_rx_data_4
        );

    \I__4959\ : Odrv4
    port map (
            O => \N__21026\,
            I => bu_rx_data_4
        );

    \I__4958\ : Odrv4
    port map (
            O => \N__21021\,
            I => bu_rx_data_4
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__21018\,
            I => bu_rx_data_4
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__21013\,
            I => bu_rx_data_4
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__21006\,
            I => bu_rx_data_4
        );

    \I__4954\ : InMux
    port map (
            O => \N__20991\,
            I => \N__20988\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__20988\,
            I => \Lab_UT.dictrl.N_13\
        );

    \I__4952\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20981\
        );

    \I__4951\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20977\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__20981\,
            I => \N__20974\
        );

    \I__4949\ : InMux
    port map (
            O => \N__20980\,
            I => \N__20971\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__20977\,
            I => \N__20959\
        );

    \I__4947\ : Span4Mux_s1_h
    port map (
            O => \N__20974\,
            I => \N__20956\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__20971\,
            I => \N__20953\
        );

    \I__4945\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20948\
        );

    \I__4944\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20948\
        );

    \I__4943\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20938\
        );

    \I__4942\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20938\
        );

    \I__4941\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20927\
        );

    \I__4940\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20927\
        );

    \I__4939\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20927\
        );

    \I__4938\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20927\
        );

    \I__4937\ : InMux
    port map (
            O => \N__20962\,
            I => \N__20927\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__20959\,
            I => \N__20924\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__20956\,
            I => \N__20921\
        );

    \I__4934\ : Span4Mux_s2_h
    port map (
            O => \N__20953\,
            I => \N__20916\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20916\
        );

    \I__4932\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20905\
        );

    \I__4931\ : InMux
    port map (
            O => \N__20946\,
            I => \N__20905\
        );

    \I__4930\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20905\
        );

    \I__4929\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20905\
        );

    \I__4928\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20905\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__20938\,
            I => bu_rx_data_5
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__20927\,
            I => bu_rx_data_5
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__20924\,
            I => bu_rx_data_5
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__20921\,
            I => bu_rx_data_5
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__20916\,
            I => bu_rx_data_5
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__20905\,
            I => bu_rx_data_5
        );

    \I__4921\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20889\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__20889\,
            I => \N__20883\
        );

    \I__4919\ : InMux
    port map (
            O => \N__20888\,
            I => \N__20880\
        );

    \I__4918\ : InMux
    port map (
            O => \N__20887\,
            I => \N__20872\
        );

    \I__4917\ : InMux
    port map (
            O => \N__20886\,
            I => \N__20869\
        );

    \I__4916\ : Span4Mux_s3_v
    port map (
            O => \N__20883\,
            I => \N__20866\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__20880\,
            I => \N__20861\
        );

    \I__4914\ : InMux
    port map (
            O => \N__20879\,
            I => \N__20858\
        );

    \I__4913\ : InMux
    port map (
            O => \N__20878\,
            I => \N__20848\
        );

    \I__4912\ : InMux
    port map (
            O => \N__20877\,
            I => \N__20845\
        );

    \I__4911\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20840\
        );

    \I__4910\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20840\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__20872\,
            I => \N__20837\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20834\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__20866\,
            I => \N__20830\
        );

    \I__4906\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20825\
        );

    \I__4905\ : InMux
    port map (
            O => \N__20864\,
            I => \N__20825\
        );

    \I__4904\ : Span4Mux_v
    port map (
            O => \N__20861\,
            I => \N__20820\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__20858\,
            I => \N__20820\
        );

    \I__4902\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20815\
        );

    \I__4901\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20815\
        );

    \I__4900\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20812\
        );

    \I__4899\ : InMux
    port map (
            O => \N__20854\,
            I => \N__20809\
        );

    \I__4898\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20806\
        );

    \I__4897\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20803\
        );

    \I__4896\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20796\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__20848\,
            I => \N__20793\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__20845\,
            I => \N__20784\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__20840\,
            I => \N__20784\
        );

    \I__4892\ : Span12Mux_s0_v
    port map (
            O => \N__20837\,
            I => \N__20784\
        );

    \I__4891\ : Sp12to4
    port map (
            O => \N__20834\,
            I => \N__20784\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__20833\,
            I => \N__20781\
        );

    \I__4889\ : Span4Mux_v
    port map (
            O => \N__20830\,
            I => \N__20774\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__20825\,
            I => \N__20774\
        );

    \I__4887\ : Span4Mux_h
    port map (
            O => \N__20820\,
            I => \N__20767\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__20815\,
            I => \N__20767\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20767\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__20809\,
            I => \N__20760\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__20806\,
            I => \N__20760\
        );

    \I__4882\ : LocalMux
    port map (
            O => \N__20803\,
            I => \N__20760\
        );

    \I__4881\ : InMux
    port map (
            O => \N__20802\,
            I => \N__20755\
        );

    \I__4880\ : InMux
    port map (
            O => \N__20801\,
            I => \N__20755\
        );

    \I__4879\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20752\
        );

    \I__4878\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20749\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20744\
        );

    \I__4876\ : Span4Mux_v
    port map (
            O => \N__20793\,
            I => \N__20744\
        );

    \I__4875\ : Span12Mux_v
    port map (
            O => \N__20784\,
            I => \N__20741\
        );

    \I__4874\ : InMux
    port map (
            O => \N__20781\,
            I => \N__20738\
        );

    \I__4873\ : InMux
    port map (
            O => \N__20780\,
            I => \N__20733\
        );

    \I__4872\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20733\
        );

    \I__4871\ : Span4Mux_h
    port map (
            O => \N__20774\,
            I => \N__20730\
        );

    \I__4870\ : Span4Mux_v
    port map (
            O => \N__20767\,
            I => \N__20723\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__20760\,
            I => \N__20723\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__20755\,
            I => \N__20723\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__20752\,
            I => bu_rx_data_1
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__20749\,
            I => bu_rx_data_1
        );

    \I__4865\ : Odrv4
    port map (
            O => \N__20744\,
            I => bu_rx_data_1
        );

    \I__4864\ : Odrv12
    port map (
            O => \N__20741\,
            I => bu_rx_data_1
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__20738\,
            I => bu_rx_data_1
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__20733\,
            I => bu_rx_data_1
        );

    \I__4861\ : Odrv4
    port map (
            O => \N__20730\,
            I => bu_rx_data_1
        );

    \I__4860\ : Odrv4
    port map (
            O => \N__20723\,
            I => bu_rx_data_1
        );

    \I__4859\ : CascadeMux
    port map (
            O => \N__20706\,
            I => \N__20699\
        );

    \I__4858\ : CascadeMux
    port map (
            O => \N__20705\,
            I => \N__20696\
        );

    \I__4857\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20693\
        );

    \I__4856\ : InMux
    port map (
            O => \N__20703\,
            I => \N__20688\
        );

    \I__4855\ : InMux
    port map (
            O => \N__20702\,
            I => \N__20688\
        );

    \I__4854\ : InMux
    port map (
            O => \N__20699\,
            I => \N__20685\
        );

    \I__4853\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20682\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__20693\,
            I => \N__20677\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__20688\,
            I => \N__20677\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__20685\,
            I => \N__20672\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__20682\,
            I => \N__20672\
        );

    \I__4848\ : Span4Mux_s3_v
    port map (
            O => \N__20677\,
            I => \N__20667\
        );

    \I__4847\ : Span4Mux_s3_h
    port map (
            O => \N__20672\,
            I => \N__20667\
        );

    \I__4846\ : Odrv4
    port map (
            O => \N__20667\,
            I => bu_rx_data_i_4_3_rep1
        );

    \I__4845\ : CascadeMux
    port map (
            O => \N__20664\,
            I => \N__20661\
        );

    \I__4844\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20657\
        );

    \I__4843\ : InMux
    port map (
            O => \N__20660\,
            I => \N__20653\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__20657\,
            I => \N__20648\
        );

    \I__4841\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20645\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20642\
        );

    \I__4839\ : InMux
    port map (
            O => \N__20652\,
            I => \N__20638\
        );

    \I__4838\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20633\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__20648\,
            I => \N__20629\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__20645\,
            I => \N__20626\
        );

    \I__4835\ : Span4Mux_h
    port map (
            O => \N__20642\,
            I => \N__20623\
        );

    \I__4834\ : InMux
    port map (
            O => \N__20641\,
            I => \N__20620\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__20638\,
            I => \N__20617\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20637\,
            I => \N__20612\
        );

    \I__4831\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20612\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20609\
        );

    \I__4829\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20606\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__20629\,
            I => bu_rx_data_i_4_2
        );

    \I__4827\ : Odrv12
    port map (
            O => \N__20626\,
            I => bu_rx_data_i_4_2
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__20623\,
            I => bu_rx_data_i_4_2
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__20620\,
            I => bu_rx_data_i_4_2
        );

    \I__4824\ : Odrv4
    port map (
            O => \N__20617\,
            I => bu_rx_data_i_4_2
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__20612\,
            I => bu_rx_data_i_4_2
        );

    \I__4822\ : Odrv12
    port map (
            O => \N__20609\,
            I => bu_rx_data_i_4_2
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__20606\,
            I => bu_rx_data_i_4_2
        );

    \I__4820\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20586\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__20586\,
            I => m46_i_0_a3_2
        );

    \I__4818\ : InMux
    port map (
            O => \N__20583\,
            I => \N__20578\
        );

    \I__4817\ : InMux
    port map (
            O => \N__20582\,
            I => \N__20573\
        );

    \I__4816\ : InMux
    port map (
            O => \N__20581\,
            I => \N__20573\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__20578\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__20573\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__4813\ : CascadeMux
    port map (
            O => \N__20568\,
            I => \N__20565\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20559\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20552\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20563\,
            I => \N__20552\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20552\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20559\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__4807\ : LocalMux
    port map (
            O => \N__20552\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20547\,
            I => \N__20542\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20546\,
            I => \N__20537\
        );

    \I__4804\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20537\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20542\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__4802\ : LocalMux
    port map (
            O => \N__20537\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__4801\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20526\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20526\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__20526\,
            I => \N__20523\
        );

    \I__4798\ : Span4Mux_s2_h
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__4797\ : Odrv4
    port map (
            O => \N__20520\,
            I => \Lab_UT.dictrl.N_90\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20511\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20506\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20510\,
            I => \N__20501\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20509\,
            I => \N__20501\
        );

    \I__4791\ : Span4Mux_v
    port map (
            O => \N__20506\,
            I => \N__20498\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20501\,
            I => \N__20495\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__20498\,
            I => \Lab_UT.dictrl.N_119\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__20495\,
            I => \Lab_UT.dictrl.N_119\
        );

    \I__4787\ : CascadeMux
    port map (
            O => \N__20490\,
            I => \Lab_UT.dictrl.N_139_cascade_\
        );

    \I__4786\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20482\
        );

    \I__4785\ : InMux
    port map (
            O => \N__20486\,
            I => \N__20476\
        );

    \I__4784\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20476\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__20482\,
            I => \N__20473\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20470\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20465\
        );

    \I__4780\ : Span4Mux_v
    port map (
            O => \N__20473\,
            I => \N__20460\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20460\
        );

    \I__4778\ : InMux
    port map (
            O => \N__20469\,
            I => \N__20455\
        );

    \I__4777\ : InMux
    port map (
            O => \N__20468\,
            I => \N__20455\
        );

    \I__4776\ : Span4Mux_h
    port map (
            O => \N__20465\,
            I => \N__20452\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__20460\,
            I => \N__20449\
        );

    \I__4774\ : LocalMux
    port map (
            O => \N__20455\,
            I => \N__20446\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__20452\,
            I => \Lab_UT.dictrl.N_116_mux\
        );

    \I__4772\ : Odrv4
    port map (
            O => \N__20449\,
            I => \Lab_UT.dictrl.N_116_mux\
        );

    \I__4771\ : Odrv4
    port map (
            O => \N__20446\,
            I => \Lab_UT.dictrl.N_116_mux\
        );

    \I__4770\ : InMux
    port map (
            O => \N__20439\,
            I => \N__20436\
        );

    \I__4769\ : LocalMux
    port map (
            O => \N__20436\,
            I => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\
        );

    \I__4768\ : CascadeMux
    port map (
            O => \N__20433\,
            I => \N__20430\
        );

    \I__4767\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20427\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__20427\,
            I => \N__20424\
        );

    \I__4765\ : Span4Mux_s2_h
    port map (
            O => \N__20424\,
            I => \N__20421\
        );

    \I__4764\ : Odrv4
    port map (
            O => \N__20421\,
            I => \Lab_UT.dictrl.g2_2\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20415\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__20415\,
            I => \N__20410\
        );

    \I__4761\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20407\
        );

    \I__4760\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20404\
        );

    \I__4759\ : Span4Mux_s2_h
    port map (
            O => \N__20410\,
            I => \N__20401\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20407\,
            I => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__20404\,
            I => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__20401\,
            I => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20391\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20391\,
            I => \N__20388\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__20388\,
            I => \Lab_UT.dictrl.N_5_1\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20385\,
            I => \N__20382\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__20382\,
            I => \N__20379\
        );

    \I__4750\ : Span4Mux_s2_h
    port map (
            O => \N__20379\,
            I => \N__20376\
        );

    \I__4749\ : Odrv4
    port map (
            O => \N__20376\,
            I => \Lab_UT.dictrl.g2_0_0_0_0\
        );

    \I__4748\ : CascadeMux
    port map (
            O => \N__20373\,
            I => \N__20363\
        );

    \I__4747\ : CascadeMux
    port map (
            O => \N__20372\,
            I => \N__20360\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20356\
        );

    \I__4745\ : CascadeMux
    port map (
            O => \N__20370\,
            I => \N__20353\
        );

    \I__4744\ : CascadeMux
    port map (
            O => \N__20369\,
            I => \N__20348\
        );

    \I__4743\ : CascadeMux
    port map (
            O => \N__20368\,
            I => \N__20342\
        );

    \I__4742\ : CascadeMux
    port map (
            O => \N__20367\,
            I => \N__20338\
        );

    \I__4741\ : CascadeMux
    port map (
            O => \N__20366\,
            I => \N__20333\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20329\
        );

    \I__4739\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20326\
        );

    \I__4738\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20323\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20320\
        );

    \I__4736\ : InMux
    port map (
            O => \N__20353\,
            I => \N__20317\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20352\,
            I => \N__20312\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20312\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20309\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20347\,
            I => \N__20306\
        );

    \I__4731\ : CascadeMux
    port map (
            O => \N__20346\,
            I => \N__20301\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20345\,
            I => \N__20295\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20295\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20292\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20287\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20337\,
            I => \N__20287\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20336\,
            I => \N__20282\
        );

    \I__4724\ : InMux
    port map (
            O => \N__20333\,
            I => \N__20282\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__20332\,
            I => \N__20279\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__20329\,
            I => \N__20274\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20326\,
            I => \N__20274\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20323\,
            I => \N__20265\
        );

    \I__4719\ : Span4Mux_v
    port map (
            O => \N__20320\,
            I => \N__20265\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20265\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__20312\,
            I => \N__20265\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__20309\,
            I => \N__20262\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20259\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20305\,
            I => \N__20252\
        );

    \I__4713\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20252\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20252\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20249\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__20295\,
            I => \N__20246\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__20292\,
            I => \N__20241\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20287\,
            I => \N__20241\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20282\,
            I => \N__20238\
        );

    \I__4706\ : InMux
    port map (
            O => \N__20279\,
            I => \N__20235\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__20274\,
            I => \N__20230\
        );

    \I__4704\ : Span4Mux_v
    port map (
            O => \N__20265\,
            I => \N__20230\
        );

    \I__4703\ : Span4Mux_s3_h
    port map (
            O => \N__20262\,
            I => \N__20221\
        );

    \I__4702\ : Span4Mux_v
    port map (
            O => \N__20259\,
            I => \N__20221\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20252\,
            I => \N__20221\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20249\,
            I => \N__20221\
        );

    \I__4699\ : Span4Mux_h
    port map (
            O => \N__20246\,
            I => \N__20218\
        );

    \I__4698\ : Odrv12
    port map (
            O => \N__20241\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__20238\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20235\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__20230\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__20221\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__20218\,
            I => \Lab_UT.dictrl.stateZ0Z_3\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20202\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20202\,
            I => \N__20199\
        );

    \I__4690\ : Span4Mux_s2_h
    port map (
            O => \N__20199\,
            I => \N__20196\
        );

    \I__4689\ : Odrv4
    port map (
            O => \N__20196\,
            I => \Lab_UT.dictrl.N_103_0_0_0\
        );

    \I__4688\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20190\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20190\,
            I => \Lab_UT.dictrl.N_1302_1_0_0\
        );

    \I__4686\ : CascadeMux
    port map (
            O => \N__20187\,
            I => \Lab_UT.dictrl.N_119_0_0_0_cascade_\
        );

    \I__4685\ : InMux
    port map (
            O => \N__20184\,
            I => \N__20169\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20183\,
            I => \N__20169\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20165\
        );

    \I__4682\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20160\
        );

    \I__4681\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20160\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__20179\,
            I => \N__20155\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__20178\,
            I => \N__20152\
        );

    \I__4678\ : CascadeMux
    port map (
            O => \N__20177\,
            I => \N__20148\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20145\
        );

    \I__4676\ : InMux
    port map (
            O => \N__20175\,
            I => \N__20142\
        );

    \I__4675\ : CascadeMux
    port map (
            O => \N__20174\,
            I => \N__20138\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20135\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20125\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20165\,
            I => \N__20122\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20119\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20113\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20113\
        );

    \I__4668\ : InMux
    port map (
            O => \N__20155\,
            I => \N__20104\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20152\,
            I => \N__20104\
        );

    \I__4666\ : InMux
    port map (
            O => \N__20151\,
            I => \N__20104\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20148\,
            I => \N__20104\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__20145\,
            I => \N__20099\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__20142\,
            I => \N__20099\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20096\
        );

    \I__4661\ : InMux
    port map (
            O => \N__20138\,
            I => \N__20092\
        );

    \I__4660\ : Span4Mux_s3_h
    port map (
            O => \N__20135\,
            I => \N__20089\
        );

    \I__4659\ : InMux
    port map (
            O => \N__20134\,
            I => \N__20078\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20133\,
            I => \N__20078\
        );

    \I__4657\ : InMux
    port map (
            O => \N__20132\,
            I => \N__20078\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20131\,
            I => \N__20078\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20130\,
            I => \N__20078\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20073\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20073\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20125\,
            I => \N__20066\
        );

    \I__4651\ : Span4Mux_s3_h
    port map (
            O => \N__20122\,
            I => \N__20066\
        );

    \I__4650\ : Span4Mux_s3_h
    port map (
            O => \N__20119\,
            I => \N__20066\
        );

    \I__4649\ : InMux
    port map (
            O => \N__20118\,
            I => \N__20063\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20054\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20054\
        );

    \I__4646\ : Span12Mux_s9_v
    port map (
            O => \N__20099\,
            I => \N__20054\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__20096\,
            I => \N__20054\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20095\,
            I => \N__20051\
        );

    \I__4643\ : LocalMux
    port map (
            O => \N__20092\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__20089\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20078\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20073\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4639\ : Odrv4
    port map (
            O => \N__20066\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__20063\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4637\ : Odrv12
    port map (
            O => \N__20054\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__20051\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__20034\,
            I => \N__20031\
        );

    \I__4634\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20025\
        );

    \I__4633\ : InMux
    port map (
            O => \N__20030\,
            I => \N__20025\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__20022\
        );

    \I__4631\ : Span4Mux_h
    port map (
            O => \N__20022\,
            I => \N__20019\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__20019\,
            I => \Lab_UT.dictrl.g1Z0Z_4\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__20016\,
            I => \Lab_UT_dictrl_next_state_3_cascade_\
        );

    \I__4628\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20010\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20010\,
            I => \Lab_UT.dictrl.state_ret_12_RNOZ0Z_3\
        );

    \I__4626\ : InMux
    port map (
            O => \N__20007\,
            I => \N__20004\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__20004\,
            I => \Lab_UT.dictrl.next_state_0_0_2\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20001\,
            I => \N__19998\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__19998\,
            I => \Lab_UT.dictrl.state_ret_12_RNOZ0Z_4\
        );

    \I__4622\ : InMux
    port map (
            O => \N__19995\,
            I => \N__19992\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__19992\,
            I => \Lab_UT.dictrl.state_ret_12and_a0_1\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__19989\,
            I => \N__19985\
        );

    \I__4619\ : CascadeMux
    port map (
            O => \N__19988\,
            I => \N__19982\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19974\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19974\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19974\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__19974\,
            I => \N__19969\
        );

    \I__4614\ : InMux
    port map (
            O => \N__19973\,
            I => \N__19966\
        );

    \I__4613\ : InMux
    port map (
            O => \N__19972\,
            I => \N__19963\
        );

    \I__4612\ : Span4Mux_s3_h
    port map (
            O => \N__19969\,
            I => \N__19958\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19966\,
            I => \N__19958\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__19963\,
            I => \N__19955\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__19958\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__4608\ : Odrv4
    port map (
            O => \N__19955\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \Lab_UT.dictrl.state_ret_12and_0_0_cascade_\
        );

    \I__4606\ : InMux
    port map (
            O => \N__19947\,
            I => \N__19939\
        );

    \I__4605\ : InMux
    port map (
            O => \N__19946\,
            I => \N__19932\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19932\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19944\,
            I => \N__19932\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19943\,
            I => \N__19929\
        );

    \I__4601\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19926\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19923\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__19932\,
            I => \N__19920\
        );

    \I__4598\ : LocalMux
    port map (
            O => \N__19929\,
            I => \N__19917\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19914\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__19923\,
            I => \N__19911\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__19920\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__19917\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__19914\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4592\ : Odrv4
    port map (
            O => \N__19911\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4591\ : CascadeMux
    port map (
            O => \N__19902\,
            I => \N__19896\
        );

    \I__4590\ : CascadeMux
    port map (
            O => \N__19901\,
            I => \N__19890\
        );

    \I__4589\ : InMux
    port map (
            O => \N__19900\,
            I => \N__19884\
        );

    \I__4588\ : InMux
    port map (
            O => \N__19899\,
            I => \N__19879\
        );

    \I__4587\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19876\
        );

    \I__4586\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19873\
        );

    \I__4585\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19870\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__19893\,
            I => \N__19867\
        );

    \I__4583\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19860\
        );

    \I__4582\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19860\
        );

    \I__4581\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19860\
        );

    \I__4580\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19857\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__19884\,
            I => \N__19854\
        );

    \I__4578\ : InMux
    port map (
            O => \N__19883\,
            I => \N__19851\
        );

    \I__4577\ : InMux
    port map (
            O => \N__19882\,
            I => \N__19848\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__19879\,
            I => \N__19845\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__19876\,
            I => \N__19838\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__19873\,
            I => \N__19838\
        );

    \I__4573\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19838\
        );

    \I__4572\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19835\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__19860\,
            I => \N__19832\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19829\
        );

    \I__4569\ : Span4Mux_v
    port map (
            O => \N__19854\,
            I => \N__19822\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__19851\,
            I => \N__19822\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__19848\,
            I => \N__19822\
        );

    \I__4566\ : Span4Mux_v
    port map (
            O => \N__19845\,
            I => \N__19817\
        );

    \I__4565\ : Span4Mux_v
    port map (
            O => \N__19838\,
            I => \N__19817\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__19835\,
            I => \N__19814\
        );

    \I__4563\ : Span4Mux_h
    port map (
            O => \N__19832\,
            I => \N__19807\
        );

    \I__4562\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19807\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__19822\,
            I => \N__19807\
        );

    \I__4560\ : Odrv4
    port map (
            O => \N__19817\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4559\ : Odrv12
    port map (
            O => \N__19814\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__19807\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4557\ : InMux
    port map (
            O => \N__19800\,
            I => \N__19796\
        );

    \I__4556\ : InMux
    port map (
            O => \N__19799\,
            I => \N__19793\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19790\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__19793\,
            I => \N__19785\
        );

    \I__4553\ : Span4Mux_v
    port map (
            O => \N__19790\,
            I => \N__19782\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__19789\,
            I => \N__19778\
        );

    \I__4551\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19771\
        );

    \I__4550\ : Span4Mux_h
    port map (
            O => \N__19785\,
            I => \N__19766\
        );

    \I__4549\ : Span4Mux_v
    port map (
            O => \N__19782\,
            I => \N__19766\
        );

    \I__4548\ : InMux
    port map (
            O => \N__19781\,
            I => \N__19755\
        );

    \I__4547\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19755\
        );

    \I__4546\ : InMux
    port map (
            O => \N__19777\,
            I => \N__19755\
        );

    \I__4545\ : InMux
    port map (
            O => \N__19776\,
            I => \N__19755\
        );

    \I__4544\ : InMux
    port map (
            O => \N__19775\,
            I => \N__19755\
        );

    \I__4543\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19752\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__19771\,
            I => \N__19749\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__19766\,
            I => \buart__rx_bitcount_3\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__19755\,
            I => \buart__rx_bitcount_3\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__19752\,
            I => \buart__rx_bitcount_3\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__19749\,
            I => \buart__rx_bitcount_3\
        );

    \I__4537\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19737\
        );

    \I__4536\ : LocalMux
    port map (
            O => \N__19737\,
            I => \N__19733\
        );

    \I__4535\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19730\
        );

    \I__4534\ : Span4Mux_h
    port map (
            O => \N__19733\,
            I => \N__19727\
        );

    \I__4533\ : LocalMux
    port map (
            O => \N__19730\,
            I => \N__19722\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__19727\,
            I => \N__19719\
        );

    \I__4531\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19714\
        );

    \I__4530\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19714\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__19722\,
            I => \N__19711\
        );

    \I__4528\ : Odrv4
    port map (
            O => \N__19719\,
            I => \buart__rx_valid_3\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__19714\,
            I => \buart__rx_valid_3\
        );

    \I__4526\ : Odrv4
    port map (
            O => \N__19711\,
            I => \buart__rx_valid_3\
        );

    \I__4525\ : InMux
    port map (
            O => \N__19704\,
            I => \N__19693\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19703\,
            I => \N__19693\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19693\
        );

    \I__4522\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19690\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19687\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__19693\,
            I => \N__19684\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__19690\,
            I => \N__19681\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__19687\,
            I => \N__19678\
        );

    \I__4517\ : Span4Mux_h
    port map (
            O => \N__19684\,
            I => \N__19673\
        );

    \I__4516\ : Span4Mux_h
    port map (
            O => \N__19681\,
            I => \N__19670\
        );

    \I__4515\ : Span4Mux_h
    port map (
            O => \N__19678\,
            I => \N__19667\
        );

    \I__4514\ : InMux
    port map (
            O => \N__19677\,
            I => \N__19664\
        );

    \I__4513\ : InMux
    port map (
            O => \N__19676\,
            I => \N__19661\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__19673\,
            I => \Lab_UT_dictrl_next_state_3\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__19670\,
            I => \Lab_UT_dictrl_next_state_3\
        );

    \I__4510\ : Odrv4
    port map (
            O => \N__19667\,
            I => \Lab_UT_dictrl_next_state_3\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__19664\,
            I => \Lab_UT_dictrl_next_state_3\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19661\,
            I => \Lab_UT_dictrl_next_state_3\
        );

    \I__4507\ : CascadeMux
    port map (
            O => \N__19650\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__4506\ : IoInMux
    port map (
            O => \N__19647\,
            I => \N__19641\
        );

    \I__4505\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19635\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19630\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19644\,
            I => \N__19630\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__19641\,
            I => \N__19627\
        );

    \I__4501\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19620\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19639\,
            I => \N__19620\
        );

    \I__4499\ : InMux
    port map (
            O => \N__19638\,
            I => \N__19620\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19617\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19630\,
            I => \N__19614\
        );

    \I__4496\ : Span4Mux_s2_h
    port map (
            O => \N__19627\,
            I => \N__19611\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19620\,
            I => \N__19608\
        );

    \I__4494\ : Span4Mux_h
    port map (
            O => \N__19617\,
            I => \N__19605\
        );

    \I__4493\ : Span4Mux_v
    port map (
            O => \N__19614\,
            I => \N__19600\
        );

    \I__4492\ : Span4Mux_h
    port map (
            O => \N__19611\,
            I => \N__19600\
        );

    \I__4491\ : Odrv12
    port map (
            O => \N__19608\,
            I => rst
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__19605\,
            I => rst
        );

    \I__4489\ : Odrv4
    port map (
            O => \N__19600\,
            I => rst
        );

    \I__4488\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19590\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__19590\,
            I => \N__19587\
        );

    \I__4486\ : Span4Mux_v
    port map (
            O => \N__19587\,
            I => \N__19583\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19586\,
            I => \N__19580\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__19583\,
            I => \Lab_UT.dictrl.N_119_mux\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__19580\,
            I => \Lab_UT.dictrl.N_119_mux\
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__19575\,
            I => \Lab_UT.dictrl.i9_mux_cascade_\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19568\
        );

    \I__4480\ : InMux
    port map (
            O => \N__19571\,
            I => \N__19565\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__19568\,
            I => \N__19562\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19565\,
            I => \N__19559\
        );

    \I__4477\ : Odrv12
    port map (
            O => \N__19562\,
            I => \Lab_UT.dictrl.N_94\
        );

    \I__4476\ : Odrv12
    port map (
            O => \N__19559\,
            I => \Lab_UT.dictrl.N_94\
        );

    \I__4475\ : CascadeMux
    port map (
            O => \N__19554\,
            I => \N__19551\
        );

    \I__4474\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19548\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19548\,
            I => \N__19542\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19547\,
            I => \N__19539\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19546\,
            I => \N__19536\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19533\
        );

    \I__4469\ : Span4Mux_v
    port map (
            O => \N__19542\,
            I => \N__19526\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__19539\,
            I => \N__19526\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19536\,
            I => \N__19526\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19533\,
            I => \N__19523\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__19526\,
            I => \N__19520\
        );

    \I__4464\ : Span4Mux_s1_h
    port map (
            O => \N__19523\,
            I => \N__19517\
        );

    \I__4463\ : Odrv4
    port map (
            O => \N__19520\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__4462\ : Odrv4
    port map (
            O => \N__19517\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__19512\,
            I => \Lab_UT.dictrl.N_107_mux_cascade_\
        );

    \I__4460\ : InMux
    port map (
            O => \N__19509\,
            I => \N__19506\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19506\,
            I => m89_am
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__19503\,
            I => \N__19499\
        );

    \I__4457\ : InMux
    port map (
            O => \N__19502\,
            I => \N__19491\
        );

    \I__4456\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19491\
        );

    \I__4455\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19491\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19488\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__19488\,
            I => \N__19484\
        );

    \I__4452\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19481\
        );

    \I__4451\ : Sp12to4
    port map (
            O => \N__19484\,
            I => \N__19478\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__19481\,
            I => \buart__rx_hh_0\
        );

    \I__4449\ : Odrv12
    port map (
            O => \N__19478\,
            I => \buart__rx_hh_0\
        );

    \I__4448\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19463\
        );

    \I__4447\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19463\
        );

    \I__4446\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19456\
        );

    \I__4445\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19456\
        );

    \I__4444\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19456\
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19453\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19463\,
            I => \N__19448\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19456\,
            I => \N__19445\
        );

    \I__4440\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19438\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19438\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19438\
        );

    \I__4437\ : Span4Mux_h
    port map (
            O => \N__19448\,
            I => \N__19433\
        );

    \I__4436\ : Span4Mux_v
    port map (
            O => \N__19445\,
            I => \N__19433\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19430\
        );

    \I__4434\ : Span4Mux_v
    port map (
            O => \N__19433\,
            I => \N__19425\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__19430\,
            I => \N__19425\
        );

    \I__4432\ : Sp12to4
    port map (
            O => \N__19425\,
            I => \N__19422\
        );

    \I__4431\ : Odrv12
    port map (
            O => \N__19422\,
            I => \buart__rx_hh_1\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19407\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19407\
        );

    \I__4428\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19407\
        );

    \I__4427\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19407\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19407\,
            I => \Lab_UT.dictrl.N_102_mux\
        );

    \I__4425\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19396\
        );

    \I__4424\ : InMux
    port map (
            O => \N__19403\,
            I => \N__19396\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19393\
        );

    \I__4422\ : InMux
    port map (
            O => \N__19401\,
            I => \N__19390\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__19396\,
            I => \N__19385\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19385\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19390\,
            I => \buart__rx_N_27_0_i\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__19385\,
            I => \buart__rx_N_27_0_i\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__19380\,
            I => \buart__rx_startbit_cascade_\
        );

    \I__4416\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19373\
        );

    \I__4415\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19367\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__19373\,
            I => \N__19364\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19357\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19371\,
            I => \N__19357\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19357\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19367\,
            I => \buart__rx_bitcount_0\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__19364\,
            I => \buart__rx_bitcount_0\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19357\,
            I => \buart__rx_bitcount_0\
        );

    \I__4407\ : CEMux
    port map (
            O => \N__19350\,
            I => \N__19346\
        );

    \I__4406\ : CEMux
    port map (
            O => \N__19349\,
            I => \N__19342\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__19346\,
            I => \N__19339\
        );

    \I__4404\ : CEMux
    port map (
            O => \N__19345\,
            I => \N__19336\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19342\,
            I => \N__19333\
        );

    \I__4402\ : Span4Mux_h
    port map (
            O => \N__19339\,
            I => \N__19330\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__19336\,
            I => \N__19327\
        );

    \I__4400\ : Odrv12
    port map (
            O => \N__19333\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__4399\ : Odrv4
    port map (
            O => \N__19330\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__4398\ : Odrv4
    port map (
            O => \N__19327\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19317\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__19317\,
            I => \N__19314\
        );

    \I__4395\ : Span4Mux_h
    port map (
            O => \N__19314\,
            I => \N__19311\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__19311\,
            I => \Lab_UT.dictrl.i9_mux_0_0\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19308\,
            I => \N__19305\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19305\,
            I => \N__19302\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__19302\,
            I => \N__19299\
        );

    \I__4390\ : Odrv4
    port map (
            O => \N__19299\,
            I => \Lab_UT.dictrl.N_94_0_0\
        );

    \I__4389\ : CascadeMux
    port map (
            O => \N__19296\,
            I => \Lab_UT.dictrl.N_2000_0_0_cascade_\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19293\,
            I => \N__19285\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19292\,
            I => \N__19285\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19291\,
            I => \N__19280\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19280\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19274\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19280\,
            I => \N__19274\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19279\,
            I => \N__19271\
        );

    \I__4381\ : Span4Mux_v
    port map (
            O => \N__19274\,
            I => \N__19268\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__19271\,
            I => \N__19265\
        );

    \I__4379\ : Odrv4
    port map (
            O => \N__19268\,
            I => \Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3\
        );

    \I__4378\ : Odrv12
    port map (
            O => \N__19265\,
            I => \Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19247\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19247\
        );

    \I__4375\ : InMux
    port map (
            O => \N__19258\,
            I => \N__19247\
        );

    \I__4374\ : InMux
    port map (
            O => \N__19257\,
            I => \N__19247\
        );

    \I__4373\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19244\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__19247\,
            I => \N__19239\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19244\,
            I => \N__19239\
        );

    \I__4370\ : Odrv12
    port map (
            O => \N__19239\,
            I => \Lab_UT.dictrl.N_121_mux\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19236\,
            I => \N__19233\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19230\
        );

    \I__4367\ : Span4Mux_h
    port map (
            O => \N__19230\,
            I => \N__19227\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__19227\,
            I => \N__19224\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__19224\,
            I => \Lab_UT.dictrl.N_83\
        );

    \I__4364\ : CascadeMux
    port map (
            O => \N__19221\,
            I => \Lab_UT.dictrl.N_194_cascade_\
        );

    \I__4363\ : IoInMux
    port map (
            O => \N__19218\,
            I => \N__19215\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19215\,
            I => \N__19212\
        );

    \I__4361\ : IoSpan4Mux
    port map (
            O => \N__19212\,
            I => \N__19209\
        );

    \I__4360\ : Span4Mux_s2_v
    port map (
            O => \N__19209\,
            I => \N__19206\
        );

    \I__4359\ : Sp12to4
    port map (
            O => \N__19206\,
            I => \N__19203\
        );

    \I__4358\ : Odrv12
    port map (
            O => \N__19203\,
            I => \buart__rx_sample\
        );

    \I__4357\ : CascadeMux
    port map (
            O => \N__19200\,
            I => \N__19194\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19187\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19187\
        );

    \I__4354\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19187\
        );

    \I__4353\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19183\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19180\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19177\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__19183\,
            I => \N__19172\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__19180\,
            I => \N__19172\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__19177\,
            I => \buart__rx_bitcount_2\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__19172\,
            I => \buart__rx_bitcount_2\
        );

    \I__4346\ : CascadeMux
    port map (
            O => \N__19167\,
            I => \N__19162\
        );

    \I__4345\ : CascadeMux
    port map (
            O => \N__19166\,
            I => \N__19158\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19151\
        );

    \I__4343\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19151\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19151\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19148\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19151\,
            I => \N__19144\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__19148\,
            I => \N__19141\
        );

    \I__4338\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19138\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__19144\,
            I => \N__19135\
        );

    \I__4336\ : Odrv4
    port map (
            O => \N__19141\,
            I => \buart__rx_bitcount_1\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19138\,
            I => \buart__rx_bitcount_1\
        );

    \I__4334\ : Odrv4
    port map (
            O => \N__19135\,
            I => \buart__rx_bitcount_1\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__19128\,
            I => \N__19123\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19115\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19115\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19115\
        );

    \I__4329\ : CascadeMux
    port map (
            O => \N__19122\,
            I => \N__19112\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19115\,
            I => \N__19109\
        );

    \I__4327\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19106\
        );

    \I__4326\ : Span4Mux_s2_h
    port map (
            O => \N__19109\,
            I => \N__19103\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19106\,
            I => \buart__rx_bitcount_4\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__19103\,
            I => \buart__rx_bitcount_4\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19095\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19095\,
            I => m89_bm
        );

    \I__4321\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19089\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19089\,
            I => \N__19086\
        );

    \I__4319\ : Odrv4
    port map (
            O => \N__19086\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__19083\,
            I => \buart__rx_N_27_0_i_cascade_\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19072\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19072\
        );

    \I__4315\ : CascadeMux
    port map (
            O => \N__19078\,
            I => \N__19069\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__19077\,
            I => \N__19065\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19062\
        );

    \I__4312\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19057\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19057\
        );

    \I__4310\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19054\
        );

    \I__4309\ : Odrv4
    port map (
            O => \N__19062\,
            I => \Lab_UT.dictrl.N_98_mux\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19057\,
            I => \Lab_UT.dictrl.N_98_mux\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__19054\,
            I => \Lab_UT.dictrl.N_98_mux\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19041\
        );

    \I__4305\ : InMux
    port map (
            O => \N__19046\,
            I => \N__19036\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19045\,
            I => \N__19036\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19044\,
            I => \N__19033\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__19041\,
            I => \Lab_UT.dictrl.N_84\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19036\,
            I => \Lab_UT.dictrl.N_84\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19033\,
            I => \Lab_UT.dictrl.N_84\
        );

    \I__4299\ : InMux
    port map (
            O => \N__19026\,
            I => \N__19021\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \N__19018\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19013\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19021\,
            I => \N__19010\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19003\
        );

    \I__4294\ : InMux
    port map (
            O => \N__19017\,
            I => \N__19003\
        );

    \I__4293\ : InMux
    port map (
            O => \N__19016\,
            I => \N__19003\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19013\,
            I => \N__19000\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__19010\,
            I => \N__18995\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__19003\,
            I => \N__18995\
        );

    \I__4289\ : Odrv12
    port map (
            O => \N__19000\,
            I => \Lab_UT.dictrl.N_89\
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__18995\,
            I => \Lab_UT.dictrl.N_89\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18990\,
            I => \N__18987\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__18987\,
            I => \Lab_UT.dictrl.m68_1\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__18984\,
            I => \Lab_UT.dictrl.N_89_cascade_\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18981\,
            I => \N__18977\
        );

    \I__4283\ : InMux
    port map (
            O => \N__18980\,
            I => \N__18974\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18971\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__18974\,
            I => \N__18968\
        );

    \I__4280\ : Span4Mux_h
    port map (
            O => \N__18971\,
            I => \N__18965\
        );

    \I__4279\ : Odrv12
    port map (
            O => \N__18968\,
            I => \Lab_UT.dictrl.N_99_mux\
        );

    \I__4278\ : Odrv4
    port map (
            O => \N__18965\,
            I => \Lab_UT.dictrl.N_99_mux\
        );

    \I__4277\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18954\
        );

    \I__4276\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18954\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18954\,
            I => \Lab_UT.dictrl.N_102\
        );

    \I__4274\ : InMux
    port map (
            O => \N__18951\,
            I => \N__18948\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__4272\ : Span4Mux_s3_v
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__18942\,
            I => \Lab_UT.dictrl.g1_1Z0Z_0\
        );

    \I__4270\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18936\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__18936\,
            I => \Lab_UT.dictrl.g1_2Z0Z_1\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18930\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__18930\,
            I => \Lab_UT.dictrl.N_102_0\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__18927\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__18924\,
            I => \buart__rx_ser_clk_cascade_\
        );

    \I__4264\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18918\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__18918\,
            I => \N__18915\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__18915\,
            I => \Lab_UT.dictrl.g1_0_0_0\
        );

    \I__4261\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18909\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__18909\,
            I => \N__18906\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__18906\,
            I => \N__18903\
        );

    \I__4258\ : Odrv4
    port map (
            O => \N__18903\,
            I => \Lab_UT.dictrl.N_88_2\
        );

    \I__4257\ : CascadeMux
    port map (
            O => \N__18900\,
            I => \N__18894\
        );

    \I__4256\ : CascadeMux
    port map (
            O => \N__18899\,
            I => \N__18890\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__18898\,
            I => \N__18884\
        );

    \I__4254\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18877\
        );

    \I__4253\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18877\
        );

    \I__4252\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18874\
        );

    \I__4251\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18871\
        );

    \I__4250\ : InMux
    port map (
            O => \N__18889\,
            I => \N__18868\
        );

    \I__4249\ : CascadeMux
    port map (
            O => \N__18888\,
            I => \N__18865\
        );

    \I__4248\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18860\
        );

    \I__4247\ : InMux
    port map (
            O => \N__18884\,
            I => \N__18860\
        );

    \I__4246\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18855\
        );

    \I__4245\ : InMux
    port map (
            O => \N__18882\,
            I => \N__18855\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__18877\,
            I => \N__18845\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18874\,
            I => \N__18845\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__18871\,
            I => \N__18845\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18868\,
            I => \N__18845\
        );

    \I__4240\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18842\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__18860\,
            I => \N__18839\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__18855\,
            I => \N__18836\
        );

    \I__4237\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18833\
        );

    \I__4236\ : Span4Mux_v
    port map (
            O => \N__18845\,
            I => \N__18826\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__18842\,
            I => \N__18826\
        );

    \I__4234\ : Span4Mux_s3_h
    port map (
            O => \N__18839\,
            I => \N__18826\
        );

    \I__4233\ : Span4Mux_v
    port map (
            O => \N__18836\,
            I => \N__18821\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18821\
        );

    \I__4231\ : Span4Mux_h
    port map (
            O => \N__18826\,
            I => \N__18818\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__18821\,
            I => \N__18815\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__18818\,
            I => bu_rx_data_i_4_3
        );

    \I__4228\ : Odrv4
    port map (
            O => \N__18815\,
            I => bu_rx_data_i_4_3
        );

    \I__4227\ : CascadeMux
    port map (
            O => \N__18810\,
            I => \Lab_UT.dictrl.N_95_0_cascade_\
        );

    \I__4226\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18804\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__18804\,
            I => \N__18801\
        );

    \I__4224\ : Odrv12
    port map (
            O => \N__18801\,
            I => \Lab_UT.dictrl.N_103_0\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__18798\,
            I => \N__18795\
        );

    \I__4222\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18792\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__18792\,
            I => \N__18789\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__18789\,
            I => \Lab_UT.dictrl.g1_2_1_0\
        );

    \I__4219\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18783\
        );

    \I__4218\ : LocalMux
    port map (
            O => \N__18783\,
            I => \N__18780\
        );

    \I__4217\ : Odrv4
    port map (
            O => \N__18780\,
            I => \Lab_UT.dictrl.g1_3\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18773\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18770\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__18773\,
            I => \N__18767\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__18770\,
            I => \Lab_UT.dictrl.N_88\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__18767\,
            I => \Lab_UT.dictrl.N_88\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__18762\,
            I => \N__18759\
        );

    \I__4210\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18756\
        );

    \I__4209\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18753\
        );

    \I__4208\ : Odrv12
    port map (
            O => \N__18753\,
            I => \Lab_UT.dictrl.N_95\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18747\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__18747\,
            I => \N__18744\
        );

    \I__4205\ : Odrv4
    port map (
            O => \N__18744\,
            I => \Lab_UT.dictrl.N_103\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18733\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18733\
        );

    \I__4202\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18730\
        );

    \I__4201\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18726\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__18733\,
            I => \N__18721\
        );

    \I__4199\ : LocalMux
    port map (
            O => \N__18730\,
            I => \N__18721\
        );

    \I__4198\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18711\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18708\
        );

    \I__4196\ : Span4Mux_s2_v
    port map (
            O => \N__18721\,
            I => \N__18704\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18720\,
            I => \N__18701\
        );

    \I__4194\ : InMux
    port map (
            O => \N__18719\,
            I => \N__18696\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18696\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18717\,
            I => \N__18688\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18716\,
            I => \N__18688\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18688\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18714\,
            I => \N__18685\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__18711\,
            I => \N__18682\
        );

    \I__4187\ : Span4Mux_s3_v
    port map (
            O => \N__18708\,
            I => \N__18679\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18707\,
            I => \N__18676\
        );

    \I__4185\ : Span4Mux_v
    port map (
            O => \N__18704\,
            I => \N__18673\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18670\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__18696\,
            I => \N__18663\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18660\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__18688\,
            I => \N__18655\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__18685\,
            I => \N__18655\
        );

    \I__4179\ : Span4Mux_s3_v
    port map (
            O => \N__18682\,
            I => \N__18652\
        );

    \I__4178\ : Span4Mux_v
    port map (
            O => \N__18679\,
            I => \N__18647\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__18676\,
            I => \N__18647\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__18673\,
            I => \N__18644\
        );

    \I__4175\ : Span12Mux_s10_v
    port map (
            O => \N__18670\,
            I => \N__18641\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18669\,
            I => \N__18632\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18668\,
            I => \N__18632\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18632\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18666\,
            I => \N__18632\
        );

    \I__4170\ : Span4Mux_v
    port map (
            O => \N__18663\,
            I => \N__18625\
        );

    \I__4169\ : LocalMux
    port map (
            O => \N__18660\,
            I => \N__18625\
        );

    \I__4168\ : Span4Mux_h
    port map (
            O => \N__18655\,
            I => \N__18625\
        );

    \I__4167\ : Span4Mux_v
    port map (
            O => \N__18652\,
            I => \N__18620\
        );

    \I__4166\ : Span4Mux_h
    port map (
            O => \N__18647\,
            I => \N__18620\
        );

    \I__4165\ : Odrv4
    port map (
            O => \N__18644\,
            I => bu_rx_data_3
        );

    \I__4164\ : Odrv12
    port map (
            O => \N__18641\,
            I => bu_rx_data_3
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__18632\,
            I => bu_rx_data_3
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__18625\,
            I => bu_rx_data_3
        );

    \I__4161\ : Odrv4
    port map (
            O => \N__18620\,
            I => bu_rx_data_3
        );

    \I__4160\ : InMux
    port map (
            O => \N__18609\,
            I => \N__18606\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__18606\,
            I => \N__18603\
        );

    \I__4158\ : Odrv12
    port map (
            O => \N__18603\,
            I => \Lab_UT.dictrl.m63_0Z0Z_1\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18600\,
            I => \N__18597\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18597\,
            I => \Lab_UT.dictrl.N_95_0_0_1\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \Lab_UT.dictrl.N_99_0_cascade_\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18588\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__18588\,
            I => \Lab_UT.dictrl.N_96_0_0\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18585\,
            I => \N__18582\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__18582\,
            I => \N__18579\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__18579\,
            I => \Lab_UT.dictrl.g2\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__18576\,
            I => \N__18573\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18573\,
            I => \N__18570\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18570\,
            I => \N__18567\
        );

    \I__4146\ : Span4Mux_h
    port map (
            O => \N__18567\,
            I => \N__18564\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__18564\,
            I => \Lab_UT.dictrl.g0_0_0_a3_5\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18561\,
            I => \N__18558\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__18558\,
            I => \N__18555\
        );

    \I__4142\ : Span4Mux_h
    port map (
            O => \N__18555\,
            I => \N__18552\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__18552\,
            I => \Lab_UT.dictrl.N_98_mux_2\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18545\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18541\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18545\,
            I => \N__18538\
        );

    \I__4137\ : CascadeMux
    port map (
            O => \N__18544\,
            I => \N__18533\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18529\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__18538\,
            I => \N__18526\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18537\,
            I => \N__18521\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18536\,
            I => \N__18521\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18533\,
            I => \N__18516\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18532\,
            I => \N__18516\
        );

    \I__4130\ : Span4Mux_h
    port map (
            O => \N__18529\,
            I => \N__18513\
        );

    \I__4129\ : Span4Mux_v
    port map (
            O => \N__18526\,
            I => \N__18510\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18521\,
            I => \N__18505\
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18505\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__18513\,
            I => bu_rx_data_i_4_5
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__18510\,
            I => bu_rx_data_i_4_5
        );

    \I__4124\ : Odrv12
    port map (
            O => \N__18505\,
            I => bu_rx_data_i_4_5
        );

    \I__4123\ : InMux
    port map (
            O => \N__18498\,
            I => \N__18495\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__18495\,
            I => \N__18492\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__18492\,
            I => \N__18489\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__18489\,
            I => \resetGen.escKeyZ0Z_4\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__18486\,
            I => \resetGen.escKeyZ0Z_5_cascade_\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18468\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18468\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18468\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18480\,
            I => \N__18468\
        );

    \I__4114\ : InMux
    port map (
            O => \N__18479\,
            I => \N__18468\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__4112\ : Span12Mux_s8_h
    port map (
            O => \N__18465\,
            I => \N__18462\
        );

    \I__4111\ : Odrv12
    port map (
            O => \N__18462\,
            I => \resetGen.escKeyZ0\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \Lab_UT.dictrl.N_120_0_cascade_\
        );

    \I__4109\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18444\
        );

    \I__4108\ : InMux
    port map (
            O => \N__18455\,
            I => \N__18444\
        );

    \I__4107\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18444\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18453\,
            I => \N__18444\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18444\,
            I => \Lab_UT.dictrl.N_1302_0\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__18441\,
            I => \N__18437\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__18440\,
            I => \N__18434\
        );

    \I__4102\ : InMux
    port map (
            O => \N__18437\,
            I => \N__18423\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18423\
        );

    \I__4100\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18423\
        );

    \I__4099\ : InMux
    port map (
            O => \N__18432\,
            I => \N__18423\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18423\,
            I => \Lab_UT.dictrl.N_119_0\
        );

    \I__4097\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18416\
        );

    \I__4096\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18413\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18416\,
            I => \N__18410\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18413\,
            I => \N__18405\
        );

    \I__4093\ : Span4Mux_s3_h
    port map (
            O => \N__18410\,
            I => \N__18405\
        );

    \I__4092\ : Odrv4
    port map (
            O => \N__18405\,
            I => \Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18402\,
            I => \N__18398\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18395\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18390\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__18395\,
            I => \N__18390\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__18390\,
            I => \Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18387\,
            I => \N__18384\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18384\,
            I => \N__18381\
        );

    \I__4084\ : Odrv4
    port map (
            O => \N__18381\,
            I => \Lab_UT.dictrl.N_120\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18378\,
            I => \N__18375\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18375\,
            I => \N__18371\
        );

    \I__4081\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18368\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__18371\,
            I => \Lab_UT.dictrl.N_99\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__18368\,
            I => \Lab_UT.dictrl.N_99\
        );

    \I__4078\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18360\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__4076\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__18356\,
            I => \Lab_UT.dictrl.N_96\
        );

    \I__4074\ : LocalMux
    port map (
            O => \N__18353\,
            I => \Lab_UT.dictrl.N_96\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__18348\,
            I => \Lab_UT.dictrl.N_99_cascade_\
        );

    \I__4072\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18342\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18339\
        );

    \I__4070\ : Odrv4
    port map (
            O => \N__18339\,
            I => \Lab_UT.dictrl.N_101\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__18336\,
            I => \Lab_UT.dictrl.N_100_cascade_\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18330\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18330\,
            I => \N__18327\
        );

    \I__4066\ : Odrv4
    port map (
            O => \N__18327\,
            I => \Lab_UT.dictrl.next_state_0_1\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__18324\,
            I => \Lab_UT.dictrl.N_104_cascade_\
        );

    \I__4064\ : CascadeMux
    port map (
            O => \N__18321\,
            I => \Lab_UT.dictrl.N_101_cascade_\
        );

    \I__4063\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18314\
        );

    \I__4062\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18311\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__18314\,
            I => \N__18306\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18306\
        );

    \I__4059\ : Odrv4
    port map (
            O => \N__18306\,
            I => \Lab_UT.dictrl.N_5_0\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__18303\,
            I => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18297\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__18297\,
            I => \N__18294\
        );

    \I__4055\ : Span4Mux_h
    port map (
            O => \N__18294\,
            I => \N__18291\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__18291\,
            I => \Lab_UT.dictrl.state_fast_3\
        );

    \I__4053\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18283\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18276\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18286\,
            I => \N__18276\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18283\,
            I => \N__18273\
        );

    \I__4049\ : InMux
    port map (
            O => \N__18282\,
            I => \N__18268\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18281\,
            I => \N__18268\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__18276\,
            I => \N__18265\
        );

    \I__4046\ : Span4Mux_h
    port map (
            O => \N__18273\,
            I => \N__18262\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__18268\,
            I => \N__18257\
        );

    \I__4044\ : Span4Mux_h
    port map (
            O => \N__18265\,
            I => \N__18257\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__18262\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__18257\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__4041\ : CEMux
    port map (
            O => \N__18252\,
            I => \N__18237\
        );

    \I__4040\ : CEMux
    port map (
            O => \N__18251\,
            I => \N__18237\
        );

    \I__4039\ : CEMux
    port map (
            O => \N__18250\,
            I => \N__18237\
        );

    \I__4038\ : CEMux
    port map (
            O => \N__18249\,
            I => \N__18237\
        );

    \I__4037\ : CEMux
    port map (
            O => \N__18248\,
            I => \N__18237\
        );

    \I__4036\ : GlobalMux
    port map (
            O => \N__18237\,
            I => \N__18234\
        );

    \I__4035\ : gio2CtrlBuf
    port map (
            O => \N__18234\,
            I => bu_rx_data_rdy_0_g
        );

    \I__4034\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18228\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18228\,
            I => \N__18220\
        );

    \I__4032\ : InMux
    port map (
            O => \N__18227\,
            I => \N__18217\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18211\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18208\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18205\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__18223\,
            I => \N__18202\
        );

    \I__4027\ : Span4Mux_s1_v
    port map (
            O => \N__18220\,
            I => \N__18195\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18195\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18192\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18188\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18214\,
            I => \N__18185\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18211\,
            I => \N__18180\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18208\,
            I => \N__18180\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18205\,
            I => \N__18177\
        );

    \I__4019\ : InMux
    port map (
            O => \N__18202\,
            I => \N__18174\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18201\,
            I => \N__18169\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18169\
        );

    \I__4016\ : Span4Mux_v
    port map (
            O => \N__18195\,
            I => \N__18164\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__18192\,
            I => \N__18164\
        );

    \I__4014\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18161\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18188\,
            I => \N__18158\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18185\,
            I => \N__18155\
        );

    \I__4011\ : Span4Mux_v
    port map (
            O => \N__18180\,
            I => \N__18147\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__18177\,
            I => \N__18147\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__18174\,
            I => \N__18147\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__18169\,
            I => \N__18144\
        );

    \I__4007\ : Span4Mux_v
    port map (
            O => \N__18164\,
            I => \N__18141\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__18161\,
            I => \N__18138\
        );

    \I__4005\ : Span12Mux_s11_v
    port map (
            O => \N__18158\,
            I => \N__18132\
        );

    \I__4004\ : Span12Mux_s6_v
    port map (
            O => \N__18155\,
            I => \N__18129\
        );

    \I__4003\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18126\
        );

    \I__4002\ : Span4Mux_v
    port map (
            O => \N__18147\,
            I => \N__18123\
        );

    \I__4001\ : Span4Mux_v
    port map (
            O => \N__18144\,
            I => \N__18116\
        );

    \I__4000\ : Span4Mux_h
    port map (
            O => \N__18141\,
            I => \N__18116\
        );

    \I__3999\ : Span4Mux_h
    port map (
            O => \N__18138\,
            I => \N__18116\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18113\
        );

    \I__3997\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18108\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18108\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__18132\,
            I => bu_rx_data_0
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__18129\,
            I => bu_rx_data_0
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18126\,
            I => bu_rx_data_0
        );

    \I__3992\ : Odrv4
    port map (
            O => \N__18123\,
            I => bu_rx_data_0
        );

    \I__3991\ : Odrv4
    port map (
            O => \N__18116\,
            I => bu_rx_data_0
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18113\,
            I => bu_rx_data_0
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__18108\,
            I => bu_rx_data_0
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18087\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__3985\ : Odrv12
    port map (
            O => \N__18084\,
            I => \Lab_UT.dictrl.g0_9Z0Z_1\
        );

    \I__3984\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18073\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18077\,
            I => \N__18068\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18076\,
            I => \N__18068\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__18073\,
            I => \N__18064\
        );

    \I__3979\ : LocalMux
    port map (
            O => \N__18068\,
            I => \N__18061\
        );

    \I__3978\ : InMux
    port map (
            O => \N__18067\,
            I => \N__18058\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__18064\,
            I => \Lab_UT.dictrl.m25Z0Z_4\
        );

    \I__3976\ : Odrv4
    port map (
            O => \N__18061\,
            I => \Lab_UT.dictrl.m25Z0Z_4\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18058\,
            I => \Lab_UT.dictrl.m25Z0Z_4\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__18051\,
            I => \Lab_UT.dictrl.N_116_mux_1_cascade_\
        );

    \I__3973\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18045\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18045\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__3971\ : InMux
    port map (
            O => \N__18042\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__18036\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18033\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18030\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18027\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__3965\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__18021\
        );

    \I__3964\ : InMux
    port map (
            O => \N__18021\,
            I => \N__18017\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18020\,
            I => \N__18014\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18017\,
            I => \N__18011\
        );

    \I__3961\ : LocalMux
    port map (
            O => \N__18014\,
            I => \N__18006\
        );

    \I__3960\ : Span4Mux_h
    port map (
            O => \N__18011\,
            I => \N__18006\
        );

    \I__3959\ : Odrv4
    port map (
            O => \N__18006\,
            I => \Lab_UT.dictrl.state_i_4_0\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__18003\,
            I => \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17997\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17997\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__17994\,
            I => \N__17990\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17985\
        );

    \I__3953\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17978\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17978\
        );

    \I__3951\ : InMux
    port map (
            O => \N__17988\,
            I => \N__17978\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17985\,
            I => \Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__17978\,
            I => \Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2\
        );

    \I__3948\ : InMux
    port map (
            O => \N__17973\,
            I => \N__17970\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__17967\,
            I => \N__17964\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__17961\,
            I => \Lab_UT.dictrl.dicLdStens_1\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__17958\,
            I => \N__17954\
        );

    \I__3942\ : InMux
    port map (
            O => \N__17957\,
            I => \N__17949\
        );

    \I__3941\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17949\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__17949\,
            I => \N__17944\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17941\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17938\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__17944\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__17941\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17938\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3934\ : CascadeMux
    port map (
            O => \N__17931\,
            I => \Lab_UT.didp.countrce2.q_5_1_cascade_\
        );

    \I__3933\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17922\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17915\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17926\,
            I => \N__17915\
        );

    \I__3930\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17912\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17922\,
            I => \N__17909\
        );

    \I__3928\ : InMux
    port map (
            O => \N__17921\,
            I => \N__17904\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17904\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__17915\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__17912\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3924\ : Odrv12
    port map (
            O => \N__17909\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__17904\,
            I => \Lab_UT.didp.di_Stens_1\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17895\,
            I => \N__17891\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17887\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17883\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17876\
        );

    \I__3918\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17876\
        );

    \I__3917\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17876\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__17883\,
            I => \Lab_UT.LdStens\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__17876\,
            I => \Lab_UT.LdStens\
        );

    \I__3914\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17868\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17868\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3912\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17862\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__17862\,
            I => \Lab_UT.LdStens_i_4\
        );

    \I__3910\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17853\
        );

    \I__3909\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17853\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17853\,
            I => \N__17848\
        );

    \I__3907\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17845\
        );

    \I__3906\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17842\
        );

    \I__3905\ : Odrv4
    port map (
            O => \N__17848\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__17845\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__17842\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__17835\,
            I => \N__17830\
        );

    \I__3901\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17825\
        );

    \I__3900\ : InMux
    port map (
            O => \N__17833\,
            I => \N__17825\
        );

    \I__3899\ : InMux
    port map (
            O => \N__17830\,
            I => \N__17822\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__17825\,
            I => \N__17819\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17816\
        );

    \I__3896\ : Span4Mux_s2_v
    port map (
            O => \N__17819\,
            I => \N__17812\
        );

    \I__3895\ : Span4Mux_s2_v
    port map (
            O => \N__17816\,
            I => \N__17809\
        );

    \I__3894\ : InMux
    port map (
            O => \N__17815\,
            I => \N__17806\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__17812\,
            I => \Lab_UT.LdSones\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__17809\,
            I => \Lab_UT.LdSones\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__17806\,
            I => \Lab_UT.LdSones\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17796\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__17796\,
            I => \N__17787\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17782\
        );

    \I__3887\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17782\
        );

    \I__3886\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17779\
        );

    \I__3885\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17772\
        );

    \I__3884\ : InMux
    port map (
            O => \N__17791\,
            I => \N__17772\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17772\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__17787\,
            I => \N__17767\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__17782\,
            I => \N__17767\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17779\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__17772\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__17767\,
            I => \Lab_UT.didp.di_Sones_0\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17757\,
            I => \N__17754\
        );

    \I__3875\ : Span4Mux_s2_v
    port map (
            O => \N__17754\,
            I => \N__17751\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__17751\,
            I => \Lab_UT.didp.countrce1.q_5_0\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__17748\,
            I => \N__17742\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__17747\,
            I => \N__17739\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17746\,
            I => \N__17732\
        );

    \I__3870\ : InMux
    port map (
            O => \N__17745\,
            I => \N__17732\
        );

    \I__3869\ : InMux
    port map (
            O => \N__17742\,
            I => \N__17732\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17739\,
            I => \N__17729\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17732\,
            I => \N__17726\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17729\,
            I => \N__17723\
        );

    \I__3865\ : Span4Mux_s3_v
    port map (
            O => \N__17726\,
            I => \N__17717\
        );

    \I__3864\ : Span4Mux_s3_h
    port map (
            O => \N__17723\,
            I => \N__17717\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17714\
        );

    \I__3862\ : Odrv4
    port map (
            O => \N__17717\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__17714\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17706\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17706\,
            I => \N__17703\
        );

    \I__3858\ : Span4Mux_s3_v
    port map (
            O => \N__17703\,
            I => \N__17700\
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__17700\,
            I => \Lab_UT.LdSones_i_4\
        );

    \I__3856\ : CascadeMux
    port map (
            O => \N__17697\,
            I => \Lab_UT.didp.countrce2.un13_qPone_cascade_\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__17694\,
            I => \Lab_UT.didp.countrce2.un20_qPone_cascade_\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__17691\,
            I => \Lab_UT.didp.countrce2.q_5_3_cascade_\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__17688\,
            I => \N__17684\
        );

    \I__3852\ : CascadeMux
    port map (
            O => \N__17687\,
            I => \N__17681\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17684\,
            I => \N__17678\
        );

    \I__3850\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17672\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17678\,
            I => \N__17669\
        );

    \I__3848\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17666\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17663\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17660\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17672\,
            I => \N__17657\
        );

    \I__3844\ : Span4Mux_h
    port map (
            O => \N__17669\,
            I => \N__17654\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17666\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__17663\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17660\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3840\ : Odrv12
    port map (
            O => \N__17657\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__17654\,
            I => \Lab_UT.didp.di_Stens_3\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17640\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__17640\,
            I => \Lab_UT.didp.countrce2.q_5_0\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17630\
        );

    \I__3835\ : InMux
    port map (
            O => \N__17636\,
            I => \N__17627\
        );

    \I__3834\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17624\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17634\,
            I => \N__17621\
        );

    \I__3832\ : InMux
    port map (
            O => \N__17633\,
            I => \N__17617\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__17630\,
            I => \N__17610\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__17627\,
            I => \N__17610\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17624\,
            I => \N__17607\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17621\,
            I => \N__17604\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17601\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17597\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17591\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17591\
        );

    \I__3823\ : Span4Mux_s2_v
    port map (
            O => \N__17610\,
            I => \N__17588\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__17607\,
            I => \N__17581\
        );

    \I__3821\ : Span4Mux_s2_v
    port map (
            O => \N__17604\,
            I => \N__17581\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__17601\,
            I => \N__17581\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17600\,
            I => \N__17578\
        );

    \I__3818\ : Span4Mux_h
    port map (
            O => \N__17597\,
            I => \N__17575\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17572\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__17591\,
            I => \N__17567\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__17588\,
            I => \N__17567\
        );

    \I__3814\ : Span4Mux_v
    port map (
            O => \N__17581\,
            I => \N__17558\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17578\,
            I => \N__17558\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__17575\,
            I => \N__17555\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17552\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__17567\,
            I => \N__17549\
        );

    \I__3809\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17540\
        );

    \I__3808\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17540\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17540\
        );

    \I__3806\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17540\
        );

    \I__3805\ : Span4Mux_v
    port map (
            O => \N__17558\,
            I => \N__17537\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__17555\,
            I => bu_rx_data_2
        );

    \I__3803\ : Odrv4
    port map (
            O => \N__17552\,
            I => bu_rx_data_2
        );

    \I__3802\ : Odrv4
    port map (
            O => \N__17549\,
            I => bu_rx_data_2
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__17540\,
            I => bu_rx_data_2
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__17537\,
            I => bu_rx_data_2
        );

    \I__3799\ : InMux
    port map (
            O => \N__17526\,
            I => \N__17523\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__17523\,
            I => \Lab_UT.didp.countrce2.un13_qPone\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__17520\,
            I => \Lab_UT.didp.countrce2.q_5_2_cascade_\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__17517\,
            I => \N__17511\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__17516\,
            I => \N__17507\
        );

    \I__3794\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17504\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17500\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17511\,
            I => \N__17497\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17510\,
            I => \N__17494\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17491\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17504\,
            I => \N__17488\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17485\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17500\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17497\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17494\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17491\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3783\ : Odrv12
    port map (
            O => \N__17488\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17485\,
            I => \Lab_UT.didp.di_Stens_2\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17467\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17464\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17470\,
            I => \N__17457\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17467\,
            I => \N__17452\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__17464\,
            I => \N__17452\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17463\,
            I => \N__17447\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17447\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17442\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17460\,
            I => \N__17442\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17457\,
            I => \N__17437\
        );

    \I__3771\ : Span4Mux_h
    port map (
            O => \N__17452\,
            I => \N__17437\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17447\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17442\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__17437\,
            I => \Lab_UT.didp.di_Stens_0\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17430\,
            I => \N__17424\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17429\,
            I => \N__17421\
        );

    \I__3765\ : CascadeMux
    port map (
            O => \N__17428\,
            I => \N__17417\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__17427\,
            I => \N__17414\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__17424\,
            I => \N__17409\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17421\,
            I => \N__17409\
        );

    \I__3761\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17402\
        );

    \I__3760\ : InMux
    port map (
            O => \N__17417\,
            I => \N__17402\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17402\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__17409\,
            I => \N__17397\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17402\,
            I => \N__17397\
        );

    \I__3756\ : Span4Mux_h
    port map (
            O => \N__17397\,
            I => \N__17394\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__17394\,
            I => \buart__rx_shifter_0_fast_3\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17388\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__17388\,
            I => \N__17384\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17381\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__17384\,
            I => \N__17372\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17381\,
            I => \N__17369\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17362\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17362\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17362\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17377\,
            I => \N__17355\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17376\,
            I => \N__17355\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17355\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__17372\,
            I => bu_rx_data_5_rep1
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__17369\,
            I => bu_rx_data_5_rep1
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__17362\,
            I => bu_rx_data_5_rep1
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__17355\,
            I => bu_rx_data_5_rep1
        );

    \I__3739\ : InMux
    port map (
            O => \N__17346\,
            I => \N__17343\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17343\,
            I => \N__17339\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17342\,
            I => \N__17332\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__17339\,
            I => \N__17329\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17320\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17320\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17336\,
            I => \N__17320\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17335\,
            I => \N__17320\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17332\,
            I => bu_rx_data_4_rep1
        );

    \I__3730\ : Odrv4
    port map (
            O => \N__17329\,
            I => bu_rx_data_4_rep1
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17320\,
            I => bu_rx_data_4_rep1
        );

    \I__3728\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17308\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__17312\,
            I => \N__17303\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17311\,
            I => \N__17300\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__17308\,
            I => \N__17297\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17292\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17306\,
            I => \N__17292\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17289\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__17300\,
            I => \N__17286\
        );

    \I__3720\ : Odrv4
    port map (
            O => \N__17297\,
            I => bu_rx_data_fast_5
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17292\,
            I => bu_rx_data_fast_5
        );

    \I__3718\ : LocalMux
    port map (
            O => \N__17289\,
            I => bu_rx_data_fast_5
        );

    \I__3717\ : Odrv4
    port map (
            O => \N__17286\,
            I => bu_rx_data_fast_5
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__17277\,
            I => \N__17272\
        );

    \I__3715\ : CascadeMux
    port map (
            O => \N__17276\,
            I => \N__17266\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17263\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17256\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17271\,
            I => \N__17256\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17256\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17251\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17251\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17263\,
            I => bu_rx_data_i_4_7_rep1
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__17256\,
            I => bu_rx_data_i_4_7_rep1
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__17251\,
            I => bu_rx_data_i_4_7_rep1
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17244\,
            I => \N__17241\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17241\,
            I => \N__17238\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17238\,
            I => \Lab_UT.dictrl.g0_28_1Z0Z_0\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17235\,
            I => \N__17229\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17226\
        );

    \I__3700\ : InMux
    port map (
            O => \N__17233\,
            I => \N__17223\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17220\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__17229\,
            I => \N__17217\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__17226\,
            I => \N__17210\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17223\,
            I => \N__17210\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17220\,
            I => \N__17210\
        );

    \I__3694\ : Span4Mux_h
    port map (
            O => \N__17217\,
            I => \N__17207\
        );

    \I__3693\ : Odrv4
    port map (
            O => \N__17210\,
            I => bu_rx_data_fast_6
        );

    \I__3692\ : Odrv4
    port map (
            O => \N__17207\,
            I => bu_rx_data_fast_6
        );

    \I__3691\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17199\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__17199\,
            I => \Lab_UT.dictrl.m31_xZ0Z0\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17185\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17185\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17194\,
            I => \N__17185\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17180\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17192\,
            I => \N__17180\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17185\,
            I => \N__17177\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17180\,
            I => \N__17171\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__17177\,
            I => \N__17171\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17176\,
            I => \N__17168\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__17171\,
            I => bu_rx_data_6_rep1
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__17168\,
            I => bu_rx_data_6_rep1
        );

    \I__3678\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17160\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17160\,
            I => \N__17157\
        );

    \I__3676\ : Odrv4
    port map (
            O => \N__17157\,
            I => \Lab_UT.dictrl.g0_43_xZ0\
        );

    \I__3675\ : CascadeMux
    port map (
            O => \N__17154\,
            I => \Lab_UT.dictrl.N_84_cascade_\
        );

    \I__3674\ : InMux
    port map (
            O => \N__17151\,
            I => \N__17148\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__17148\,
            I => \N__17144\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17141\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__17144\,
            I => \N__17138\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__17141\,
            I => \N__17135\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__17138\,
            I => \Lab_UT.dictrl.alarmstate8_2\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__17135\,
            I => \Lab_UT.dictrl.alarmstate8_2\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__17130\,
            I => \N__17127\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17124\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17124\,
            I => \Lab_UT.dictrl.g1_0_0_0_0\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17118\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17118\,
            I => \N__17115\
        );

    \I__3662\ : Odrv4
    port map (
            O => \N__17115\,
            I => \Lab_UT.dictrl.g0_4_a4Z0Z_5\
        );

    \I__3661\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17108\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__17111\,
            I => \N__17105\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17101\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17096\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17104\,
            I => \N__17096\
        );

    \I__3656\ : Sp12to4
    port map (
            O => \N__17101\,
            I => \N__17091\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__17096\,
            I => \N__17091\
        );

    \I__3654\ : Odrv12
    port map (
            O => \N__17091\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__17088\,
            I => \N__17083\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__17087\,
            I => \N__17079\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17075\
        );

    \I__3650\ : InMux
    port map (
            O => \N__17083\,
            I => \N__17068\
        );

    \I__3649\ : InMux
    port map (
            O => \N__17082\,
            I => \N__17068\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17068\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__17078\,
            I => \N__17065\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17060\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17068\,
            I => \N__17060\
        );

    \I__3644\ : InMux
    port map (
            O => \N__17065\,
            I => \N__17057\
        );

    \I__3643\ : Span4Mux_h
    port map (
            O => \N__17060\,
            I => \N__17054\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17057\,
            I => bu_rx_data_i_4_0
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__17054\,
            I => bu_rx_data_i_4_0
        );

    \I__3640\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17046\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__17046\,
            I => \Lab_UT.dictrl.g1_5\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17040\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__17040\,
            I => \Lab_UT.dictrl.g0_5_4\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__17037\,
            I => \N__17031\
        );

    \I__3635\ : CascadeMux
    port map (
            O => \N__17036\,
            I => \N__17027\
        );

    \I__3634\ : CascadeMux
    port map (
            O => \N__17035\,
            I => \N__17022\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__17034\,
            I => \N__17018\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17007\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17030\,
            I => \N__17007\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17007\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17007\
        );

    \I__3628\ : InMux
    port map (
            O => \N__17025\,
            I => \N__17007\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17022\,
            I => \N__16999\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17021\,
            I => \N__16999\
        );

    \I__3625\ : InMux
    port map (
            O => \N__17018\,
            I => \N__16999\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__17007\,
            I => \N__16995\
        );

    \I__3623\ : InMux
    port map (
            O => \N__17006\,
            I => \N__16990\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__16999\,
            I => \N__16987\
        );

    \I__3621\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16984\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__16995\,
            I => \N__16981\
        );

    \I__3619\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16978\
        );

    \I__3618\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16975\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__16990\,
            I => \N__16972\
        );

    \I__3616\ : Span4Mux_v
    port map (
            O => \N__16987\,
            I => \N__16967\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16967\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__16981\,
            I => \Lab_UT.dicLdMones_1\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__16978\,
            I => \Lab_UT.dicLdMones_1\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__16975\,
            I => \Lab_UT.dicLdMones_1\
        );

    \I__3611\ : Odrv4
    port map (
            O => \N__16972\,
            I => \Lab_UT.dicLdMones_1\
        );

    \I__3610\ : Odrv4
    port map (
            O => \N__16967\,
            I => \Lab_UT.dicLdMones_1\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__16956\,
            I => \Lab_UT.dictrl.N_1300_0_cascade_\
        );

    \I__3608\ : InMux
    port map (
            O => \N__16953\,
            I => \N__16950\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16950\,
            I => \Lab_UT.dictrl.g1_2_0\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__16947\,
            I => \Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_\
        );

    \I__3605\ : InMux
    port map (
            O => \N__16944\,
            I => \N__16934\
        );

    \I__3604\ : InMux
    port map (
            O => \N__16943\,
            I => \N__16934\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16934\
        );

    \I__3602\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16931\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__16934\,
            I => \N__16928\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__16931\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3599\ : Odrv4
    port map (
            O => \N__16928\,
            I => \buart__rx_shifter_0_fast_2\
        );

    \I__3598\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16920\
        );

    \I__3597\ : LocalMux
    port map (
            O => \N__16920\,
            I => \Lab_UT.dictrl.g0_5_5\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16914\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__16914\,
            I => \Lab_UT.dictrl.N_7\
        );

    \I__3594\ : InMux
    port map (
            O => \N__16911\,
            I => \N__16908\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__16908\,
            I => \Lab_UT.dictrl.g0_4_a4_4\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16902\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__16902\,
            I => \Lab_UT.dictrl.N_5_2\
        );

    \I__3590\ : InMux
    port map (
            O => \N__16899\,
            I => \N__16896\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16896\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6\
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__16893\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__16890\,
            I => \Lab_UT.dictrl.N_96_1_cascade_\
        );

    \I__3586\ : InMux
    port map (
            O => \N__16887\,
            I => \N__16884\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__16884\,
            I => \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3\
        );

    \I__3584\ : InMux
    port map (
            O => \N__16881\,
            I => \N__16877\
        );

    \I__3583\ : InMux
    port map (
            O => \N__16880\,
            I => \N__16874\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__16877\,
            I => \N__16871\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16874\,
            I => \Lab_UT.dictrl.m36_0\
        );

    \I__3580\ : Odrv4
    port map (
            O => \N__16871\,
            I => \Lab_UT.dictrl.m36_0\
        );

    \I__3579\ : InMux
    port map (
            O => \N__16866\,
            I => \N__16860\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16865\,
            I => \N__16860\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__16860\,
            I => \N__16857\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__16857\,
            I => \Lab_UT.dictrl.g1_5_0\
        );

    \I__3575\ : InMux
    port map (
            O => \N__16854\,
            I => \N__16851\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__16851\,
            I => \Lab_UT.dictrl.m45_1\
        );

    \I__3573\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16843\
        );

    \I__3572\ : InMux
    port map (
            O => \N__16847\,
            I => \N__16838\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16846\,
            I => \N__16838\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__16843\,
            I => \N__16832\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__16838\,
            I => \N__16832\
        );

    \I__3568\ : InMux
    port map (
            O => \N__16837\,
            I => \N__16829\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__16832\,
            I => \N__16824\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__16829\,
            I => \N__16821\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16828\,
            I => \N__16818\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16815\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__16824\,
            I => \Lab_UT.dictrl.m25Z0Z_0\
        );

    \I__3562\ : Odrv4
    port map (
            O => \N__16821\,
            I => \Lab_UT.dictrl.m25Z0Z_0\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__16818\,
            I => \Lab_UT.dictrl.m25Z0Z_0\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__16815\,
            I => \Lab_UT.dictrl.m25Z0Z_0\
        );

    \I__3559\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16803\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16803\,
            I => \N__16800\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__16800\,
            I => \Lab_UT.dictrl.N_6_0\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16794\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__16794\,
            I => \N__16791\
        );

    \I__3554\ : Odrv4
    port map (
            O => \N__16791\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__16788\,
            I => \N__16785\
        );

    \I__3552\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16782\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16779\
        );

    \I__3550\ : Odrv12
    port map (
            O => \N__16779\,
            I => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\
        );

    \I__3549\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16773\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__16773\,
            I => \Lab_UT.dictrl.state_i_4_2\
        );

    \I__3547\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16750\
        );

    \I__3546\ : InMux
    port map (
            O => \N__16769\,
            I => \N__16750\
        );

    \I__3545\ : InMux
    port map (
            O => \N__16768\,
            I => \N__16750\
        );

    \I__3544\ : InMux
    port map (
            O => \N__16767\,
            I => \N__16750\
        );

    \I__3543\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16750\
        );

    \I__3542\ : InMux
    port map (
            O => \N__16765\,
            I => \N__16745\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16764\,
            I => \N__16745\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16763\,
            I => \N__16738\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16738\
        );

    \I__3538\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16738\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__16750\,
            I => \N__16733\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16745\,
            I => \N__16733\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__16738\,
            I => \N__16730\
        );

    \I__3534\ : Span4Mux_h
    port map (
            O => \N__16733\,
            I => \N__16727\
        );

    \I__3533\ : Odrv4
    port map (
            O => \N__16730\,
            I => \Lab_UT.dicLdAMones_2\
        );

    \I__3532\ : Odrv4
    port map (
            O => \N__16727\,
            I => \Lab_UT.dicLdAMones_2\
        );

    \I__3531\ : InMux
    port map (
            O => \N__16722\,
            I => \N__16719\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16719\,
            I => \N__16715\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16712\
        );

    \I__3528\ : Span4Mux_h
    port map (
            O => \N__16715\,
            I => \N__16709\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__16712\,
            I => \Lab_UT.dictrl.N_94_0\
        );

    \I__3526\ : Odrv4
    port map (
            O => \N__16709\,
            I => \Lab_UT.dictrl.N_94_0\
        );

    \I__3525\ : InMux
    port map (
            O => \N__16704\,
            I => \N__16701\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16701\,
            I => \Lab_UT.dictrl.N_2000_0\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16695\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__16695\,
            I => \N__16692\
        );

    \I__3521\ : Odrv4
    port map (
            O => \N__16692\,
            I => \Lab_UT.dictrl.g1\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16689\,
            I => \N__16686\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__16686\,
            I => \Lab_UT.dictrl.g1_3_1\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16679\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16676\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__16679\,
            I => \N__16673\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16676\,
            I => \N__16670\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__16673\,
            I => \N__16667\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__16670\,
            I => \N__16664\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__16667\,
            I => \Lab_UT.dictrl.N_88_0\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__16664\,
            I => \Lab_UT.dictrl.N_88_0\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__16659\,
            I => \Lab_UT.dictrl.g1Z0Z_1_cascade_\
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__16656\,
            I => \Lab_UT.dictrl.i9_mux_0_1_0_cascade_\
        );

    \I__3508\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16650\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__16650\,
            I => \Lab_UT.dictrl.N_94_0_1_0\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__16647\,
            I => \Lab_UT.dictrl.N_2000_0_1_0_cascade_\
        );

    \I__3505\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16641\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16641\,
            I => \N__16638\
        );

    \I__3503\ : Span4Mux_h
    port map (
            O => \N__16638\,
            I => \N__16630\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16627\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16624\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16611\
        );

    \I__3499\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16611\
        );

    \I__3498\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16611\
        );

    \I__3497\ : Span4Mux_v
    port map (
            O => \N__16630\,
            I => \N__16608\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__16627\,
            I => \N__16605\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__16624\,
            I => \N__16602\
        );

    \I__3494\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16595\
        );

    \I__3493\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16595\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16595\
        );

    \I__3491\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16590\
        );

    \I__3490\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16590\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16587\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__16611\,
            I => \N__16582\
        );

    \I__3487\ : Span4Mux_h
    port map (
            O => \N__16608\,
            I => \N__16582\
        );

    \I__3486\ : Odrv12
    port map (
            O => \N__16605\,
            I => \uu0.un4_l_count_0\
        );

    \I__3485\ : Odrv4
    port map (
            O => \N__16602\,
            I => \uu0.un4_l_count_0\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__16595\,
            I => \uu0.un4_l_count_0\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16590\,
            I => \uu0.un4_l_count_0\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16587\,
            I => \uu0.un4_l_count_0\
        );

    \I__3481\ : Odrv4
    port map (
            O => \N__16582\,
            I => \uu0.un4_l_count_0\
        );

    \I__3480\ : IoInMux
    port map (
            O => \N__16569\,
            I => \N__16566\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16563\
        );

    \I__3478\ : IoSpan4Mux
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__3477\ : Span4Mux_s1_h
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__3476\ : Span4Mux_h
    port map (
            O => \N__16557\,
            I => \N__16554\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__16554\,
            I => \uu0.un11_l_count_i\
        );

    \I__3474\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16538\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16538\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16538\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16538\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16547\,
            I => \N__16535\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16532\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16529\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__16532\,
            I => \N__16524\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__16529\,
            I => \N__16524\
        );

    \I__3465\ : Odrv4
    port map (
            O => \N__16524\,
            I => \Lab_UT.dicLdASones_0\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__16521\,
            I => \N__16518\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16518\,
            I => \N__16515\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16515\,
            I => \Lab_UT.dictrl.g3_1\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16512\,
            I => \Lab_UT.dictrl.i9_mux_0_cascade_\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__16509\,
            I => \Lab_UT.dictrl.N_2000_0_cascade_\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \resetGen.un241_ci_cascade_\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__16503\,
            I => \N__16500\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16494\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16494\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__16494\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__16491\,
            I => \resetGen.reset_count_2_0_4_cascade_\
        );

    \I__3453\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16485\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__16485\,
            I => \resetGen.un241_ci\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__16482\,
            I => \N__16475\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16471\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16480\,
            I => \N__16460\
        );

    \I__3448\ : InMux
    port map (
            O => \N__16479\,
            I => \N__16460\
        );

    \I__3447\ : InMux
    port map (
            O => \N__16478\,
            I => \N__16460\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16460\
        );

    \I__3445\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16460\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__16471\,
            I => \N__16457\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16460\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__16457\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__16452\,
            I => \N__16446\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__16451\,
            I => \N__16441\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \N__16437\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16433\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16446\,
            I => \N__16418\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16418\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16418\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16441\,
            I => \N__16418\
        );

    \I__3433\ : InMux
    port map (
            O => \N__16440\,
            I => \N__16418\
        );

    \I__3432\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16418\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16436\,
            I => \N__16418\
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__16433\,
            I => \N__16414\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__16418\,
            I => \N__16411\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__16417\,
            I => \N__16408\
        );

    \I__3427\ : Span4Mux_h
    port map (
            O => \N__16414\,
            I => \N__16404\
        );

    \I__3426\ : Span4Mux_v
    port map (
            O => \N__16411\,
            I => \N__16401\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16398\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16395\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__16404\,
            I => \N__16392\
        );

    \I__3422\ : Odrv4
    port map (
            O => \N__16401\,
            I => \Lab_UT.dicRun_1\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16398\,
            I => \Lab_UT.dicRun_1\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16395\,
            I => \Lab_UT.dicRun_1\
        );

    \I__3419\ : Odrv4
    port map (
            O => \N__16392\,
            I => \Lab_UT.dicRun_1\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16376\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16382\,
            I => \N__16376\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16373\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__16376\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16373\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16368\,
            I => \N__16364\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16359\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16356\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16351\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16351\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__16359\,
            I => \N__16348\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16356\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__16351\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__16348\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16336\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16331\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16331\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16336\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16331\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16323\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16323\,
            I => \resetGen.un252_ci\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16317\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__16317\,
            I => \N__16313\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16310\
        );

    \I__3394\ : Sp12to4
    port map (
            O => \N__16313\,
            I => \N__16307\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__16310\,
            I => \N__16304\
        );

    \I__3392\ : Span12Mux_s9_v
    port map (
            O => \N__16307\,
            I => \N__16301\
        );

    \I__3391\ : Odrv4
    port map (
            O => \N__16304\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__3390\ : Odrv12
    port map (
            O => \N__16301\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16293\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16293\,
            I => \N__16290\
        );

    \I__3387\ : Span4Mux_h
    port map (
            O => \N__16290\,
            I => \N__16287\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__16287\,
            I => \N__16284\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__16284\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__16281\,
            I => \N__16277\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16280\,
            I => \N__16274\
        );

    \I__3382\ : InMux
    port map (
            O => \N__16277\,
            I => \N__16271\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16274\,
            I => \N__16264\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16271\,
            I => \N__16264\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16261\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16258\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__16264\,
            I => \N__16255\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16261\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16258\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__16255\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16245\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__3371\ : Span4Mux_s2_v
    port map (
            O => \N__16242\,
            I => \N__16238\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16235\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__16238\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__16235\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3367\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16225\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16220\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16220\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__16225\,
            I => \Lab_UT.didp.countrce3.ce_12_2_3\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__16220\,
            I => \Lab_UT.didp.countrce3.ce_12_2_3\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16215\,
            I => \N__16210\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__16214\,
            I => \N__16206\
        );

    \I__3360\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16202\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16197\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16209\,
            I => \N__16197\
        );

    \I__3357\ : InMux
    port map (
            O => \N__16206\,
            I => \N__16190\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16205\,
            I => \N__16190\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16190\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__16197\,
            I => \N__16185\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16190\,
            I => \N__16185\
        );

    \I__3352\ : Odrv12
    port map (
            O => \N__16185\,
            I => \Lab_UT.didp.un24_ce_2\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16182\,
            I => \N__16179\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16179\,
            I => \Lab_UT.didp.reset_12_1_3\
        );

    \I__3349\ : InMux
    port map (
            O => \N__16176\,
            I => \N__16172\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16168\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__16172\,
            I => \N__16165\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16160\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16168\,
            I => \N__16154\
        );

    \I__3344\ : Span4Mux_s3_v
    port map (
            O => \N__16165\,
            I => \N__16154\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16149\
        );

    \I__3342\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16149\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__16160\,
            I => \N__16146\
        );

    \I__3340\ : InMux
    port map (
            O => \N__16159\,
            I => \N__16143\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__16154\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16149\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__16146\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16143\,
            I => \Lab_UT.didp.di_Mtens_1\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__16134\,
            I => \Lab_UT.didp.ce_12_3_cascade_\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16125\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__16130\,
            I => \N__16122\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__16129\,
            I => \N__16119\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__16128\,
            I => \N__16115\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__16125\,
            I => \N__16112\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16109\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16106\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16103\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16100\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__16112\,
            I => \N__16093\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__16109\,
            I => \N__16093\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16106\,
            I => \N__16093\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__16103\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__16100\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__16093\,
            I => \Lab_UT.didp.di_Mtens_3\
        );

    \I__3319\ : InMux
    port map (
            O => \N__16086\,
            I => \N__16083\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__16083\,
            I => \N__16077\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16070\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16070\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16070\
        );

    \I__3314\ : Span4Mux_h
    port map (
            O => \N__16077\,
            I => \N__16065\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16070\,
            I => \N__16065\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__16065\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16041\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16041\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16041\
        );

    \I__3308\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16041\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16058\,
            I => \N__16041\
        );

    \I__3306\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16041\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16041\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16038\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__16038\,
            I => \Lab_UT.didp.un18_ce\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16014\
        );

    \I__3301\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16014\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16014\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16014\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16014\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16030\,
            I => \N__16014\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16014\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16014\,
            I => \N__16009\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__16013\,
            I => \N__16004\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16012\,
            I => \N__16001\
        );

    \I__3292\ : Span4Mux_h
    port map (
            O => \N__16009\,
            I => \N__15998\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16008\,
            I => \N__15995\
        );

    \I__3290\ : CascadeMux
    port map (
            O => \N__16007\,
            I => \N__15990\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16004\,
            I => \N__15985\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__16001\,
            I => \N__15982\
        );

    \I__3287\ : Span4Mux_v
    port map (
            O => \N__15998\,
            I => \N__15977\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__15995\,
            I => \N__15977\
        );

    \I__3285\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15972\
        );

    \I__3284\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15972\
        );

    \I__3283\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15969\
        );

    \I__3282\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15964\
        );

    \I__3281\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15964\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__15985\,
            I => \N__15961\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__15982\,
            I => \N__15958\
        );

    \I__3278\ : Span4Mux_v
    port map (
            O => \N__15977\,
            I => \N__15953\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__15972\,
            I => \N__15953\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__15969\,
            I => \N__15948\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__15964\,
            I => \N__15948\
        );

    \I__3274\ : Span4Mux_v
    port map (
            O => \N__15961\,
            I => \N__15945\
        );

    \I__3273\ : Span4Mux_h
    port map (
            O => \N__15958\,
            I => \N__15942\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__15953\,
            I => \N__15939\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__15948\,
            I => \oneSecStrb\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__15945\,
            I => \oneSecStrb\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__15942\,
            I => \oneSecStrb\
        );

    \I__3268\ : Odrv4
    port map (
            O => \N__15939\,
            I => \oneSecStrb\
        );

    \I__3267\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15924\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15924\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__15924\,
            I => \N__15919\
        );

    \I__3264\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15914\
        );

    \I__3263\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15914\
        );

    \I__3262\ : Span4Mux_h
    port map (
            O => \N__15919\,
            I => \N__15909\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15914\,
            I => \N__15909\
        );

    \I__3260\ : Span4Mux_s0_v
    port map (
            O => \N__15909\,
            I => \N__15906\
        );

    \I__3259\ : Odrv4
    port map (
            O => \N__15906\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3258\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15897\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15892\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15889\
        );

    \I__3255\ : InMux
    port map (
            O => \N__15900\,
            I => \N__15886\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__15897\,
            I => \N__15883\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15878\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15878\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15892\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15889\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__15886\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3248\ : Odrv4
    port map (
            O => \N__15883\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__15878\,
            I => \Lab_UT.didp.di_Mones_1\
        );

    \I__3246\ : InMux
    port map (
            O => \N__15867\,
            I => \N__15861\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15866\,
            I => \N__15861\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__15861\,
            I => \N__15854\
        );

    \I__3243\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15851\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15844\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15844\
        );

    \I__3240\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15844\
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__15854\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__15851\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__15844\,
            I => \Lab_UT.didp.di_Mones_0\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__15837\,
            I => \Lab_UT.didp.countrce3.un13_qPone_cascade_\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__15834\,
            I => \Lab_UT.didp.countrce3.q_5_2_cascade_\
        );

    \I__3234\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15828\
        );

    \I__3233\ : LocalMux
    port map (
            O => \N__15828\,
            I => \Lab_UT.didp.countrce3.un13_qPone\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__15825\,
            I => \N__15817\
        );

    \I__3231\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15814\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__15823\,
            I => \N__15811\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15802\
        );

    \I__3228\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15802\
        );

    \I__3227\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15802\
        );

    \I__3226\ : InMux
    port map (
            O => \N__15817\,
            I => \N__15802\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__15814\,
            I => \N__15799\
        );

    \I__3224\ : InMux
    port map (
            O => \N__15811\,
            I => \N__15796\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__15802\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__15799\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__15796\,
            I => \Lab_UT.didp.di_Mones_2\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15783\
        );

    \I__3219\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15780\
        );

    \I__3218\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15777\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__15786\,
            I => \N__15773\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15783\,
            I => \N__15765\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__15780\,
            I => \N__15765\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__15777\,
            I => \N__15765\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15758\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15758\
        );

    \I__3211\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15758\
        );

    \I__3210\ : Span4Mux_h
    port map (
            O => \N__15765\,
            I => \N__15755\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__15758\,
            I => \N__15752\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__15755\,
            I => \N__15749\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__15752\,
            I => \N__15746\
        );

    \I__3206\ : Odrv4
    port map (
            O => \N__15749\,
            I => \Lab_UT.LdMones\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__15746\,
            I => \Lab_UT.LdMones\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__15741\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__15738\,
            I => \Lab_UT.didp.countrce3.q_5_3_cascade_\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15729\
        );

    \I__3201\ : InMux
    port map (
            O => \N__15734\,
            I => \N__15729\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__15729\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15719\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15725\,
            I => \N__15716\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15724\,
            I => \N__15709\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15709\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15709\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__15719\,
            I => \N__15706\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15703\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__15709\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3191\ : Odrv4
    port map (
            O => \N__15706\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__15703\,
            I => \Lab_UT.didp.di_Mones_3\
        );

    \I__3189\ : InMux
    port map (
            O => \N__15696\,
            I => \N__15690\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15690\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__15690\,
            I => \N__15687\
        );

    \I__3186\ : Span4Mux_v
    port map (
            O => \N__15687\,
            I => \N__15684\
        );

    \I__3185\ : Odrv4
    port map (
            O => \N__15684\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15674\
        );

    \I__3183\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15671\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15668\
        );

    \I__3181\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15663\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15663\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15674\,
            I => \N__15658\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__15671\,
            I => \N__15658\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15668\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__15663\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__15658\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15648\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__15648\,
            I => \N__15645\
        );

    \I__3172\ : Odrv12
    port map (
            O => \N__15645\,
            I => \Lab_UT.dictrl.g0_5_2\
        );

    \I__3171\ : CascadeMux
    port map (
            O => \N__15642\,
            I => \N__15637\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__15641\,
            I => \N__15632\
        );

    \I__3169\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15629\
        );

    \I__3168\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15626\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15621\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15621\
        );

    \I__3165\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15618\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15615\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__15626\,
            I => bu_rx_data_i_4_fast_7
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15621\,
            I => bu_rx_data_i_4_fast_7
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__15618\,
            I => bu_rx_data_i_4_fast_7
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__15615\,
            I => bu_rx_data_i_4_fast_7
        );

    \I__3159\ : CEMux
    port map (
            O => \N__15606\,
            I => \N__15579\
        );

    \I__3158\ : CEMux
    port map (
            O => \N__15605\,
            I => \N__15579\
        );

    \I__3157\ : CEMux
    port map (
            O => \N__15604\,
            I => \N__15579\
        );

    \I__3156\ : CEMux
    port map (
            O => \N__15603\,
            I => \N__15579\
        );

    \I__3155\ : CEMux
    port map (
            O => \N__15602\,
            I => \N__15579\
        );

    \I__3154\ : CEMux
    port map (
            O => \N__15601\,
            I => \N__15579\
        );

    \I__3153\ : CEMux
    port map (
            O => \N__15600\,
            I => \N__15579\
        );

    \I__3152\ : CEMux
    port map (
            O => \N__15599\,
            I => \N__15579\
        );

    \I__3151\ : CEMux
    port map (
            O => \N__15598\,
            I => \N__15579\
        );

    \I__3150\ : GlobalMux
    port map (
            O => \N__15579\,
            I => \N__15576\
        );

    \I__3149\ : gio2CtrlBuf
    port map (
            O => \N__15576\,
            I => \buart__rx_sample_g\
        );

    \I__3148\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15569\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__15572\,
            I => \N__15566\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__15569\,
            I => \N__15563\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15560\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__15563\,
            I => \N__15555\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__15560\,
            I => \N__15552\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15559\,
            I => \N__15549\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15558\,
            I => \N__15546\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__15555\,
            I => \N__15543\
        );

    \I__3139\ : Span4Mux_s2_v
    port map (
            O => \N__15552\,
            I => \N__15540\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15549\,
            I => \N__15537\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__15546\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__15543\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3135\ : Odrv4
    port map (
            O => \N__15540\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__15537\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15521\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__15524\,
            I => \N__15518\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15521\,
            I => \N__15513\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15510\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15517\,
            I => \N__15507\
        );

    \I__3127\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15504\
        );

    \I__3126\ : Span4Mux_h
    port map (
            O => \N__15513\,
            I => \N__15501\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15510\,
            I => \N__15498\
        );

    \I__3124\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15495\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15492\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__15501\,
            I => \N__15487\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__15498\,
            I => \N__15487\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15484\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__15492\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__15487\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3117\ : Odrv4
    port map (
            O => \N__15484\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15474\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__15468\,
            I => \Lab_UT.didp.did_alarmMatch_2\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15458\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15464\,
            I => \N__15454\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15463\,
            I => \N__15447\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15447\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15447\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15458\,
            I => \N__15444\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15457\,
            I => \N__15441\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__15454\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15447\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__15444\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__15441\,
            I => \Lab_UT.didp.di_Sones_1\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15425\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15422\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15419\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15416\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15413\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15425\,
            I => \N__15410\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15422\,
            I => \N__15405\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__15419\,
            I => \N__15405\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__15416\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15413\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__15410\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__15405\,
            I => \Lab_UT.didp.di_Sones_3\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__15396\,
            I => \N__15391\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15385\
        );

    \I__3087\ : InMux
    port map (
            O => \N__15394\,
            I => \N__15385\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15391\,
            I => \N__15382\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15390\,
            I => \N__15379\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__15385\,
            I => \N__15372\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15372\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__15379\,
            I => \N__15369\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15378\,
            I => \N__15364\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15364\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__15372\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__15369\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15364\,
            I => \Lab_UT.didp.di_Sones_2\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15354\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__15354\,
            I => \Lab_UT.dictrl.g1_1_1_0\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15351\,
            I => \N__15345\
        );

    \I__3073\ : InMux
    port map (
            O => \N__15350\,
            I => \N__15345\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__15345\,
            I => \N__15340\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15337\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15334\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__15340\,
            I => bu_rx_data_fast_4
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__15337\,
            I => bu_rx_data_fast_4
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__15334\,
            I => bu_rx_data_fast_4
        );

    \I__3066\ : InMux
    port map (
            O => \N__15327\,
            I => \N__15324\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15324\,
            I => \Lab_UT.dictrl.N_98_mux_0\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__15321\,
            I => \Lab_UT.dictrl.g0_3_1_0_cascade_\
        );

    \I__3063\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15315\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__15315\,
            I => \Lab_UT.dictrl.g0_4Z0Z_1\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__15312\,
            I => \N__15307\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15302\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15302\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15299\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__15302\,
            I => \buart__rx_shifter_ret_1_fast\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15299\,
            I => \buart__rx_shifter_ret_1_fast\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \Lab_UT.dictrl.m25_xZ0Z1_cascade_\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \Lab_UT.dictrl.N_116_mux_cascade_\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__15288\,
            I => \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15282\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15282\,
            I => \N__15279\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__15279\,
            I => \Lab_UT.dictrl.g0_0_0_a3_4\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15276\,
            I => \Lab_UT.dictrl.N_98_mux_4_cascade_\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__15273\,
            I => \Lab_UT.dictrl.N_1304_0_0_cascade_\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15267\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15267\,
            I => \N__15264\
        );

    \I__3045\ : Span4Mux_v
    port map (
            O => \N__15264\,
            I => \N__15261\
        );

    \I__3044\ : Odrv4
    port map (
            O => \N__15261\,
            I => \Lab_UT.dictrl.N_88_0_0\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15258\,
            I => \Lab_UT.dictrl.g1_1_1_cascade_\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15252\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__15252\,
            I => \Lab_UT.dictrl.g1_0\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__15249\,
            I => \Lab_UT.dictrl.N_116_mux_0_cascade_\
        );

    \I__3039\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15243\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__15243\,
            I => \Lab_UT.dictrl.N_116_mux_0_0_0\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__15240\,
            I => \Lab_UT.dictrl.N_1304_0_1_0_cascade_\
        );

    \I__3036\ : InMux
    port map (
            O => \N__15237\,
            I => \N__15234\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15234\,
            I => \Lab_UT.dictrl.N_1304_0\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \Lab_UT.didp.countrce4.q_5_0_cascade_\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15228\,
            I => \N__15222\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15219\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__15226\,
            I => \N__15216\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15211\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15222\,
            I => \N__15206\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15219\,
            I => \N__15206\
        );

    \I__3027\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15199\
        );

    \I__3026\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15199\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15199\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15211\,
            I => \N__15196\
        );

    \I__3023\ : Span4Mux_s1_v
    port map (
            O => \N__15206\,
            I => \N__15193\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__15199\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__15196\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__15193\,
            I => \Lab_UT.didp.di_Mtens_0\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__15186\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15180\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15180\,
            I => \Lab_UT.didp.countrce4.un20_qPone\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__15177\,
            I => \Lab_UT.didp.countrce4.q_5_3_cascade_\
        );

    \I__3015\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15166\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15173\,
            I => \N__15163\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15154\
        );

    \I__3012\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15154\
        );

    \I__3011\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15154\
        );

    \I__3010\ : InMux
    port map (
            O => \N__15169\,
            I => \N__15154\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__15166\,
            I => \N__15147\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__15163\,
            I => \N__15147\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15154\,
            I => \N__15147\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__15147\,
            I => \N__15144\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__15144\,
            I => \Lab_UT.LdMtens\
        );

    \I__3004\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15136\
        );

    \I__3003\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15131\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15131\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__15136\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__15131\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15123\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15123\,
            I => \N__15120\
        );

    \I__2997\ : IoSpan4Mux
    port map (
            O => \N__15120\,
            I => \N__15117\
        );

    \I__2996\ : Odrv4
    port map (
            O => \N__15117\,
            I => \Lab_UT.didp.did_alarmMatch_3\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__15114\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_\
        );

    \I__2994\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15108\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15108\,
            I => \N__15105\
        );

    \I__2992\ : Span4Mux_h
    port map (
            O => \N__15105\,
            I => \N__15102\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__15102\,
            I => \Lab_UT.didp.did_alarmMatch_1\
        );

    \I__2990\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15096\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15096\,
            I => \N__15093\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__15093\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_12\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15090\,
            I => \N__15086\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__15089\,
            I => \N__15083\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__15086\,
            I => \N__15080\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15075\
        );

    \I__2983\ : Span12Mux_s6_h
    port map (
            O => \N__15080\,
            I => \N__15072\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15067\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15078\,
            I => \N__15067\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__15075\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2979\ : Odrv12
    port map (
            O => \N__15072\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__15067\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__15060\,
            I => \N__15056\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__15059\,
            I => \N__15052\
        );

    \I__2975\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15039\
        );

    \I__2974\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15039\
        );

    \I__2973\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15039\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15039\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15050\,
            I => \N__15036\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15049\,
            I => \N__15032\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__15048\,
            I => \N__15027\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__15039\,
            I => \N__15018\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15015\
        );

    \I__2966\ : InMux
    port map (
            O => \N__15035\,
            I => \N__15010\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15010\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15031\,
            I => \N__15003\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15003\
        );

    \I__2962\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15003\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15026\,
            I => \N__14990\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15025\,
            I => \N__14990\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15024\,
            I => \N__14990\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15023\,
            I => \N__14990\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15022\,
            I => \N__14990\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15021\,
            I => \N__14990\
        );

    \I__2955\ : Span4Mux_s2_v
    port map (
            O => \N__15018\,
            I => \N__14987\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__15015\,
            I => \Lab_UT.loadalarm_1\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__15010\,
            I => \Lab_UT.loadalarm_1\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15003\,
            I => \Lab_UT.loadalarm_1\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__14990\,
            I => \Lab_UT.loadalarm_1\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__14987\,
            I => \Lab_UT.loadalarm_1\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14970\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14963\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14963\
        );

    \I__2946\ : InMux
    port map (
            O => \N__14973\,
            I => \N__14963\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__14970\,
            I => \N__14955\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14963\,
            I => \N__14955\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__14962\,
            I => \N__14945\
        );

    \I__2942\ : InMux
    port map (
            O => \N__14961\,
            I => \N__14941\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14938\
        );

    \I__2940\ : Span4Mux_s2_v
    port map (
            O => \N__14955\,
            I => \N__14935\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14930\
        );

    \I__2938\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14930\
        );

    \I__2937\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14917\
        );

    \I__2936\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14917\
        );

    \I__2935\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14917\
        );

    \I__2934\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14917\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14917\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14917\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14914\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__14941\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14938\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__14935\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__14930\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__14917\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__14914\,
            I => \Lab_UT.loadalarm_0_0\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__14901\,
            I => \N__14896\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__14900\,
            I => \N__14893\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__14899\,
            I => \N__14890\
        );

    \I__2921\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14876\
        );

    \I__2920\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14876\
        );

    \I__2919\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14876\
        );

    \I__2918\ : InMux
    port map (
            O => \N__14889\,
            I => \N__14876\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14888\,
            I => \N__14876\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__14887\,
            I => \N__14872\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__14876\,
            I => \N__14869\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14875\,
            I => \N__14864\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14872\,
            I => \N__14864\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__14869\,
            I => \N__14861\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__14864\,
            I => \N__14858\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__14861\,
            I => \Lab_UT.min1_3\
        );

    \I__2909\ : Odrv12
    port map (
            O => \N__14858\,
            I => \Lab_UT.min1_3\
        );

    \I__2908\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14850\,
            I => \N__14847\
        );

    \I__2906\ : Span4Mux_s0_v
    port map (
            O => \N__14847\,
            I => \N__14844\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14844\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14838\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__14838\,
            I => \N__14835\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__14835\,
            I => \N__14830\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14826\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14823\
        );

    \I__2899\ : Span4Mux_h
    port map (
            O => \N__14830\,
            I => \N__14820\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14817\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__14826\,
            I => \N__14814\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__14823\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2895\ : Odrv4
    port map (
            O => \N__14820\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14817\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__14814\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__2892\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14802\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__14802\,
            I => \N__14799\
        );

    \I__2890\ : Span4Mux_v
    port map (
            O => \N__14799\,
            I => \N__14795\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14798\,
            I => \N__14790\
        );

    \I__2888\ : Span4Mux_h
    port map (
            O => \N__14795\,
            I => \N__14787\
        );

    \I__2887\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14784\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14781\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__14790\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__14787\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__14784\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__14781\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__14772\,
            I => \N__14767\
        );

    \I__2880\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14760\
        );

    \I__2879\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14757\
        );

    \I__2878\ : InMux
    port map (
            O => \N__14767\,
            I => \N__14754\
        );

    \I__2877\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14745\
        );

    \I__2876\ : InMux
    port map (
            O => \N__14765\,
            I => \N__14745\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14764\,
            I => \N__14745\
        );

    \I__2874\ : InMux
    port map (
            O => \N__14763\,
            I => \N__14745\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__14760\,
            I => \N__14740\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__14757\,
            I => \N__14740\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__14754\,
            I => \Lab_UT.dicRun_2\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__14745\,
            I => \Lab_UT.dicRun_2\
        );

    \I__2869\ : Odrv4
    port map (
            O => \N__14740\,
            I => \Lab_UT.dicRun_2\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__14733\,
            I => \N__14729\
        );

    \I__2867\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14726\
        );

    \I__2866\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14723\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__14726\,
            I => \N__14719\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14716\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14712\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__14719\,
            I => \N__14709\
        );

    \I__2861\ : Span4Mux_h
    port map (
            O => \N__14716\,
            I => \N__14706\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14715\,
            I => \N__14703\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14712\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__14709\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__14706\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__14703\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__14694\,
            I => \N__14691\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14685\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14690\,
            I => \N__14685\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14685\,
            I => \Lab_UT.didp.countrce4.un13_qPone\
        );

    \I__2851\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14678\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__14681\,
            I => \N__14675\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14678\,
            I => \N__14672\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14668\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__14672\,
            I => \N__14665\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \N__14661\
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__14668\,
            I => \N__14656\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__14665\,
            I => \N__14656\
        );

    \I__2843\ : InMux
    port map (
            O => \N__14664\,
            I => \N__14653\
        );

    \I__2842\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14650\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__14656\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14653\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__14650\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2838\ : InMux
    port map (
            O => \N__14643\,
            I => \N__14640\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__14640\,
            I => \N__14637\
        );

    \I__2836\ : Span4Mux_v
    port map (
            O => \N__14637\,
            I => \N__14632\
        );

    \I__2835\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14627\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14627\
        );

    \I__2833\ : Span4Mux_v
    port map (
            O => \N__14632\,
            I => \N__14623\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14627\,
            I => \N__14620\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14617\
        );

    \I__2830\ : Span4Mux_v
    port map (
            O => \N__14623\,
            I => \N__14612\
        );

    \I__2829\ : Span4Mux_s2_v
    port map (
            O => \N__14620\,
            I => \N__14612\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__14617\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__14612\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14604\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14604\,
            I => \N__14600\
        );

    \I__2824\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14597\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__14600\,
            I => \N__14594\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14591\
        );

    \I__2821\ : Span4Mux_v
    port map (
            O => \N__14594\,
            I => \N__14585\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14591\,
            I => \N__14585\
        );

    \I__2819\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14581\
        );

    \I__2818\ : Span4Mux_s2_v
    port map (
            O => \N__14585\,
            I => \N__14578\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14584\,
            I => \N__14575\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__14581\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__14578\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14575\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__2813\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14557\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14557\
        );

    \I__2811\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14546\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14546\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14546\
        );

    \I__2808\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14546\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14546\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14557\,
            I => \N__14543\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14546\,
            I => \Lab_UT.min1_0\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__14543\,
            I => \Lab_UT.min1_0\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14538\,
            I => \N__14527\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14537\,
            I => \N__14527\
        );

    \I__2801\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14516\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14516\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14516\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14533\,
            I => \N__14516\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14532\,
            I => \N__14516\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__14527\,
            I => \N__14513\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14516\,
            I => \Lab_UT.min1_1\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__14513\,
            I => \Lab_UT.min1_1\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__14508\,
            I => \N__14504\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14507\,
            I => \N__14500\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14497\
        );

    \I__2790\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14494\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14500\,
            I => \N__14490\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__14497\,
            I => \N__14487\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__14494\,
            I => \N__14484\
        );

    \I__2786\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14481\
        );

    \I__2785\ : Span12Mux_s5_h
    port map (
            O => \N__14490\,
            I => \N__14478\
        );

    \I__2784\ : Span12Mux_s6_v
    port map (
            O => \N__14487\,
            I => \N__14475\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__14484\,
            I => \N__14472\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__14481\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2781\ : Odrv12
    port map (
            O => \N__14478\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2780\ : Odrv12
    port map (
            O => \N__14475\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2779\ : Odrv4
    port map (
            O => \N__14472\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14463\,
            I => \Lab_UT.didp.countrce1.q_5_1_cascade_\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__14460\,
            I => \N__14456\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__14459\,
            I => \N__14453\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14448\
        );

    \I__2774\ : InMux
    port map (
            O => \N__14453\,
            I => \N__14448\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__14448\,
            I => \Lab_UT.didp.countrce1.un13_qPone\
        );

    \I__2772\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14438\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14444\,
            I => \N__14438\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14435\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__14438\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__14435\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__14430\,
            I => \Lab_UT.didp.un1_dicLdSones_0_cascade_\
        );

    \I__2766\ : InMux
    port map (
            O => \N__14427\,
            I => \N__14424\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__14424\,
            I => \N__14419\
        );

    \I__2764\ : InMux
    port map (
            O => \N__14423\,
            I => \N__14416\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__14422\,
            I => \N__14410\
        );

    \I__2762\ : Span4Mux_s2_v
    port map (
            O => \N__14419\,
            I => \N__14407\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__14416\,
            I => \N__14404\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14395\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14395\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14395\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14395\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__14407\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__2755\ : Odrv12
    port map (
            O => \N__14404\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__14395\,
            I => \Lab_UT.didp.di_Mtens_2\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__14388\,
            I => \N__14384\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__14387\,
            I => \N__14380\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14376\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14383\,
            I => \N__14373\
        );

    \I__2749\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14370\
        );

    \I__2748\ : InMux
    port map (
            O => \N__14379\,
            I => \N__14367\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14364\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__14373\,
            I => \N__14361\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__14370\,
            I => \N__14356\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14367\,
            I => \N__14356\
        );

    \I__2743\ : Span4Mux_s3_v
    port map (
            O => \N__14364\,
            I => \N__14353\
        );

    \I__2742\ : Span4Mux_s3_v
    port map (
            O => \N__14361\,
            I => \N__14350\
        );

    \I__2741\ : Odrv4
    port map (
            O => \N__14356\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__14353\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__14350\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__2738\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14340\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14337\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__14337\,
            I => \N__14334\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__14334\,
            I => \Lab_UT.didp.did_alarmMatch_5\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__14331\,
            I => \Lab_UT.didp.un1_dicLdMones_0_cascade_\
        );

    \I__2733\ : InMux
    port map (
            O => \N__14328\,
            I => \N__14325\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__14325\,
            I => \N__14322\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__14322\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14319\,
            I => \N__14316\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__14316\,
            I => bu_rx_data_i_4_fast_3
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__14313\,
            I => \N__14309\
        );

    \I__2727\ : CascadeMux
    port map (
            O => \N__14312\,
            I => \N__14306\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14309\,
            I => \N__14303\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14306\,
            I => \N__14300\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14303\,
            I => \buart__rx_shifter_ret_5_fast\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14300\,
            I => \buart__rx_shifter_ret_5_fast\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__14295\,
            I => \Lab_UT.dictrl.g1_1Z0Z_4_cascade_\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__14292\,
            I => \N__14289\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14286\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__14286\,
            I => \Lab_UT.dictrl.N_98_mux_1\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14280\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__14280\,
            I => \Lab_UT.dictrl.N_98_mux_0_0\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14277\,
            I => \Lab_UT.dictrl.g0_3_1_cascade_\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__14274\,
            I => \N__14268\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14259\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14272\,
            I => \N__14259\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14271\,
            I => \N__14259\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14259\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__14259\,
            I => bu_rx_data_7
        );

    \I__2709\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14253\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__14253\,
            I => \N__14250\
        );

    \I__2707\ : Odrv12
    port map (
            O => \N__14250\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_6\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__14247\,
            I => \N__14244\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14241\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14238\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__14238\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_7\
        );

    \I__2702\ : CascadeMux
    port map (
            O => \N__14235\,
            I => \Lab_UT.dictrl.N_127_0_0_cascade_\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14226\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14226\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__14226\,
            I => \Lab_UT.dictrl.justentered_0\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__14223\,
            I => \N__14215\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14222\,
            I => \N__14211\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14208\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14197\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14219\,
            I => \N__14197\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14197\
        );

    \I__2692\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14197\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14197\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14211\,
            I => \Lab_UT.shifter_ret_3_RNIK5FS8_0\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__14208\,
            I => \Lab_UT.shifter_ret_3_RNIK5FS8_0\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14197\,
            I => \Lab_UT.shifter_ret_3_RNIK5FS8_0\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14190\,
            I => \N__14181\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14189\,
            I => \N__14178\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14167\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14187\,
            I => \N__14167\
        );

    \I__2683\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14167\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14185\,
            I => \N__14167\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14167\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14181\,
            I => \Lab_UT.shifter_ret_3_RNIQBH29_0\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__14178\,
            I => \Lab_UT.shifter_ret_3_RNIQBH29_0\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14167\,
            I => \Lab_UT.shifter_ret_3_RNIQBH29_0\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14154\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14154\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__14154\,
            I => \Lab_UT.armed\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__14151\,
            I => \Lab_UT.armed_cascade_\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14148\,
            I => \N__14141\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14147\,
            I => \N__14141\
        );

    \I__2671\ : InMux
    port map (
            O => \N__14146\,
            I => \N__14138\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14135\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__14138\,
            I => \N__14132\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__14135\,
            I => \Lab_UT.alarmMatch\
        );

    \I__2667\ : Odrv12
    port map (
            O => \N__14132\,
            I => \Lab_UT.alarmMatch\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14124\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14124\,
            I => \G_203\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14118\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__14118\,
            I => \Lab_UT.dictrl.alarmstate8_2_reti\
        );

    \I__2662\ : CascadeMux
    port map (
            O => \N__14115\,
            I => \Lab_UT.dictrl.alarmstate8_10_3_cascade_\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14109\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14109\,
            I => \N__14105\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14102\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__14105\,
            I => \Lab_UT.dictrl.alarmstate8\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__14102\,
            I => \Lab_UT.dictrl.alarmstate8\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__14097\,
            I => \Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_\
        );

    \I__2655\ : CascadeMux
    port map (
            O => \N__14094\,
            I => \Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_\
        );

    \I__2654\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14088\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14088\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14079\
        );

    \I__2651\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14079\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14079\,
            I => \Lab_UT.dictrl.alarmstate_0_sqmuxa_1\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__14076\,
            I => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14073\,
            I => \N__14070\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__14070\,
            I => \Lab_UT.dictrl.alarmstate_1_0_i_0\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__14067\,
            I => \Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_\
        );

    \I__2645\ : InMux
    port map (
            O => \N__14064\,
            I => \N__14061\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14061\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_0\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__14058\,
            I => \N__14055\
        );

    \I__2642\ : InMux
    port map (
            O => \N__14055\,
            I => \N__14052\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14052\,
            I => \Lab_UT.dictrl.N_127_0_0\
        );

    \I__2640\ : InMux
    port map (
            O => \N__14049\,
            I => \N__14044\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14048\,
            I => \N__14039\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14047\,
            I => \N__14039\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__14044\,
            I => \Lab_UT.trig\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14039\,
            I => \Lab_UT.trig\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14030\
        );

    \I__2634\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14027\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14030\,
            I => \N__14024\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14027\,
            I => \N__14019\
        );

    \I__2631\ : Span4Mux_s2_v
    port map (
            O => \N__14024\,
            I => \N__14016\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14013\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14010\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__14019\,
            I => \N__14005\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__14016\,
            I => \N__14005\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__14013\,
            I => \N__14002\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__14010\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__2624\ : Odrv4
    port map (
            O => \N__14005\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__2623\ : Odrv12
    port map (
            O => \N__14002\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__13995\,
            I => \N__13992\
        );

    \I__2621\ : InMux
    port map (
            O => \N__13992\,
            I => \N__13988\
        );

    \I__2620\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13983\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13988\,
            I => \N__13980\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__13987\,
            I => \N__13977\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__13986\,
            I => \N__13974\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13971\
        );

    \I__2615\ : Span4Mux_s2_v
    port map (
            O => \N__13980\,
            I => \N__13968\
        );

    \I__2614\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13965\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13962\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__13971\,
            I => \N__13957\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__13968\,
            I => \N__13957\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__13965\,
            I => \N__13954\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__13962\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__2608\ : Odrv4
    port map (
            O => \N__13957\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__2607\ : Odrv12
    port map (
            O => \N__13954\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__2606\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13942\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13937\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13937\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__13942\,
            I => \N__13933\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13937\,
            I => \N__13930\
        );

    \I__2601\ : InMux
    port map (
            O => \N__13936\,
            I => \N__13927\
        );

    \I__2600\ : Span4Mux_v
    port map (
            O => \N__13933\,
            I => \N__13922\
        );

    \I__2599\ : Span4Mux_s2_v
    port map (
            O => \N__13930\,
            I => \N__13922\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13927\,
            I => \N__13917\
        );

    \I__2597\ : Span4Mux_v
    port map (
            O => \N__13922\,
            I => \N__13917\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__13917\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__13914\,
            I => \N__13908\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13905\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13902\
        );

    \I__2592\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13899\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13896\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__13905\,
            I => \N__13893\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__13902\,
            I => \N__13888\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__13899\,
            I => \N__13888\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__13896\,
            I => \N__13885\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__13893\,
            I => \N__13882\
        );

    \I__2585\ : Span4Mux_s2_v
    port map (
            O => \N__13888\,
            I => \N__13879\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__13885\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__13882\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__13879\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__13872\,
            I => \N__13867\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \N__13864\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__13870\,
            I => \N__13858\
        );

    \I__2578\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13846\
        );

    \I__2577\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13846\
        );

    \I__2576\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13846\
        );

    \I__2575\ : InMux
    port map (
            O => \N__13862\,
            I => \N__13846\
        );

    \I__2574\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13846\
        );

    \I__2573\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13841\
        );

    \I__2572\ : InMux
    port map (
            O => \N__13857\,
            I => \N__13841\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__13846\,
            I => \N__13838\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__13841\,
            I => \Lab_UT.min1_2\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__13838\,
            I => \Lab_UT.min1_2\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__13830\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2566\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__13824\,
            I => \N__13820\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13806\
        );

    \I__2563\ : Span4Mux_h
    port map (
            O => \N__13820\,
            I => \N__13801\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13798\
        );

    \I__2561\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13791\
        );

    \I__2560\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13791\
        );

    \I__2559\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13791\
        );

    \I__2558\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13784\
        );

    \I__2557\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13784\
        );

    \I__2556\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13784\
        );

    \I__2555\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13775\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13775\
        );

    \I__2553\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13775\
        );

    \I__2552\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13775\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13772\
        );

    \I__2550\ : InMux
    port map (
            O => \N__13805\,
            I => \N__13769\
        );

    \I__2549\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13766\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__13801\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__13798\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__13791\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__13784\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__13775\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2543\ : Odrv12
    port map (
            O => \N__13772\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__13769\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__13766\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__13749\,
            I => \N__13746\
        );

    \I__2539\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13743\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__13743\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13737\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__13737\,
            I => \N__13734\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__13734\,
            I => \N__13731\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__13731\,
            I => \uu2.bitmap_pmux_26_bm_1\
        );

    \I__2533\ : InMux
    port map (
            O => \N__13728\,
            I => \N__13725\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13725\,
            I => \N__13722\
        );

    \I__2531\ : Span4Mux_h
    port map (
            O => \N__13722\,
            I => \N__13717\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13714\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13711\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__13717\,
            I => \N__13693\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__13714\,
            I => \N__13690\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13711\,
            I => \N__13687\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13684\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13677\
        );

    \I__2523\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13677\
        );

    \I__2522\ : InMux
    port map (
            O => \N__13707\,
            I => \N__13677\
        );

    \I__2521\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13668\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13668\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13668\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13668\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13665\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13662\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13657\
        );

    \I__2514\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13657\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13698\,
            I => \N__13650\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13650\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13696\,
            I => \N__13650\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__13693\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2509\ : Odrv12
    port map (
            O => \N__13690\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__13687\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13684\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13677\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13668\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__13665\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13662\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__13657\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__13650\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13626\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__13623\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__13617\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__13611\,
            I => \N__13608\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__13608\,
            I => \uu2.N_217\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__13605\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13602\,
            I => \N__13599\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__13599\,
            I => \N__13596\
        );

    \I__2489\ : Odrv12
    port map (
            O => \N__13596\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_11\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__13593\,
            I => \Lab_UT.didp.countrce4.q_5_2_cascade_\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__13590\,
            I => \N__13584\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13581\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13578\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13587\,
            I => \N__13575\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13572\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__13581\,
            I => \N__13569\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__13578\,
            I => \N__13564\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13575\,
            I => \N__13564\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__13572\,
            I => \N__13559\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__13569\,
            I => \N__13559\
        );

    \I__2477\ : Span4Mux_s2_v
    port map (
            O => \N__13564\,
            I => \N__13556\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__13559\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__13556\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__13551\,
            I => \uu2.o_adder_vbuf_w_addr_displaying_6_cascade_\
        );

    \I__2473\ : CEMux
    port map (
            O => \N__13548\,
            I => \N__13544\
        );

    \I__2472\ : CEMux
    port map (
            O => \N__13547\,
            I => \N__13541\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__13544\,
            I => \N__13538\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__13541\,
            I => \N__13535\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__13538\,
            I => \N__13532\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__13535\,
            I => \N__13529\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__13532\,
            I => \N__13526\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__13529\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__13526\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__2464\ : CascadeMux
    port map (
            O => \N__13521\,
            I => \N__13518\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13515\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13512\
        );

    \I__2461\ : Span4Mux_v
    port map (
            O => \N__13512\,
            I => \N__13509\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__13509\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13503\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13503\,
            I => \N__13499\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__13502\,
            I => \N__13495\
        );

    \I__2456\ : Span4Mux_v
    port map (
            O => \N__13499\,
            I => \N__13490\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13487\
        );

    \I__2454\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13482\
        );

    \I__2453\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13482\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__13493\,
            I => \N__13479\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__13490\,
            I => \N__13468\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__13487\,
            I => \N__13468\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13468\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13461\
        );

    \I__2447\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13461\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13461\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13476\,
            I => \N__13458\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13475\,
            I => \N__13455\
        );

    \I__2443\ : Span4Mux_h
    port map (
            O => \N__13468\,
            I => \N__13452\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__13461\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13458\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13455\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2439\ : Odrv4
    port map (
            O => \N__13452\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__13443\,
            I => \N__13438\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13435\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13432\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13428\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__13435\,
            I => \N__13425\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__13432\,
            I => \N__13421\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__13431\,
            I => \N__13417\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__13428\,
            I => \N__13412\
        );

    \I__2430\ : Span4Mux_h
    port map (
            O => \N__13425\,
            I => \N__13412\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13409\
        );

    \I__2428\ : Span4Mux_h
    port map (
            O => \N__13421\,
            I => \N__13406\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13420\,
            I => \N__13401\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13417\,
            I => \N__13401\
        );

    \I__2425\ : Span4Mux_v
    port map (
            O => \N__13412\,
            I => \N__13398\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13409\,
            I => \uu2.un15_w_data_displaying_6\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__13406\,
            I => \uu2.un15_w_data_displaying_6\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13401\,
            I => \uu2.un15_w_data_displaying_6\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__13398\,
            I => \uu2.un15_w_data_displaying_6\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13386\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__13386\,
            I => \N__13381\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13374\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13371\
        );

    \I__2416\ : Span4Mux_h
    port map (
            O => \N__13381\,
            I => \N__13368\
        );

    \I__2415\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13359\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13379\,
            I => \N__13359\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13378\,
            I => \N__13359\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13359\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__13374\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__13371\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__13368\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__13359\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13350\,
            I => \N__13347\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13347\,
            I => \N__13343\
        );

    \I__2405\ : CascadeMux
    port map (
            O => \N__13346\,
            I => \N__13339\
        );

    \I__2404\ : Span4Mux_v
    port map (
            O => \N__13343\,
            I => \N__13333\
        );

    \I__2403\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13330\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13327\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13324\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13314\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13314\
        );

    \I__2398\ : Span4Mux_h
    port map (
            O => \N__13333\,
            I => \N__13308\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13301\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__13327\,
            I => \N__13301\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__13324\,
            I => \N__13301\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13298\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13295\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13321\,
            I => \N__13292\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13287\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13287\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__13314\,
            I => \N__13284\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13313\,
            I => \N__13277\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13277\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13311\,
            I => \N__13277\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__13308\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__13301\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__13298\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13295\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13292\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__13287\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__13284\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__13277\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2377\ : InMux
    port map (
            O => \N__13260\,
            I => \N__13257\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13254\
        );

    \I__2375\ : Span4Mux_h
    port map (
            O => \N__13254\,
            I => \N__13247\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__13253\,
            I => \N__13243\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__13252\,
            I => \N__13240\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__13251\,
            I => \N__13237\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13234\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__13247\,
            I => \N__13231\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13246\,
            I => \N__13226\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13243\,
            I => \N__13226\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13240\,
            I => \N__13221\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13221\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13234\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__13231\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13226\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__13221\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13209\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__13209\,
            I => \N__13206\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__13206\,
            I => \N__13203\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__13203\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13197\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13197\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__2355\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13191\,
            I => \uu2.bitmap_pmux_25_am_1\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__13182\,
            I => \N__13179\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__13179\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__13176\,
            I => \N__13173\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13165\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13172\,
            I => \N__13162\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13171\,
            I => \N__13156\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13170\,
            I => \N__13152\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13145\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13145\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13140\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13140\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13133\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13133\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13133\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13156\,
            I => \N__13130\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13127\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13152\,
            I => \N__13124\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__13151\,
            I => \N__13121\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13110\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13145\,
            I => \N__13101\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__13140\,
            I => \N__13101\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__13133\,
            I => \N__13101\
        );

    \I__2329\ : Span4Mux_h
    port map (
            O => \N__13130\,
            I => \N__13101\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13127\,
            I => \N__13096\
        );

    \I__2327\ : Span4Mux_s0_v
    port map (
            O => \N__13124\,
            I => \N__13096\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13093\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13088\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13088\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13118\,
            I => \N__13079\
        );

    \I__2322\ : InMux
    port map (
            O => \N__13117\,
            I => \N__13079\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13079\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13079\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13074\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13074\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13110\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__13101\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__13096\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13093\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__13088\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13079\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13074\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2310\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13056\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13053\
        );

    \I__2308\ : Span4Mux_h
    port map (
            O => \N__13053\,
            I => \N__13050\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__13050\,
            I => \uu2.bitmap_RNIV8902Z0Z_66\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__13047\,
            I => \Lab_UT.didp.un2_did_alarmMatch_0_cascade_\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13038\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13038\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13038\,
            I => \N__13030\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13037\,
            I => \N__13019\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13036\,
            I => \N__13019\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13035\,
            I => \N__13019\
        );

    \I__2299\ : InMux
    port map (
            O => \N__13034\,
            I => \N__13019\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13019\
        );

    \I__2297\ : Span4Mux_s2_v
    port map (
            O => \N__13030\,
            I => \N__13016\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__13019\,
            I => \N__13013\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__13016\,
            I => \Lab_UT.sec2_0\
        );

    \I__2294\ : Odrv4
    port map (
            O => \N__13013\,
            I => \Lab_UT.sec2_0\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__13008\,
            I => \Lab_UT.loadalarm_0_0_cascade_\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12987\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12987\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13003\,
            I => \N__12987\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12987\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12987\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12987\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12983\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12980\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__12983\,
            I => \N__12977\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__12980\,
            I => \N__12974\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__12977\,
            I => \Lab_UT.sec1_0\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__12974\,
            I => \Lab_UT.sec1_0\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12966\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__12966\,
            I => \Lab_UT.didp.did_alarmMatch_7\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__12963\,
            I => \N__12957\
        );

    \I__2277\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12950\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12950\
        );

    \I__2275\ : InMux
    port map (
            O => \N__12960\,
            I => \N__12950\
        );

    \I__2274\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12947\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__12950\,
            I => \N__12942\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__12947\,
            I => \N__12942\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__12942\,
            I => \N__12936\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12929\
        );

    \I__2269\ : InMux
    port map (
            O => \N__12940\,
            I => \N__12929\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12929\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__12936\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12929\,
            I => \uu2.un15_w_data_displaying_5\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__12924\,
            I => \N__12921\
        );

    \I__2264\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12915\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12915\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12915\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12909\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__12909\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__12906\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \Lab_UT.didp.countrce1.q_5_3_cascade_\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__12900\,
            I => \Lab_UT.didp.countrce1.q_5_2_cascade_\
        );

    \I__2256\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__12894\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__2254\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__12888\,
            I => \N__12884\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12881\
        );

    \I__2251\ : Span4Mux_s3_v
    port map (
            O => \N__12884\,
            I => \N__12875\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__12881\,
            I => \N__12875\
        );

    \I__2249\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12872\
        );

    \I__2248\ : Span4Mux_v
    port map (
            O => \N__12875\,
            I => \N__12869\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__12872\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__12869\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__2245\ : CascadeMux
    port map (
            O => \N__12864\,
            I => \N__12861\
        );

    \I__2244\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12857\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__12860\,
            I => \N__12854\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__12857\,
            I => \N__12851\
        );

    \I__2241\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12848\
        );

    \I__2240\ : Span4Mux_s3_v
    port map (
            O => \N__12851\,
            I => \N__12843\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__12848\,
            I => \N__12843\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__12843\,
            I => \N__12838\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12842\,
            I => \N__12833\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12841\,
            I => \N__12833\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__12838\,
            I => \N__12830\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__12833\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__12830\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__2232\ : InMux
    port map (
            O => \N__12825\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__2231\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12818\
        );

    \I__2230\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12815\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__12818\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__12815\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__2227\ : InMux
    port map (
            O => \N__12810\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__2226\ : InMux
    port map (
            O => \N__12807\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__2225\ : InMux
    port map (
            O => \N__12804\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12791\
        );

    \I__2223\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12791\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12799\,
            I => \N__12791\
        );

    \I__2221\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12788\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__12791\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__12788\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12783\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__2216\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12771\
        );

    \I__2215\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12771\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__12771\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__12768\,
            I => \N__12765\
        );

    \I__2212\ : InMux
    port map (
            O => \N__12765\,
            I => \N__12759\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12759\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__12759\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__12756\,
            I => \N__12752\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12749\
        );

    \I__2207\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12746\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12749\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__12746\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__12741\,
            I => \Lab_UT.dispString.N_41_cascade_\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12732\,
            I => \Lab_UT.dispString.dOut_RNO_0Z0Z_0\
        );

    \I__2200\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12717\
        );

    \I__2199\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12717\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12717\
        );

    \I__2197\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12717\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__12717\,
            I => \L3_tx_data_0\
        );

    \I__2195\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12709\
        );

    \I__2194\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12704\
        );

    \I__2193\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12704\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__12709\,
            I => \Lab_UT.alarmchar_1\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__12704\,
            I => \Lab_UT.alarmchar_1\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__12699\,
            I => \N__12691\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__12698\,
            I => \N__12688\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12682\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12676\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12676\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12669\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12669\
        );

    \I__2183\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12669\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12659\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12686\,
            I => \N__12659\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12685\,
            I => \N__12659\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12682\,
            I => \N__12656\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12681\,
            I => \N__12653\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12676\,
            I => \N__12648\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12669\,
            I => \N__12648\
        );

    \I__2175\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12641\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12641\
        );

    \I__2173\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12641\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__12659\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__12656\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12653\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2169\ : Odrv4
    port map (
            O => \N__12648\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__12641\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12630\,
            I => \Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__12624\,
            I => \Lab_UT.dispString.dOut_RNO_0Z0Z_2\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12615\
        );

    \I__2163\ : InMux
    port map (
            O => \N__12620\,
            I => \N__12608\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12608\
        );

    \I__2161\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12608\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12615\,
            I => \L3_tx_data_2\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12608\,
            I => \L3_tx_data_2\
        );

    \I__2158\ : InMux
    port map (
            O => \N__12603\,
            I => \N__12591\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12602\,
            I => \N__12591\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12586\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12586\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12579\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12579\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12579\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12576\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__12591\,
            I => \N__12561\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__12586\,
            I => \N__12561\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12579\,
            I => \N__12561\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12576\,
            I => \N__12558\
        );

    \I__2146\ : InMux
    port map (
            O => \N__12575\,
            I => \N__12549\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12574\,
            I => \N__12549\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12549\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12549\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12571\,
            I => \N__12540\
        );

    \I__2141\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12540\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12540\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12568\,
            I => \N__12540\
        );

    \I__2138\ : Odrv4
    port map (
            O => \N__12561\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__12558\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__12549\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__12540\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12528\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12528\,
            I => \Lab_UT.dispString.N_32\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__12525\,
            I => \N__12514\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \N__12508\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__12523\,
            I => \N__12499\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__12522\,
            I => \N__12496\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__12521\,
            I => \N__12493\
        );

    \I__2127\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12485\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12519\,
            I => \N__12485\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12518\,
            I => \N__12485\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__12517\,
            I => \N__12482\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12514\,
            I => \N__12471\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12471\
        );

    \I__2121\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12471\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12471\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12471\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__12507\,
            I => \N__12468\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__12506\,
            I => \N__12465\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12505\,
            I => \N__12462\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__12504\,
            I => \N__12459\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12456\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12449\
        );

    \I__2112\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12449\
        );

    \I__2111\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12449\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12446\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__12492\,
            I => \N__12443\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12485\,
            I => \N__12438\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12435\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__12471\,
            I => \N__12432\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12423\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12465\,
            I => \N__12423\
        );

    \I__2103\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12423\
        );

    \I__2102\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12423\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12456\,
            I => \N__12420\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12417\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12414\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12407\
        );

    \I__2097\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12407\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12441\,
            I => \N__12407\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__12438\,
            I => \N__12400\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__12435\,
            I => \N__12400\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__12432\,
            I => \N__12400\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__12423\,
            I => \N__12395\
        );

    \I__2091\ : Span4Mux_s3_h
    port map (
            O => \N__12420\,
            I => \N__12395\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__12417\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2089\ : Odrv12
    port map (
            O => \N__12414\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__12407\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__12400\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__12395\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12381\,
            I => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\
        );

    \I__2083\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12373\
        );

    \I__2082\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12368\
        );

    \I__2081\ : InMux
    port map (
            O => \N__12376\,
            I => \N__12368\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__12373\,
            I => \N__12365\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__12368\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__12365\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12357\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__12357\,
            I => \N__12353\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__12356\,
            I => \N__12349\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__12353\,
            I => \N__12345\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12342\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12337\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12337\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__12345\,
            I => \uu2.N_115\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__12342\,
            I => \uu2.N_115\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__12337\,
            I => \uu2.N_115\
        );

    \I__2067\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12321\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12321\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12321\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12321\,
            I => \N__12312\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12303\
        );

    \I__2062\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12303\
        );

    \I__2061\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12303\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12303\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12300\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12297\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__12312\,
            I => \N__12292\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12292\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12300\,
            I => \uu2.N_144\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12297\,
            I => \uu2.N_144\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__12292\,
            I => \uu2.N_144\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12277\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12284\,
            I => \N__12272\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12283\,
            I => \N__12272\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12269\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12266\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__12280\,
            I => \N__12263\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12277\,
            I => \N__12254\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12254\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12269\,
            I => \N__12254\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12266\,
            I => \N__12254\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12251\
        );

    \I__2041\ : Span4Mux_v
    port map (
            O => \N__12254\,
            I => \N__12248\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12251\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2039\ : Odrv4
    port map (
            O => \N__12248\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2038\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12240\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__12240\,
            I => \N__12235\
        );

    \I__2036\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12231\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12228\
        );

    \I__2034\ : Span4Mux_h
    port map (
            O => \N__12235\,
            I => \N__12225\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12222\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12231\,
            I => \o_One_Sec_Pulse\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12228\,
            I => \o_One_Sec_Pulse\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__12225\,
            I => \o_One_Sec_Pulse\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__12222\,
            I => \o_One_Sec_Pulse\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12210\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12203\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12200\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12203\,
            I => \N__12193\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12200\,
            I => \N__12193\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12190\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12198\,
            I => \N__12187\
        );

    \I__2020\ : Span12Mux_s11_h
    port map (
            O => \N__12193\,
            I => \N__12184\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12190\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12187\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2017\ : Odrv12
    port map (
            O => \N__12184\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2016\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12174\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__12174\,
            I => \N__12171\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__12171\,
            I => \N__12167\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12164\
        );

    \I__2012\ : Span4Mux_h
    port map (
            O => \N__12167\,
            I => \N__12161\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__12164\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__12161\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12156\,
            I => \N__12153\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__12153\,
            I => \N__12150\
        );

    \I__2007\ : Span4Mux_v
    port map (
            O => \N__12150\,
            I => \N__12147\
        );

    \I__2006\ : Span4Mux_h
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__12144\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12138\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12138\,
            I => \Lab_UT.dispString.dOutP_1_iv_0_4\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__12135\,
            I => \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\
        );

    \I__2001\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12129\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12129\,
            I => \N__12125\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__12128\,
            I => \N__12120\
        );

    \I__1998\ : Span4Mux_h
    port map (
            O => \N__12125\,
            I => \N__12116\
        );

    \I__1997\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12107\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12107\
        );

    \I__1995\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12107\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12107\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__12116\,
            I => \L3_tx_data_1\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__12107\,
            I => \L3_tx_data_1\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12099\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_5\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12092\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12089\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12086\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__12089\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__1985\ : Odrv12
    port map (
            O => \N__12086\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12078\,
            I => \N__12075\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__12075\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__12072\,
            I => \uu2.N_383_cascade_\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12069\,
            I => \N__12066\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__12063\,
            I => \uu2.N_215\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12057\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__12054\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__1971\ : Odrv12
    port map (
            O => \N__12042\,
            I => \uu2.bitmap_RNIS4UH1Z0Z_314\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12036\,
            I => \uu2.N_397\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12030\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12030\,
            I => \uu2.bitmap_pmux_sn_N_15\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__12027\,
            I => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\
        );

    \I__1965\ : InMux
    port map (
            O => \N__12024\,
            I => \N__12021\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__12021\,
            I => \uu2.bitmap_RNIELSJ2Z0Z_111\
        );

    \I__1963\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12014\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12007\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__12014\,
            I => \N__12004\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__12013\,
            I => \N__12001\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__12012\,
            I => \N__11993\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__12011\,
            I => \N__11989\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__12010\,
            I => \N__11983\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__12007\,
            I => \N__11980\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__12004\,
            I => \N__11977\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12001\,
            I => \N__11968\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11968\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11968\
        );

    \I__1951\ : InMux
    port map (
            O => \N__11998\,
            I => \N__11968\
        );

    \I__1950\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11959\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11959\
        );

    \I__1948\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11959\
        );

    \I__1947\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11959\
        );

    \I__1946\ : InMux
    port map (
            O => \N__11989\,
            I => \N__11954\
        );

    \I__1945\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11954\
        );

    \I__1944\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11951\
        );

    \I__1943\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11946\
        );

    \I__1942\ : InMux
    port map (
            O => \N__11983\,
            I => \N__11946\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__11980\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__11977\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__11968\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__11959\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__11954\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11951\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11946\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__11931\,
            I => \N__11926\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__11930\,
            I => \N__11921\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11917\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11914\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11905\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11905\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11905\
        );

    \I__1927\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11905\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__11917\,
            I => \N__11902\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11914\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__11905\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__11902\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__1922\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11890\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__11894\,
            I => \N__11883\
        );

    \I__1920\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11878\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__11890\,
            I => \N__11875\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11870\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11870\
        );

    \I__1916\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11861\
        );

    \I__1915\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11861\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11861\
        );

    \I__1913\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11861\
        );

    \I__1912\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11856\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11853\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__11875\,
            I => \N__11850\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__11870\,
            I => \N__11847\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__11861\,
            I => \N__11844\
        );

    \I__1907\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11839\
        );

    \I__1906\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11839\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__11856\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1904\ : Odrv12
    port map (
            O => \N__11853\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__11850\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__11847\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__11844\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__11839\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__1899\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11821\
        );

    \I__1898\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11818\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__11824\,
            I => \N__11815\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11808\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__11818\,
            I => \N__11805\
        );

    \I__1894\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11802\
        );

    \I__1893\ : InMux
    port map (
            O => \N__11814\,
            I => \N__11793\
        );

    \I__1892\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11793\
        );

    \I__1891\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11793\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11793\
        );

    \I__1889\ : Span4Mux_h
    port map (
            O => \N__11808\,
            I => \N__11788\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__11805\,
            I => \N__11788\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11802\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__11793\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__11788\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11776\
        );

    \I__1883\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \N__11772\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11769\
        );

    \I__1881\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11765\
        );

    \I__1880\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11758\
        );

    \I__1879\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11758\
        );

    \I__1878\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11758\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__11768\,
            I => \N__11755\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__11765\,
            I => \N__11749\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__11758\,
            I => \N__11749\
        );

    \I__1874\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11746\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11743\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__11749\,
            I => \N__11740\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__11746\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11743\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__11740\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__11733\,
            I => \N__11729\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11726\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11723\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11726\,
            I => \uu2.un33_w_data_displaying\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11723\,
            I => \uu2.un33_w_data_displaying\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11714\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__11717\,
            I => \N__11701\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__11714\,
            I => \N__11696\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11693\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11690\
        );

    \I__1858\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11685\
        );

    \I__1857\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11685\
        );

    \I__1856\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11680\
        );

    \I__1855\ : InMux
    port map (
            O => \N__11708\,
            I => \N__11680\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11707\,
            I => \N__11675\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11675\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11670\
        );

    \I__1851\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11670\
        );

    \I__1850\ : InMux
    port map (
            O => \N__11701\,
            I => \N__11667\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11662\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11662\
        );

    \I__1847\ : Span4Mux_h
    port map (
            O => \N__11696\,
            I => \N__11653\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11693\,
            I => \N__11653\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11690\,
            I => \N__11653\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11685\,
            I => \N__11653\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11680\,
            I => \N__11650\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__11675\,
            I => \N__11645\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__11670\,
            I => \N__11645\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__11667\,
            I => \N__11640\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__11662\,
            I => \N__11640\
        );

    \I__1838\ : Span4Mux_v
    port map (
            O => \N__11653\,
            I => \N__11635\
        );

    \I__1837\ : Span4Mux_v
    port map (
            O => \N__11650\,
            I => \N__11635\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__11645\,
            I => \N__11632\
        );

    \I__1835\ : Odrv12
    port map (
            O => \N__11640\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__11635\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__11632\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__11625\,
            I => \uu2.un21_w_addr_displaying_i_cascade_\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11619\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11619\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11613\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11613\,
            I => \N__11610\
        );

    \I__1827\ : Odrv12
    port map (
            O => \N__11610\,
            I => \uu2.bitmap_pmux_sn_N_65\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__11607\,
            I => \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__11604\,
            I => \N__11600\
        );

    \I__1824\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11594\
        );

    \I__1823\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11594\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11591\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__11594\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__11591\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1819\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11583\,
            I => \uu2.bitmap_pmux_sn_i7_mux_0\
        );

    \I__1817\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11577\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11572\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11567\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11567\
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__11572\,
            I => \uu2.un15_w_data_displaying_2\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__11567\,
            I => \uu2.un15_w_data_displaying_2\
        );

    \I__1811\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11559\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11559\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__11556\,
            I => \N__11553\
        );

    \I__1808\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11550\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__11550\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__11547\,
            I => \uu2.un437_ci_0_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11539\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__11543\,
            I => \N__11536\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__11542\,
            I => \N__11533\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11530\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11525\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11525\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__11530\,
            I => \N__11522\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11525\,
            I => \N__11519\
        );

    \I__1797\ : Odrv4
    port map (
            O => \N__11522\,
            I => \L3_tx_data_6\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__11519\,
            I => \L3_tx_data_6\
        );

    \I__1795\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11511\,
            I => \N__11508\
        );

    \I__1793\ : Span4Mux_h
    port map (
            O => \N__11508\,
            I => \N__11505\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__11505\,
            I => \uu2.mem0.w_data_6\
        );

    \I__1791\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11499\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__11499\,
            I => \uu2.un31_w_data_displaying_2\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__11496\,
            I => \N__11493\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11490\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11490\,
            I => \N__11487\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__11487\,
            I => \N__11484\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__11484\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11478\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11478\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__1781\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11469\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__11469\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__11466\,
            I => \uu2.bitmap_pmux_24_i_m2_bm_1_cascade_\
        );

    \I__1778\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11460\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__11460\,
            I => \uu2.bitmap_RNI1UT12Z0Z_75\
        );

    \I__1776\ : InMux
    port map (
            O => \N__11457\,
            I => \N__11454\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__11454\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11451\,
            I => \N__11448\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__11448\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11442\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__11442\,
            I => \N__11439\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__11439\,
            I => \N__11430\
        );

    \I__1769\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11417\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11417\
        );

    \I__1767\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11417\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11417\
        );

    \I__1765\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11417\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11417\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__11430\,
            I => \Lab_UT.min2_2\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__11417\,
            I => \Lab_UT.min2_2\
        );

    \I__1761\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11409\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11403\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__11408\,
            I => \N__11399\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__11407\,
            I => \N__11396\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__11406\,
            I => \N__11393\
        );

    \I__1756\ : Sp12to4
    port map (
            O => \N__11403\,
            I => \N__11388\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11375\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11375\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11375\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11375\
        );

    \I__1751\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11375\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11375\
        );

    \I__1749\ : Odrv12
    port map (
            O => \N__11388\,
            I => \Lab_UT.min2_1\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__11375\,
            I => \Lab_UT.min2_1\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__11370\,
            I => \N__11367\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11364\,
            I => \N__11358\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11363\,
            I => \N__11355\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11349\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__11361\,
            I => \N__11346\
        );

    \I__1741\ : Span4Mux_v
    port map (
            O => \N__11358\,
            I => \N__11343\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11355\,
            I => \N__11330\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11330\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11330\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11352\,
            I => \N__11330\
        );

    \I__1736\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11330\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11330\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__11343\,
            I => \Lab_UT.min2_3\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__11330\,
            I => \Lab_UT.min2_3\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11322\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__11322\,
            I => \N__11319\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__11319\,
            I => \N__11310\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11297\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11297\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11297\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11297\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11297\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11313\,
            I => \N__11297\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__11310\,
            I => \Lab_UT.min2_0\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__11297\,
            I => \Lab_UT.min2_0\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11292\,
            I => \N__11285\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11291\,
            I => \N__11282\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__11290\,
            I => \N__11278\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__11289\,
            I => \N__11274\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11269\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11269\
        );

    \I__1715\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11258\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11258\
        );

    \I__1713\ : InMux
    port map (
            O => \N__11278\,
            I => \N__11258\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11258\
        );

    \I__1711\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11258\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__11269\,
            I => \Lab_UT.sec2_3\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__11258\,
            I => \Lab_UT.sec2_3\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__11253\,
            I => \N__11248\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \N__11244\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11230\
        );

    \I__1705\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11230\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11230\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11230\
        );

    \I__1702\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11230\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11225\
        );

    \I__1700\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11225\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11230\,
            I => \N__11222\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__11225\,
            I => \Lab_UT.sec2_2\
        );

    \I__1697\ : Odrv4
    port map (
            O => \N__11222\,
            I => \Lab_UT.sec2_2\
        );

    \I__1696\ : CascadeMux
    port map (
            O => \N__11217\,
            I => \N__11209\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11197\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11197\
        );

    \I__1693\ : InMux
    port map (
            O => \N__11214\,
            I => \N__11197\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11213\,
            I => \N__11197\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11212\,
            I => \N__11197\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11209\,
            I => \N__11192\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11208\,
            I => \N__11192\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11197\,
            I => \N__11189\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11192\,
            I => \Lab_UT.sec2_1\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__11189\,
            I => \Lab_UT.sec2_1\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11184\,
            I => \N__11181\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__11181\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__11175\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__11172\,
            I => \uu2.N_216_cascade_\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11151\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11151\
        );

    \I__1678\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11151\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11151\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11151\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11151\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__11151\,
            I => \N__11148\
        );

    \I__1673\ : IoSpan4Mux
    port map (
            O => \N__11148\,
            I => \N__11144\
        );

    \I__1672\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11141\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__11144\,
            I => \Lab_UT.sec1_1\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__11141\,
            I => \Lab_UT.sec1_1\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__11136\,
            I => \N__11130\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \N__11127\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__11134\,
            I => \N__11124\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__11133\,
            I => \N__11121\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11105\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11127\,
            I => \N__11105\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11124\,
            I => \N__11105\
        );

    \I__1662\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11105\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11105\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11105\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__11118\,
            I => \N__11102\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__11105\,
            I => \N__11099\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11096\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__11099\,
            I => \Lab_UT.sec1_2\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11096\,
            I => \Lab_UT.sec1_2\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__11091\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__11088\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__11085\,
            I => \buart.Z_tx.un1_bitcount_c2_cascade_\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11077\
        );

    \I__1650\ : InMux
    port map (
            O => \N__11081\,
            I => \N__11072\
        );

    \I__1649\ : InMux
    port map (
            O => \N__11080\,
            I => \N__11072\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__11077\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11072\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11067\,
            I => \N__11061\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11058\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11051\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11051\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11046\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__11046\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11041\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11041\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11051\,
            I => \N__11036\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__11046\,
            I => \N__11036\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11041\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1635\ : Odrv4
    port map (
            O => \N__11036\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__11031\,
            I => \N__11028\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11019\
        );

    \I__1632\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11019\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11019\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__11016\,
            I => \N__11004\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11015\,
            I => \N__10993\
        );

    \I__1627\ : InMux
    port map (
            O => \N__11014\,
            I => \N__10993\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11013\,
            I => \N__10993\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11012\,
            I => \N__10993\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11011\,
            I => \N__10993\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10990\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10985\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10985\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__11007\,
            I => \N__10978\
        );

    \I__1619\ : Span4Mux_v
    port map (
            O => \N__11004\,
            I => \N__10975\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__10993\,
            I => \N__10968\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10968\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10968\
        );

    \I__1615\ : InMux
    port map (
            O => \N__10984\,
            I => \N__10959\
        );

    \I__1614\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10959\
        );

    \I__1613\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10959\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10959\
        );

    \I__1611\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10956\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__10975\,
            I => \N__10953\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__10968\,
            I => \N__10948\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10948\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__10956\,
            I => vbuf_tx_data_rdy
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__10953\,
            I => vbuf_tx_data_rdy
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__10948\,
            I => vbuf_tx_data_rdy
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__10941\,
            I => \N__10937\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10940\,
            I => \N__10929\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10929\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10924\
        );

    \I__1600\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10924\
        );

    \I__1599\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10921\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__10929\,
            I => \N__10916\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__10924\,
            I => \N__10916\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__10921\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__10916\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1594\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10899\
        );

    \I__1593\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10899\
        );

    \I__1592\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10899\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10899\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__10899\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10893\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__10893\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__10890\,
            I => \N__10887\
        );

    \I__1586\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10884\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__10884\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10878\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__10878\,
            I => \uu2.bitmap_pmux_25_bm_1\
        );

    \I__1582\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10872\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__10872\,
            I => \Lab_UT.dispString.N_50\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__10869\,
            I => \Lab_UT.dispString.N_28_cascade_\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10866\,
            I => \N__10863\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__10863\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_3\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__10860\,
            I => \buart.Z_tx.un1_bitcount_c3_cascade_\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10853\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10850\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10853\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10850\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__10845\,
            I => \N__10841\
        );

    \I__1571\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10838\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10834\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__10838\,
            I => \N__10831\
        );

    \I__1568\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10828\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10834\,
            I => \N__10825\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__10831\,
            I => \uu2.N_361\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__10828\,
            I => \uu2.N_361\
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__10825\,
            I => \uu2.N_361\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__10818\,
            I => \uu2.mem0.w_data_0_a2_0_4_cascade_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10812\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__10812\,
            I => \N__10809\
        );

    \I__1560\ : Span4Mux_s3_h
    port map (
            O => \N__10809\,
            I => \N__10806\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__10806\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1558\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10798\
        );

    \I__1557\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10795\
        );

    \I__1556\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10792\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__10798\,
            I => \N__10789\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10784\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10784\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__10789\,
            I => \L3_tx_data_5\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__10784\,
            I => \L3_tx_data_5\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10779\,
            I => \N__10773\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10773\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10770\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__10770\,
            I => \L3_tx_data_4\
        );

    \I__1546\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10755\
        );

    \I__1545\ : InMux
    port map (
            O => \N__10766\,
            I => \N__10755\
        );

    \I__1544\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10755\
        );

    \I__1543\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10755\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__10755\,
            I => \uu2.N_109\
        );

    \I__1541\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10746\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__10746\,
            I => \uu2.N_111\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__10743\,
            I => \uu2.N_109_cascade_\
        );

    \I__1537\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10730\
        );

    \I__1536\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10730\
        );

    \I__1535\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10727\
        );

    \I__1534\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10720\
        );

    \I__1533\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10720\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10720\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10717\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__10727\,
            I => \L3_tx_data_rdy\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__10720\,
            I => \L3_tx_data_rdy\
        );

    \I__1528\ : Odrv4
    port map (
            O => \N__10717\,
            I => \L3_tx_data_rdy\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__10710\,
            I => \N__10705\
        );

    \I__1526\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10701\
        );

    \I__1525\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10694\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10694\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10704\,
            I => \N__10694\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10691\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__10694\,
            I => \N__10688\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__10691\,
            I => \N__10685\
        );

    \I__1519\ : Odrv4
    port map (
            O => \N__10688\,
            I => \Lab_UT.dispString.N_61\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__10685\,
            I => \Lab_UT.dispString.N_61\
        );

    \I__1517\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10674\
        );

    \I__1515\ : Span4Mux_h
    port map (
            O => \N__10674\,
            I => \N__10671\
        );

    \I__1514\ : Odrv4
    port map (
            O => \N__10671\,
            I => \Lab_UT.dispString.un46_dOutP_i_m_3\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__10668\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_3_cascade_\
        );

    \I__1512\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__10662\,
            I => \Lab_UT.dispString.dOutP_6\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10656\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10653\
        );

    \I__1508\ : Span12Mux_s4_v
    port map (
            O => \N__10653\,
            I => \N__10648\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10643\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10643\
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__10648\,
            I => \L3_tx_data_3\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__10643\,
            I => \L3_tx_data_3\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__10638\,
            I => \uu2.N_111_cascade_\
        );

    \I__1502\ : SRMux
    port map (
            O => \N__10635\,
            I => \N__10631\
        );

    \I__1501\ : CEMux
    port map (
            O => \N__10634\,
            I => \N__10628\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10631\,
            I => \N__10625\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__10628\,
            I => \N__10622\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__10625\,
            I => \N__10617\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__10622\,
            I => \N__10617\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__10617\,
            I => \N__10614\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__10614\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__10611\,
            I => \uu2.mem0.w_data_i_a2_1_0_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__10605\,
            I => \N__10602\
        );

    \I__1491\ : Span4Mux_s3_h
    port map (
            O => \N__10602\,
            I => \N__10599\
        );

    \I__1490\ : Odrv4
    port map (
            O => \N__10599\,
            I => \uu2.mem0.N_82_i\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10593\,
            I => \N__10590\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10590\,
            I => \uu2.mem0.N_110\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10579\
        );

    \I__1485\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10576\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10567\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10567\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10567\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10567\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__10579\,
            I => \N__10564\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10561\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__10567\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1477\ : Odrv4
    port map (
            O => \N__10564\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__10561\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10549\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10546\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10543\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__10549\,
            I => \N__10540\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10535\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10543\,
            I => \N__10535\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__10540\,
            I => \N__10532\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__10535\,
            I => \uu2.N_225\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__10532\,
            I => \uu2.N_225\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__10527\,
            I => \uu2.N_144_cascade_\
        );

    \I__1465\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10521\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__10521\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__10518\,
            I => \uu2.bitmap_RNI1PH82Z0Z_40_cascade_\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__10515\,
            I => \uu2.N_401_cascade_\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10512\,
            I => \N__10509\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10509\,
            I => \uu2.N_406\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10503\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10503\,
            I => \N__10500\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__10500\,
            I => \uu2.un31_w_data_displaying_1\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__10497\,
            I => \N__10494\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10490\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10493\,
            I => \N__10487\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10490\,
            I => \N__10484\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__10487\,
            I => \uu2.un49_w_data_displaying_1\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__10484\,
            I => \uu2.un49_w_data_displaying_1\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__10479\,
            I => \N__10476\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10473\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__10473\,
            I => \N__10470\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__10470\,
            I => \uu2.mem0.N_81_i\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__10467\,
            I => \N__10464\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10464\,
            I => \N__10461\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10461\,
            I => \N__10458\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__10458\,
            I => \N__10455\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__10455\,
            I => \uu2.mem0.N_80_i\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10449\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10449\,
            I => \N__10446\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__1438\ : Odrv4
    port map (
            O => \N__10443\,
            I => \uu2.mem0.N_72_i\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__10440\,
            I => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__10437\,
            I => \uu2.bitmap_pmux_sn_i5_mux_cascade_\
        );

    \I__1435\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10431\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10431\,
            I => \N__10428\
        );

    \I__1433\ : Odrv12
    port map (
            O => \N__10428\,
            I => \uu2.N_404\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__10425\,
            I => \uu2.bitmap_pmux_29_0_cascade_\
        );

    \I__1431\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10416\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10416\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__10416\,
            I => \uu2.bitmap_pmux\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10410\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__10410\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10404\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__10404\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__10401\,
            I => \N__10393\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__10400\,
            I => \N__10390\
        );

    \I__1422\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10376\
        );

    \I__1421\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10376\
        );

    \I__1420\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10376\
        );

    \I__1419\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10376\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10376\
        );

    \I__1417\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10376\
        );

    \I__1416\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10373\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10370\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10367\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__10370\,
            I => \Lab_UT.sec1_3\
        );

    \I__1412\ : Odrv12
    port map (
            O => \N__10367\,
            I => \Lab_UT.sec1_3\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10359\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__10359\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__1409\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10353\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10347\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10347\,
            I => \uu2.bitmap_pmux_24_i_m2_am_1\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__10344\,
            I => \uu2.un51_w_data_displaying_cascade_\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10341\,
            I => \N__10338\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__10338\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10331\
        );

    \I__1401\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10328\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__10331\,
            I => \N__10325\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10322\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__10325\,
            I => \uu2.w_addr_displaying_4_1\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__10322\,
            I => \uu2.w_addr_displaying_4_1\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10314\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__10314\,
            I => \uu2.un51_w_data_displaying\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10311\,
            I => \N__10308\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__10308\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10302\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10302\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10299\,
            I => \uu2.bitmap_RNIAE522Z0Z_93_cascade_\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__10296\,
            I => \N__10293\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10290\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10287\,
            I => \uu2.bitmap_RNIKL222Z0Z_212_cascade_\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10281\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10281\,
            I => \uu2.bitmap_pmux_27_ns_1\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10275\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10275\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10269\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10266\
        );

    \I__1379\ : Odrv4
    port map (
            O => \N__10266\,
            I => vbuf_tx_data_3
        );

    \I__1378\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10260\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10260\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10257\,
            I => \N__10254\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10254\,
            I => \N__10251\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__10251\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10245\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10242\
        );

    \I__1371\ : Odrv12
    port map (
            O => \N__10242\,
            I => vbuf_tx_data_4
        );

    \I__1370\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__10236\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1368\ : CEMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10226\
        );

    \I__1366\ : CEMux
    port map (
            O => \N__10229\,
            I => \N__10223\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__10226\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10223\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1363\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10215\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__10215\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__1361\ : CascadeMux
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10206\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__10203\,
            I => \N__10199\
        );

    \I__1357\ : InMux
    port map (
            O => \N__10202\,
            I => \N__10196\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__10196\,
            I => \N__10190\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10193\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__10190\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10179\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10184\,
            I => \N__10172\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10172\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10172\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__10179\,
            I => \N__10169\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10172\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__10169\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10157\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10157\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10154\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10157\,
            I => \N__10151\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10154\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__10151\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10141\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__10145\,
            I => \N__10137\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__10144\,
            I => \N__10134\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10141\,
            I => \N__10131\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10128\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10123\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10123\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__10131\,
            I => \uu0.un154_ci_9\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__10128\,
            I => \uu0.un154_ci_9\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__10123\,
            I => \uu0.un154_ci_9\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10113\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10113\,
            I => \N__10110\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__10110\,
            I => \uu0.un165_ci_0\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10107\,
            I => \N__10104\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__10101\,
            I => vbuf_tx_data_0
        );

    \I__1323\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10095\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10095\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10089\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1319\ : IoInMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10080\
        );

    \I__1317\ : Span12Mux_s1_h
    port map (
            O => \N__10080\,
            I => \N__10077\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__10077\,
            I => o_serial_data_c
        );

    \I__1315\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10071\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10068\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__10068\,
            I => vbuf_tx_data_1
        );

    \I__1312\ : InMux
    port map (
            O => \N__10065\,
            I => \N__10062\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10062\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1310\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10056\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__10053\,
            I => vbuf_tx_data_2
        );

    \I__1307\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10047\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10047\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10041\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__10041\,
            I => \N__10038\
        );

    \I__1303\ : Sp12to4
    port map (
            O => \N__10038\,
            I => \N__10035\
        );

    \I__1302\ : Odrv12
    port map (
            O => \N__10035\,
            I => \uu2.r_data_wire_1\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10032\,
            I => \N__10029\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10026\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__10026\,
            I => \N__10023\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__10023\,
            I => \uu2.r_data_wire_2\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10020\,
            I => \N__10017\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__10017\,
            I => \N__10014\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__10014\,
            I => \N__10011\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__10011\,
            I => \uu2.r_data_wire_3\
        );

    \I__1293\ : InMux
    port map (
            O => \N__10008\,
            I => \N__10005\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__10002\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__10002\,
            I => \N__9999\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__9999\,
            I => \uu2.r_data_wire_4\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9993\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__9987\,
            I => \uu2.r_data_wire_5\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9981\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__9981\,
            I => vbuf_tx_data_5
        );

    \I__1283\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9975\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__9975\,
            I => \N__9972\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__9972\,
            I => \N__9969\
        );

    \I__1280\ : Odrv4
    port map (
            O => \N__9969\,
            I => \uu2.r_data_wire_6\
        );

    \I__1279\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9963\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9963\,
            I => vbuf_tx_data_6
        );

    \I__1277\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9957\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__1275\ : Span12Mux_s2_h
    port map (
            O => \N__9954\,
            I => \N__9951\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__9951\,
            I => \uu2.r_data_wire_7\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9945\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__9945\,
            I => vbuf_tx_data_7
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__9942\,
            I => \N__9938\
        );

    \I__1270\ : InMux
    port map (
            O => \N__9941\,
            I => \N__9935\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9932\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__9935\,
            I => \N__9929\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9932\,
            I => \N__9923\
        );

    \I__1266\ : Span12Mux_s5_v
    port map (
            O => \N__9929\,
            I => \N__9920\
        );

    \I__1265\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9917\
        );

    \I__1264\ : InMux
    port map (
            O => \N__9927\,
            I => \N__9912\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9912\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__9923\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1261\ : Odrv12
    port map (
            O => \N__9920\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9917\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__9912\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9900\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__1256\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9891\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9898\,
            I => \N__9886\
        );

    \I__1254\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9886\
        );

    \I__1253\ : Odrv12
    port map (
            O => \N__9894\,
            I => \uu2.un404_ci\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__9891\,
            I => \uu2.un404_ci\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9886\,
            I => \uu2.un404_ci\
        );

    \I__1250\ : InMux
    port map (
            O => \N__9879\,
            I => \N__9876\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__9876\,
            I => \N__9869\
        );

    \I__1248\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9860\
        );

    \I__1247\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9860\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9860\
        );

    \I__1245\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9860\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__9869\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__9860\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__9855\,
            I => \N__9851\
        );

    \I__1241\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9848\
        );

    \I__1240\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9845\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__9848\,
            I => \N__9841\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__9845\,
            I => \N__9838\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__9844\,
            I => \N__9834\
        );

    \I__1236\ : Span4Mux_v
    port map (
            O => \N__9841\,
            I => \N__9829\
        );

    \I__1235\ : Span4Mux_h
    port map (
            O => \N__9838\,
            I => \N__9829\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9826\
        );

    \I__1233\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9823\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__9829\,
            I => \N__9820\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9817\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__9823\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__9820\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1228\ : Odrv12
    port map (
            O => \N__9817\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1227\ : CEMux
    port map (
            O => \N__9810\,
            I => \N__9807\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__9804\,
            I => \N__9801\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__9801\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9788\
        );

    \I__1221\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9779\
        );

    \I__1220\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9779\
        );

    \I__1219\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9779\
        );

    \I__1218\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9779\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__9788\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__9779\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__9774\,
            I => \uu2.N_115_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9765\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__9770\,
            I => \N__9761\
        );

    \I__1212\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9756\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9756\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9765\,
            I => \N__9753\
        );

    \I__1209\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9748\
        );

    \I__1208\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9748\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9756\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__9753\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__9748\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1204\ : CEMux
    port map (
            O => \N__9741\,
            I => \N__9738\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__9738\,
            I => \N__9735\
        );

    \I__1202\ : Span4Mux_v
    port map (
            O => \N__9735\,
            I => \N__9731\
        );

    \I__1201\ : CEMux
    port map (
            O => \N__9734\,
            I => \N__9728\
        );

    \I__1200\ : Span4Mux_s1_h
    port map (
            O => \N__9731\,
            I => \N__9725\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9728\,
            I => \N__9722\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__9725\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__1197\ : Odrv12
    port map (
            O => \N__9722\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__1196\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9714\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__9714\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9708\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__9708\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__9705\,
            I => \N__9701\
        );

    \I__1191\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9696\
        );

    \I__1190\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9689\
        );

    \I__1189\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9689\
        );

    \I__1188\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9689\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__9696\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9689\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9678\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__1182\ : Span4Mux_h
    port map (
            O => \N__9675\,
            I => \N__9672\
        );

    \I__1181\ : Span4Mux_v
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__9669\,
            I => \uu2.mem0.N_78_i\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__9666\,
            I => \N__9663\
        );

    \I__1178\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9660\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9657\
        );

    \I__1176\ : Span4Mux_v
    port map (
            O => \N__9657\,
            I => \N__9654\
        );

    \I__1175\ : Odrv4
    port map (
            O => \N__9654\,
            I => \uu2.mem0.N_77_i\
        );

    \I__1174\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9648\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__1172\ : Sp12to4
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__1171\ : Odrv12
    port map (
            O => \N__9642\,
            I => \uu2.r_data_wire_0\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__9639\,
            I => \N__9636\
        );

    \I__1169\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9633\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__9633\,
            I => \N__9630\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__9627\,
            I => \uu2.mem0.N_75_i\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__9615\,
            I => \N__9612\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__9612\,
            I => \uu2.mem0.N_74_i\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__9609\,
            I => \N__9605\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9600\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9595\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9595\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9592\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__9600\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9595\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__9592\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9581\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9584\,
            I => \N__9577\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9574\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9571\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__9577\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__9574\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9571\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1145\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9561\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9561\,
            I => \uu2.N_186\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9555\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__9555\,
            I => \uu2.w_addr_user_3_i_a2_2_6\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__9552\,
            I => \uu2.N_150_cascade_\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__9540\,
            I => \uu2.mem0.N_79_i\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9533\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9530\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9527\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9530\,
            I => \N__9524\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__9527\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__9524\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9516\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9516\,
            I => \uu0.sec_clkDZ0\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__9513\,
            I => \oneSecStrb_cascade_\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__9510\,
            I => \uu2.N_118_cascade_\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9504\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__9504\,
            I => \uu2.N_117\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__9501\,
            I => \uu2.N_117_cascade_\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__9498\,
            I => \uu2.un404_ci_cascade_\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9492\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__9492\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__9489\,
            I => \N__9486\
        );

    \I__1119\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9481\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9476\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9476\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9481\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9476\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9468\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9468\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__9465\,
            I => \N__9461\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__9464\,
            I => \N__9457\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9453\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9450\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9445\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9445\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__9453\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__9450\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9445\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__9438\,
            I => \N__9435\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9431\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__9434\,
            I => \N__9428\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9425\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9420\
        );

    \I__1098\ : Span4Mux_h
    port map (
            O => \N__9425\,
            I => \N__9417\
        );

    \I__1097\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9412\
        );

    \I__1096\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9412\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__9420\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__9417\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9412\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__9405\,
            I => \N__9402\
        );

    \I__1091\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9399\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__9399\,
            I => \N__9392\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9387\
        );

    \I__1088\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9387\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9382\
        );

    \I__1086\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9382\
        );

    \I__1085\ : Odrv4
    port map (
            O => \N__9392\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9387\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__9382\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9368\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__9371\,
            I => \N__9364\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9368\,
            I => \N__9358\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9351\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9351\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9351\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9346\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9361\,
            I => \N__9346\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__9358\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9351\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9346\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1070\ : CascadeMux
    port map (
            O => \N__9339\,
            I => \N__9334\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__9338\,
            I => \N__9331\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9328\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9325\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9320\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9320\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9325\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9320\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1062\ : CEMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9312\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__9309\,
            I => \N__9306\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9303\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9303\,
            I => \uu2.mem0.N_76_i\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__9300\,
            I => \N__9297\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9294\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9294\,
            I => \N__9291\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__9291\,
            I => \uu2.mem0.N_73_i\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__9288\,
            I => \N__9282\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9275\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9286\,
            I => \N__9272\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9269\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9262\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9262\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9262\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__9279\,
            I => \N__9258\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__9278\,
            I => \N__9255\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9245\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9272\,
            I => \N__9245\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9269\,
            I => \N__9245\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9262\,
            I => \N__9245\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9236\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9236\
        );

    \I__1038\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9236\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9236\
        );

    \I__1036\ : Odrv12
    port map (
            O => \N__9245\,
            I => \uu0.un110_ci\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__9236\,
            I => \uu0.un110_ci\
        );

    \I__1034\ : CEMux
    port map (
            O => \N__9231\,
            I => \N__9213\
        );

    \I__1033\ : CEMux
    port map (
            O => \N__9230\,
            I => \N__9213\
        );

    \I__1032\ : CEMux
    port map (
            O => \N__9229\,
            I => \N__9213\
        );

    \I__1031\ : CEMux
    port map (
            O => \N__9228\,
            I => \N__9213\
        );

    \I__1030\ : CEMux
    port map (
            O => \N__9227\,
            I => \N__9213\
        );

    \I__1029\ : CEMux
    port map (
            O => \N__9226\,
            I => \N__9213\
        );

    \I__1028\ : GlobalMux
    port map (
            O => \N__9213\,
            I => \N__9210\
        );

    \I__1027\ : gio2CtrlBuf
    port map (
            O => \N__9210\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__9207\,
            I => \uu2.trig_rd_is_det_cascade_\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9204\,
            I => \N__9198\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9198\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9198\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9192\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__9192\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__9189\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__9186\,
            I => \N__9183\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9179\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9176\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9179\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__9176\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9166\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9163\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9160\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9166\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9163\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9160\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__9153\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__9150\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__9147\,
            I => \N__9143\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9140\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9137\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__9140\,
            I => \N__9129\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9129\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9122\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9122\
        );

    \I__999\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9122\
        );

    \I__998\ : Odrv12
    port map (
            O => \N__9129\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__9122\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__996\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9105\
        );

    \I__995\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9105\
        );

    \I__994\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9105\
        );

    \I__993\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9105\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9105\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__991\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9099\,
            I => \N__9093\
        );

    \I__989\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9088\
        );

    \I__988\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9088\
        );

    \I__987\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9085\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__9093\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9088\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9085\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__9078\,
            I => \N__9073\
        );

    \I__982\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9070\
        );

    \I__981\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9065\
        );

    \I__980\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9065\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9070\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__9065\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__977\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9057\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9057\,
            I => \uu0.un4_l_count_13\
        );

    \I__975\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9051\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9051\,
            I => \N__9046\
        );

    \I__973\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9043\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__9049\,
            I => \N__9039\
        );

    \I__971\ : Span4Mux_s2_v
    port map (
            O => \N__9046\,
            I => \N__9034\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9043\,
            I => \N__9034\
        );

    \I__969\ : InMux
    port map (
            O => \N__9042\,
            I => \N__9031\
        );

    \I__968\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9028\
        );

    \I__967\ : Odrv4
    port map (
            O => \N__9034\,
            I => \uu0.un66_ci\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9031\,
            I => \uu0.un66_ci\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9028\,
            I => \uu0.un66_ci\
        );

    \I__964\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9017\
        );

    \I__963\ : InMux
    port map (
            O => \N__9020\,
            I => \N__9012\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__9009\
        );

    \I__961\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9004\
        );

    \I__960\ : InMux
    port map (
            O => \N__9015\,
            I => \N__9004\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9012\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__958\ : Odrv12
    port map (
            O => \N__9009\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__9004\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__956\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8994\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__8994\,
            I => \N__8990\
        );

    \I__954\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8987\
        );

    \I__953\ : Span4Mux_v
    port map (
            O => \N__8990\,
            I => \N__8981\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__8987\,
            I => \N__8981\
        );

    \I__951\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8978\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__8981\,
            I => \N__8975\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__8978\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__948\ : Odrv4
    port map (
            O => \N__8975\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__946\ : InMux
    port map (
            O => \N__8967\,
            I => \N__8958\
        );

    \I__945\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8958\
        );

    \I__944\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8954\
        );

    \I__943\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8951\
        );

    \I__942\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8948\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__8958\,
            I => \N__8945\
        );

    \I__940\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8942\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__8954\,
            I => \N__8939\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8951\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8948\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__8945\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__8942\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__934\ : Odrv12
    port map (
            O => \N__8939\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__933\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8922\
        );

    \I__932\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8915\
        );

    \I__931\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8915\
        );

    \I__930\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8915\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8922\,
            I => \N__8912\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__8915\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__8912\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__926\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__8904\,
            I => \uu0.un44_ci\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__8901\,
            I => \N__8898\
        );

    \I__923\ : InMux
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8889\
        );

    \I__921\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8884\
        );

    \I__920\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8884\
        );

    \I__919\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8881\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__8889\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__8884\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__8881\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__915\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8869\
        );

    \I__914\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8864\
        );

    \I__913\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8864\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__8869\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8864\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__8859\,
            I => \N__8856\
        );

    \I__909\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8853\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8853\,
            I => \N__8850\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__8850\,
            I => \uu0.un99_ci_0\
        );

    \I__906\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8842\
        );

    \I__905\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8837\
        );

    \I__904\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8837\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__8842\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8837\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__901\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8829\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__8829\,
            I => \uu0.un220_ci\
        );

    \I__899\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8822\
        );

    \I__898\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8817\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8814\
        );

    \I__896\ : InMux
    port map (
            O => \N__8821\,
            I => \N__8809\
        );

    \I__895\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8809\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__8817\,
            I => \N__8806\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__8814\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__8809\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__891\ : Odrv4
    port map (
            O => \N__8806\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__890\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__8796\,
            I => \uu0.un4_l_count_11\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__8793\,
            I => \N__8789\
        );

    \I__887\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8784\
        );

    \I__886\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8784\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__8784\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__884\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__8778\,
            I => \N__8775\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__8775\,
            I => \uu0.un4_l_count_18\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__8772\,
            I => \uu0.un4_l_count_16_cascade_\
        );

    \I__880\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8766\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8763\
        );

    \I__878\ : Odrv4
    port map (
            O => \N__8763\,
            I => \uu0.un4_l_count_12\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__8760\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__876\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8754\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__8754\,
            I => \uu0.un143_ci_0\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__8751\,
            I => \N__8746\
        );

    \I__873\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8739\
        );

    \I__872\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8739\
        );

    \I__871\ : InMux
    port map (
            O => \N__8746\,
            I => \N__8739\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8739\,
            I => \N__8736\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__8736\,
            I => \uu0.un198_ci_2\
        );

    \I__868\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8720\
        );

    \I__867\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8720\
        );

    \I__866\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8720\
        );

    \I__865\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8720\
        );

    \I__864\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8717\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__8720\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__8717\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \N__8707\
        );

    \I__860\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8699\
        );

    \I__859\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8699\
        );

    \I__858\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8699\
        );

    \I__857\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8696\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__8699\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__8696\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__854\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8684\
        );

    \I__853\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8684\
        );

    \I__852\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8681\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8684\,
            I => \N__8678\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8681\,
            I => \uu0.un88_ci_3\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__8678\,
            I => \uu0.un88_ci_3\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__8670\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__8667\,
            I => \N__8662\
        );

    \I__845\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8655\
        );

    \I__844\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8655\
        );

    \I__843\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8655\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__8655\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__8652\,
            I => \N__8647\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__8651\,
            I => \N__8644\
        );

    \I__839\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8637\
        );

    \I__838\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8637\
        );

    \I__837\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8637\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8637\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__835\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8619\
        );

    \I__834\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8619\
        );

    \I__833\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8619\
        );

    \I__832\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8619\
        );

    \I__831\ : InMux
    port map (
            O => \N__8630\,
            I => \N__8619\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8619\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__8616\,
            I => \N__8610\
        );

    \I__828\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8601\
        );

    \I__827\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8601\
        );

    \I__826\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8601\
        );

    \I__825\ : InMux
    port map (
            O => \N__8610\,
            I => \N__8601\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8601\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__822\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8579\
        );

    \I__821\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8579\
        );

    \I__820\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8579\
        );

    \I__819\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8579\
        );

    \I__818\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8579\
        );

    \I__817\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8576\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8579\,
            I => \N__8573\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__8576\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__814\ : Odrv12
    port map (
            O => \N__8573\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__8568\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__8565\,
            I => \uu0.un44_ci_cascade_\
        );

    \I__811\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8557\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__8561\,
            I => \N__8552\
        );

    \I__809\ : InMux
    port map (
            O => \N__8560\,
            I => \N__8549\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8546\
        );

    \I__807\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8539\
        );

    \I__806\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8539\
        );

    \I__805\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8539\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8549\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__8546\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8539\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__801\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8526\
        );

    \I__800\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8523\
        );

    \I__799\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8520\
        );

    \I__798\ : InMux
    port map (
            O => \N__8529\,
            I => \N__8515\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8510\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__8523\,
            I => \N__8510\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8507\
        );

    \I__794\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8502\
        );

    \I__793\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8502\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__8515\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__791\ : Odrv12
    port map (
            O => \N__8510\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__8507\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8502\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__8493\,
            I => \N__8490\
        );

    \I__787\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8484\
        );

    \I__786\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8484\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__8481\,
            I => \uu2.un284_ci\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__782\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8470\
        );

    \I__781\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8467\
        );

    \I__780\ : InMux
    port map (
            O => \N__8473\,
            I => \N__8464\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__8470\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__8467\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__8464\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__8457\,
            I => \N__8452\
        );

    \I__775\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8447\
        );

    \I__774\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8447\
        );

    \I__773\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8444\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8447\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__8444\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__770\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8430\
        );

    \I__769\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8430\
        );

    \I__768\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8430\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__8430\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__765\ : InMux
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8421\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__763\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8403\
        );

    \I__762\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8403\
        );

    \I__761\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8403\
        );

    \I__760\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8403\
        );

    \I__759\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8403\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8403\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__8400\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__756\ : InMux
    port map (
            O => \N__8397\,
            I => \N__8394\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8394\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__754\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8386\
        );

    \I__753\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8383\
        );

    \I__752\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8380\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8386\,
            I => \N__8377\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__8383\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8380\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__8377\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__8370\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8358\
        );

    \I__745\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8358\
        );

    \I__744\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8351\
        );

    \I__743\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8351\
        );

    \I__742\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8351\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8358\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8351\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__739\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8337\
        );

    \I__738\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8337\
        );

    \I__737\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8330\
        );

    \I__736\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8330\
        );

    \I__735\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8330\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__8337\,
            I => \uu2.un306_ci\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__8330\,
            I => \uu2.un306_ci\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__8325\,
            I => \N__8321\
        );

    \I__731\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8317\
        );

    \I__730\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8312\
        );

    \I__729\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8312\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8317\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__8312\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__726\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8301\
        );

    \I__724\ : IoSpan4Mux
    port map (
            O => \N__8301\,
            I => \N__8298\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__8298\,
            I => \uart_RXD\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__8295\,
            I => \N__8290\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__8294\,
            I => \N__8287\
        );

    \I__720\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8280\
        );

    \I__719\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8280\
        );

    \I__718\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8280\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8280\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__716\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8271\
        );

    \I__715\ : InMux
    port map (
            O => \N__8276\,
            I => \N__8271\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__8271\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__8268\,
            I => \uu2.vbuf_count.un328_ci_3_cascade_\
        );

    \I__712\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8250\
        );

    \I__711\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8250\
        );

    \I__710\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8250\
        );

    \I__709\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8250\
        );

    \I__708\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8250\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__8250\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__8247\,
            I => \N__8244\
        );

    \I__705\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__8241\,
            I => \uu2.un350_ci\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__8238\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__702\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__8232\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__700\ : IoInMux
    port map (
            O => \N__8229\,
            I => \N__8226\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8223\
        );

    \I__698\ : Span12Mux_s5_v
    port map (
            O => \N__8223\,
            I => \N__8220\
        );

    \I__697\ : Odrv12
    port map (
            O => \N__8220\,
            I => \latticehx1k_pll_inst.clk\
        );

    \I__696\ : IoInMux
    port map (
            O => \N__8217\,
            I => \N__8214\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8211\
        );

    \I__694\ : IoSpan4Mux
    port map (
            O => \N__8211\,
            I => \N__8208\
        );

    \I__693\ : Odrv4
    port map (
            O => \N__8208\,
            I => clk_in_c
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__22806\
        );

    \INVuu2.w_addr_displaying_ness_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_ness_6C_net\,
            I => \N__22814\
        );

    \INVuu2.w_addr_displaying_2C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2C_net\,
            I => \N__22799\
        );

    \INVuu2.w_addr_displaying_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_3C_net\,
            I => \N__22811\
        );

    \INVuu2.w_addr_displaying_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_8C_net\,
            I => \N__22818\
        );

    \INVuu2.bitmap_69C\ : INV
    port map (
            O => \INVuu2.bitmap_69C_net\,
            I => \N__22822\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__22831\
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__22846\
        );

    \INVuu2.bitmap_40C\ : INV
    port map (
            O => \INVuu2.bitmap_40C_net\,
            I => \N__22810\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__22830\
        );

    \INVuu2.bitmap_215C\ : INV
    port map (
            O => \INVuu2.bitmap_215C_net\,
            I => \N__22838\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__22845\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__22794\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__22802\
        );

    \INVuu2.w_addr_user_nesr_7C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_7C_net\,
            I => \N__22809\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_12_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_3_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8229\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \bu_rx_data_rdy_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22338\,
            GLOBALBUFFEROUTPUT => bu_rx_data_rdy_0_g
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16569\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \buart.Z_rx.sample_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19218\,
            GLOBALBUFFEROUTPUT => \buart__rx_sample_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__19647\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.vram_rd_clk_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12198\,
            in2 => \_gnd_net_\,
            in3 => \N__8391\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22854\,
            ce => 'H',
            sr => \N__22516\
        );

    \uu2.l_count_0_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8529\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22851\,
            ce => 'H',
            sr => \N__22495\
        );

    \uu2.trig_rd_det_0_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12199\,
            in2 => \_gnd_net_\,
            in3 => \N__9536\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22851\,
            ce => 'H',
            sr => \N__22495\
        );

    \uu2.l_count_6_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__8276\,
            in2 => \_gnd_net_\,
            in3 => \N__8264\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22843\,
            ce => 'H',
            sr => \N__22512\
        );

    \uu2.l_count_RNIBCGK1_9_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8262\,
            in1 => \N__8519\,
            in2 => \N__8295\,
            in3 => \N__8364\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__8456\,
            in1 => \N__8293\,
            in2 => \N__8247\,
            in3 => \N__8390\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22843\,
            ce => 'H',
            sr => \N__22512\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8261\,
            in1 => \N__8518\,
            in2 => \N__8294\,
            in3 => \N__8363\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_7_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8344\,
            in1 => \N__8265\,
            in2 => \N__8478\,
            in3 => \N__8277\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22843\,
            ce => 'H',
            sr => \N__22512\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8324\,
            in2 => \_gnd_net_\,
            in3 => \N__8365\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => \uu2.vbuf_count.un328_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8342\,
            in1 => \N__8474\,
            in2 => \N__8268\,
            in3 => \N__8263\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8238\,
            in3 => \N__8455\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22843\,
            ce => 'H',
            sr => \N__22512\
        );

    \uu2.l_count_RNI9S834_0_1_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8415\,
            in1 => \N__8555\,
            in2 => \N__8427\,
            in3 => \N__8235\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8489\,
            in2 => \_gnd_net_\,
            in3 => \N__8417\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22836\,
            ce => 'H',
            sr => \N__22510\
        );

    \uu2.l_count_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8418\,
            in1 => \N__8389\,
            in2 => \N__8493\,
            in3 => \N__8439\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22836\,
            ce => 'H',
            sr => \N__22510\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8438\,
            in1 => \N__8530\,
            in2 => \N__8561\,
            in3 => \N__8414\,
            lcout => \uu2.un306_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIFGGK1_3_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8473\,
            in1 => \N__8320\,
            in2 => \N__8457\,
            in3 => \N__8437\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8556\,
            in1 => \N__8416\,
            in2 => \N__8400\,
            in3 => \N__8397\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__8346\,
            in1 => \_gnd_net_\,
            in2 => \N__8370\,
            in3 => \N__8366\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22836\,
            ce => 'H',
            sr => \N__22510\
        );

    \uu2.l_count_5_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__8367\,
            in1 => \_gnd_net_\,
            in2 => \N__8325\,
            in3 => \N__8345\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22836\,
            ce => 'H',
            sr => \N__22510\
        );

    \uu0.sec_clk_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12238\,
            in2 => \_gnd_net_\,
            in3 => \N__16637\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \uu2.l_count_1_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8560\,
            in2 => \_gnd_net_\,
            in3 => \N__8532\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \buart.Z_rx.hh_0_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_hh_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \buart.Z_rx.hh_1_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19487\,
            lcout => \buart__rx_hh_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \uu0.delay_line_1_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16316\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \uu0.l_precount_0_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8590\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22827\,
            ce => 'H',
            sr => \N__22508\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8997\,
            in2 => \_gnd_net_\,
            in3 => \N__9021\,
            lcout => \uu0.un88_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8689\,
            in2 => \_gnd_net_\,
            in3 => \N__8826\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8562\,
            in2 => \_gnd_net_\,
            in3 => \N__8531\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI2Q224_6_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22556\,
            in2 => \_gnd_net_\,
            in3 => \N__12378\,
            lcout => \uu2.un28_w_addr_user_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12841\,
            in2 => \_gnd_net_\,
            in3 => \N__12880\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22816\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22816\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8631\,
            in1 => \N__8592\,
            in2 => \N__8652\,
            in3 => \N__8613\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22808\,
            ce => 'H',
            sr => \N__22509\
        );

    \uu0.l_precount_3_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8615\,
            in1 => \N__8650\,
            in2 => \N__8598\,
            in3 => \N__8634\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22808\,
            ce => 'H',
            sr => \N__22509\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8630\,
            in1 => \N__8993\,
            in2 => \N__8651\,
            in3 => \N__8706\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_1_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8593\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8632\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22808\,
            ce => 'H',
            sr => \N__22509\
        );

    \uu0.l_precount_2_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8633\,
            in1 => \N__8594\,
            in2 => \_gnd_net_\,
            in3 => \N__8614\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22808\,
            ce => 'H',
            sr => \N__22509\
        );

    \uu0.l_precount_RNI3Q7K1_2_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8965\,
            in1 => \N__8892\,
            in2 => \N__8616\,
            in3 => \N__8729\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIO2782_16_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__10185\,
            in1 => \N__8591\,
            in2 => \N__8568\,
            in3 => \N__8928\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_6_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__8691\,
            in1 => \N__8821\,
            in2 => \N__9049\,
            in3 => \N__16635\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22801\,
            ce => \N__9226\,
            sr => \N__22511\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8731\,
            lcout => \uu0.un44_ci\,
            ltout => \uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8565\,
            in3 => \N__8894\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22801\,
            ce => \N__9226\,
            sr => \N__22511\
        );

    \uu0.l_count_1_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8711\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8733\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22801\,
            ce => \N__9226\,
            sr => \N__22511\
        );

    \uu0.l_count_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8732\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16633\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22801\,
            ce => \N__9226\,
            sr => \N__22511\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8893\,
            in1 => \N__8730\,
            in2 => \N__8712\,
            in3 => \N__8874\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8690\,
            in1 => \N__8820\,
            in2 => \N__8673\,
            in3 => \N__8847\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_12_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__16634\,
            in1 => \N__10146\,
            in2 => \N__8670\,
            in3 => \N__10162\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22801\,
            ce => \N__9226\,
            sr => \N__22511\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__9134\,
            in1 => \N__8845\,
            in2 => \N__8667\,
            in3 => \N__8872\,
            lcout => \uu0.un4_l_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9102\,
            in1 => \N__8966\,
            in2 => \_gnd_net_\,
            in3 => \N__9135\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_9_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__9136\,
            in1 => \_gnd_net_\,
            in2 => \N__8970\,
            in3 => \N__9261\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22797\,
            ce => \N__9227\,
            sr => \N__22513\
        );

    \uu0.l_count_17_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8927\,
            in1 => \N__8666\,
            in2 => \N__9279\,
            in3 => \N__8750\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22797\,
            ce => \N__9227\,
            sr => \N__22513\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8665\,
            in1 => \N__9254\,
            in2 => \N__8751\,
            in3 => \N__8925\,
            lcout => \uu0.un220_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__8749\,
            in2 => \N__9278\,
            in3 => \N__16621\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22797\,
            ce => \N__9227\,
            sr => \N__22513\
        );

    \uu0.l_count_3_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__16623\,
            in1 => \N__8907\,
            in2 => \N__8901\,
            in3 => \N__8873\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22797\,
            ce => \N__9227\,
            sr => \N__22513\
        );

    \uu0.l_count_7_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8846\,
            in1 => \N__9042\,
            in2 => \N__8859\,
            in3 => \N__16622\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22797\,
            ce => \N__9227\,
            sr => \N__22513\
        );

    \uu0.l_count_18_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__8792\,
            in2 => \_gnd_net_\,
            in3 => \N__16618\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22793\,
            ce => \N__9228\,
            sr => \N__22515\
        );

    \uu0.l_count_RNIOIDD2_18_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8825\,
            in1 => \N__8799\,
            in2 => \N__8793\,
            in3 => \N__9169\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_15_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9060\,
            in1 => \N__8781\,
            in2 => \N__8772\,
            in3 => \N__8769\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_11_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__9171\,
            in1 => \N__9287\,
            in2 => \N__8760\,
            in3 => \N__8757\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22793\,
            ce => \N__9228\,
            sr => \N__22515\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__9115\,
            in2 => \N__10144\,
            in3 => \N__10182\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9097\,
            in1 => \N__8957\,
            in2 => \N__9147\,
            in3 => \N__9170\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9116\,
            in2 => \N__9153\,
            in3 => \N__10183\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9076\,
            in1 => \N__9281\,
            in2 => \N__9150\,
            in3 => \N__16619\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22789\,
            ce => \N__9229\,
            sr => \N__22517\
        );

    \uu0.l_count_14_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9280\,
            in1 => \N__9117\,
            in2 => \N__10145\,
            in3 => \N__10184\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22789\,
            ce => \N__9229\,
            sr => \N__22517\
        );

    \uu0.l_count_4_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9050\,
            in1 => \N__9016\,
            in2 => \_gnd_net_\,
            in3 => \N__16620\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22789\,
            ce => \N__9229\,
            sr => \N__22517\
        );

    \uu0.l_count_10_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9146\,
            in1 => \N__8964\,
            in2 => \N__9288\,
            in3 => \N__9098\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22789\,
            ce => \N__9229\,
            sr => \N__22517\
        );

    \uu0.l_count_RNIGTCU_15_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9114\,
            in1 => \N__9096\,
            in2 => \N__9078\,
            in3 => \N__9015\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_5_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9054\,
            in1 => \N__8986\,
            in2 => \_gnd_net_\,
            in3 => \N__9020\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22785\,
            ce => \N__9230\,
            sr => \N__22518\
        );

    \uu0.l_count_8_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9286\,
            in2 => \_gnd_net_\,
            in3 => \N__8963\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22785\,
            ce => \N__9230\,
            sr => \N__22518\
        );

    \uu0.l_count_13_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__9285\,
            in1 => \N__10116\,
            in2 => \N__10203\,
            in3 => \N__16636\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22782\,
            ce => \N__9231\,
            sr => \N__22521\
        );

    \uu2.r_addr_2_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9398\,
            in1 => \N__9367\,
            in2 => \N__9434\,
            in3 => \N__9875\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22844\,
            ce => 'H',
            sr => \N__22497\
        );

    \uu2.r_addr_1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__9873\,
            in1 => \_gnd_net_\,
            in2 => \N__9371\,
            in3 => \N__9397\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22844\,
            ce => 'H',
            sr => \N__22497\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9872\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9195\,
            in2 => \_gnd_net_\,
            in3 => \N__9203\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => \uu2.trig_rd_is_det_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_0_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9207\,
            in3 => \N__9363\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22844\,
            ce => 'H',
            sr => \N__22497\
        );

    \uu2.trig_rd_det_1_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9204\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22844\,
            ce => 'H',
            sr => \N__22497\
        );

    \uu2.r_addr_4_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9874\,
            in1 => \N__9928\,
            in2 => \_gnd_net_\,
            in3 => \N__9899\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22844\,
            ce => 'H',
            sr => \N__22497\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9837\,
            in2 => \_gnd_net_\,
            in3 => \N__9926\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9182\,
            in1 => \N__9471\,
            in2 => \N__9189\,
            in3 => \N__9898\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22837\,
            ce => \N__9315\,
            sr => \N__22496\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9423\,
            in1 => \N__9395\,
            in2 => \N__9337\,
            in3 => \N__9361\,
            lcout => \uu2.un404_ci\,
            ltout => \uu2.un404_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_7_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9485\,
            in1 => \N__9460\,
            in2 => \N__9498\,
            in3 => \N__9495\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22837\,
            ce => \N__9315\,
            sr => \N__22496\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9484\,
            in2 => \_gnd_net_\,
            in3 => \N__9456\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9927\,
            in1 => \N__9854\,
            in2 => \N__9464\,
            in3 => \N__9897\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22837\,
            ce => \N__9315\,
            sr => \N__22496\
        );

    \uu2.r_addr_esr_3_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9424\,
            in1 => \N__9396\,
            in2 => \N__9338\,
            in3 => \N__9362\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22837\,
            ce => \N__9315\,
            sr => \N__22496\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9771\,
            in1 => \N__11718\,
            in2 => \_gnd_net_\,
            in3 => \N__13389\,
            lcout => \uu2.mem0.N_76_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI84IJ2_2_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__11895\,
            in1 => \N__13171\,
            in2 => \N__13521\,
            in3 => \N__13721\,
            lcout => \uu2.bitmap_pmux_sn_N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9585\,
            in1 => \N__11713\,
            in2 => \_gnd_net_\,
            in3 => \N__13827\,
            lcout => \uu2.mem0.N_73_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12239\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.sec_clkDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22821\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9798\,
            in1 => \N__11712\,
            in2 => \_gnd_net_\,
            in3 => \N__11893\,
            lcout => \uu2.mem0.N_79_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__12207\,
            in1 => \N__9537\,
            in2 => \N__11007\,
            in3 => \N__22560\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22817\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9519\,
            in2 => \_gnd_net_\,
            in3 => \N__12234\,
            lcout => \oneSecStrb\,
            ltout => \oneSecStrb_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__12503\,
            in1 => \N__10709\,
            in2 => \N__9513\,
            in3 => \N__15090\,
            lcout => \Lab_UT.dispString.un46_dOutP_i_m_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_7_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__12319\,
            in1 => \N__9507\,
            in2 => \N__9609\,
            in3 => \N__10583\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_7C_net\,
            ce => \N__9734\,
            sr => \N__22472\
        );

    \uu2.w_addr_user_nesr_RNO_0_8_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__10582\,
            in1 => \N__9769\,
            in2 => \N__12356\,
            in3 => \N__12284\,
            lcout => OPEN,
            ltout => \uu2.N_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000100000100"
        )
    port map (
            in0 => \N__12320\,
            in1 => \N__9608\,
            in2 => \N__9510\,
            in3 => \N__9584\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_7C_net\,
            ce => \N__9734\,
            sr => \N__22472\
        );

    \uu2.w_addr_user_nesr_RNIHSS8_5_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__12348\,
            in1 => \N__9768\,
            in2 => \_gnd_net_\,
            in3 => \N__12283\,
            lcout => \uu2.N_117\,
            ltout => \uu2.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_6_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000001"
        )
    port map (
            in0 => \N__12318\,
            in1 => \N__10553\,
            in2 => \N__9501\,
            in3 => \N__10585\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_7C_net\,
            ce => \N__9734\,
            sr => \N__22472\
        );

    \uu2.w_addr_user_nesr_0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__10584\,
            in1 => \N__10552\,
            in2 => \N__11824\,
            in3 => \N__12317\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_7C_net\,
            ce => \N__9734\,
            sr => \N__22472\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10586\,
            in1 => \N__11710\,
            in2 => \_gnd_net_\,
            in3 => \N__13260\,
            lcout => \uu2.mem0.N_75_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11711\,
            in1 => \N__9604\,
            in2 => \_gnd_net_\,
            in3 => \N__13350\,
            lcout => \uu2.mem0.N_74_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIG9RA_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11811\,
            in1 => \N__9558\,
            in2 => \N__11779\,
            in3 => \N__9564\,
            lcout => \uu2.N_225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIVCU1_8_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9603\,
            in2 => \_gnd_net_\,
            in3 => \N__9580\,
            lcout => \uu2.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNINJD5_3_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12281\,
            in1 => \N__9699\,
            in2 => \N__9770\,
            in3 => \N__9791\,
            lcout => \uu2.w_addr_user_3_i_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNO_0_3_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9793\,
            in1 => \N__11775\,
            in2 => \N__9705\,
            in3 => \N__11813\,
            lcout => OPEN,
            ltout => \uu2.N_150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__12329\,
            in1 => \_gnd_net_\,
            in2 => \N__9552\,
            in3 => \N__12352\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__9741\,
            sr => \N__22473\
        );

    \uu2.w_addr_user_nesr_2_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9794\,
            in1 => \N__11814\,
            in2 => \N__11781\,
            in3 => \N__12328\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__9741\,
            sr => \N__22473\
        );

    \uu2.w_addr_user_nesr_RNIFBD5_3_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__11812\,
            in1 => \N__9700\,
            in2 => \N__11780\,
            in3 => \N__9792\,
            lcout => \uu2.N_115\,
            ltout => \uu2.N_115_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_5_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000110"
        )
    port map (
            in0 => \N__12285\,
            in1 => \N__9764\,
            in2 => \N__9774\,
            in3 => \N__12330\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__9741\,
            sr => \N__22473\
        );

    \buart.Z_tx.shifter_6_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10983\,
            in1 => \N__9717\,
            in2 => \_gnd_net_\,
            in3 => \N__9984\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22798\,
            ce => \N__10229\,
            sr => \N__22514\
        );

    \buart.Z_tx.shifter_7_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9711\,
            in1 => \N__10984\,
            in2 => \_gnd_net_\,
            in3 => \N__9966\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22798\,
            ce => \N__10229\,
            sr => \N__22514\
        );

    \buart.Z_tx.shifter_8_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9948\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22798\,
            ce => \N__10229\,
            sr => \N__22514\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__11066\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9704\,
            in1 => \N__11708\,
            in2 => \_gnd_net_\,
            in3 => \N__13728\,
            lcout => \uu2.mem0.N_78_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11709\,
            in1 => \N__12282\,
            in2 => \_gnd_net_\,
            in3 => \N__13506\,
            lcout => \uu2.mem0.N_77_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9651\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10044\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10008\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9996\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9978\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__9810\,
            sr => \_gnd_net_\
        );

    \uu2.r_addr_5_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9941\,
            in1 => \N__9903\,
            in2 => \N__9844\,
            in3 => \N__9879\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22790\,
            ce => 'H',
            sr => \N__22555\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12156\,
            in1 => \N__12177\,
            in2 => \_gnd_net_\,
            in3 => \N__22554\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11010\,
            in1 => \N__10934\,
            in2 => \_gnd_net_\,
            in3 => \N__11067\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22790\,
            ce => 'H',
            sr => \N__22555\
        );

    \uu0.l_count_RNIFAQ9_13_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10202\,
            in2 => \_gnd_net_\,
            in3 => \N__10163\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10164\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10140\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11011\,
            in1 => \N__10065\,
            in2 => \_gnd_net_\,
            in3 => \N__10107\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.shifter_0_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10098\,
            in2 => \_gnd_net_\,
            in3 => \N__11015\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.uart_tx_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11008\,
            in2 => \_gnd_net_\,
            in3 => \N__10092\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.shifter_2_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11009\,
            in1 => \N__10050\,
            in2 => \_gnd_net_\,
            in3 => \N__10074\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.shifter_3_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11012\,
            in1 => \N__10263\,
            in2 => \_gnd_net_\,
            in3 => \N__10059\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.shifter_4_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10239\,
            in1 => \N__11014\,
            in2 => \_gnd_net_\,
            in3 => \N__10272\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \buart.Z_tx.shifter_5_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11013\,
            in1 => \N__10257\,
            in2 => \_gnd_net_\,
            in3 => \N__10248\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22786\,
            ce => \N__10233\,
            sr => \N__22519\
        );

    \Lab_UT.didp.regrce1.q_RNI2NVO3_1_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14973\,
            in1 => \N__15465\,
            in2 => \N__15059\,
            in3 => \N__14034\,
            lcout => \Lab_UT.sec2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNI4PVO3_2_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14976\,
            in1 => \N__15390\,
            in2 => \N__13995\,
            in3 => \N__15055\,
            lcout => \Lab_UT.sec2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNI6RVO3_3_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14974\,
            in1 => \N__15431\,
            in2 => \N__15060\,
            in3 => \N__13946\,
            lcout => \Lab_UT.sec2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI85KT3_3_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__14636\,
            in1 => \N__15051\,
            in2 => \N__17687\,
            in3 => \N__14975\,
            lcout => \Lab_UT.sec1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNIK3221_3_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__15430\,
            in1 => \N__14635\,
            in2 => \N__17688\,
            in3 => \N__13945\,
            lcout => \Lab_UT.didp.did_alarmMatch_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__13044\,
            in1 => \N__11242\,
            in2 => \N__11217\,
            in3 => \N__11288\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__22482\
        );

    \uu2.bitmap_221_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__11241\,
            in1 => \N__11208\,
            in2 => \N__11292\,
            in3 => \N__13043\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__22482\
        );

    \uu2.bitmap_RNIAE522_93_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__13155\,
            in1 => \N__10218\,
            in2 => \N__10212\,
            in3 => \N__10881\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNIAE522Z0Z_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIMS86A_66_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__10335\,
            in1 => \N__13059\,
            in2 => \N__10299\,
            in3 => \N__10284\,
            lcout => \uu2.N_404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__11147\,
            in1 => \N__10389\,
            in2 => \N__11118\,
            in3 => \N__12986\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__22479\
        );

    \uu2.bitmap_RNIKL222_212_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111100"
        )
    port map (
            in0 => \N__10278\,
            in1 => \N__13323\,
            in2 => \N__10296\,
            in3 => \N__10350\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNIKL222Z0Z_212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI9ITA5_3_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__10334\,
            in1 => \N__11463\,
            in2 => \N__10287\,
            in3 => \N__13720\,
            lcout => \uu2.bitmap_pmux_27_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100101"
        )
    port map (
            in0 => \N__13002\,
            in1 => \N__10396\,
            in2 => \N__11133\,
            in3 => \N__11166\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_212_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__11165\,
            in1 => \N__11120\,
            in2 => \N__10401\,
            in3 => \N__13001\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_84_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000111101"
        )
    port map (
            in0 => \N__13004\,
            in1 => \N__10398\,
            in2 => \N__11135\,
            in3 => \N__11168\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_180_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__11164\,
            in1 => \N__11119\,
            in2 => \N__10400\,
            in3 => \N__13000\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_52_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101101101"
        )
    port map (
            in0 => \N__13003\,
            in1 => \N__10397\,
            in2 => \N__11134\,
            in3 => \N__11167\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_RNIU2IS_52_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13804\,
            in1 => \N__10413\,
            in2 => \_gnd_net_\,
            in3 => \N__10407\,
            lcout => \uu2.N_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011110011111"
        )
    port map (
            in0 => \N__13005\,
            in1 => \N__10399\,
            in2 => \N__11136\,
            in3 => \N__11169\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__22477\
        );

    \uu2.bitmap_RNIC6I01_84_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001101001111"
        )
    port map (
            in0 => \N__10362\,
            in1 => \N__13321\,
            in2 => \N__13151\,
            in3 => \N__10356\,
            lcout => \uu2.bitmap_pmux_24_i_m2_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAJJL8_8_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__11576\,
            in1 => \N__10493\,
            in2 => \N__11733\,
            in3 => \N__13441\,
            lcout => \uu2.un51_w_data_displaying\,
            ltout => \uu2.un51_w_data_displaying_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__10803\,
            in1 => \_gnd_net_\,
            in2 => \N__10344\,
            in3 => \N__11699\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11992\,
            in2 => \_gnd_net_\,
            in3 => \N__13115\,
            lcout => \uu2.w_addr_displaying_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000111010"
        )
    port map (
            in0 => \N__10659\,
            in1 => \N__10317\,
            in2 => \N__11717\,
            in3 => \N__10421\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI25P31_0_1_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13818\,
            in1 => \N__11997\,
            in2 => \_gnd_net_\,
            in3 => \N__13117\,
            lcout => \uu2.un49_w_data_displaying_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000101110"
        )
    port map (
            in0 => \N__12132\,
            in1 => \N__11700\,
            in2 => \N__10845\,
            in3 => \N__10422\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI25P31_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13817\,
            in1 => \N__11996\,
            in2 => \_gnd_net_\,
            in3 => \N__13116\,
            lcout => \uu2.un31_w_data_displaying_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIASLS1_1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13118\,
            in1 => \N__11575\,
            in2 => \N__12012\,
            in3 => \N__13816\,
            lcout => \uu2.un31_w_data_displaying_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8NSO_4_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13494\,
            in2 => \_gnd_net_\,
            in3 => \N__11988\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIOELE1_4_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100100110110"
        )
    port map (
            in0 => \N__13160\,
            in1 => \N__11888\,
            in2 => \N__13502\,
            in3 => \N__13707\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI6RE03_3_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100100100"
        )
    port map (
            in0 => \N__13709\,
            in1 => \N__11599\,
            in2 => \N__10440\,
            in3 => \N__13161\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_i5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI1U7M3_7_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010100000"
        )
    port map (
            in0 => \N__13342\,
            in1 => \_gnd_net_\,
            in2 => \N__10437\,
            in3 => \N__13819\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_29_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI30QB21_7_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__11586\,
            in1 => \N__10434\,
            in2 => \N__10425\,
            in3 => \N__10512\,
            lcout => \uu2.bitmap_pmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNICAPH1_2_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13159\,
            in1 => \N__11889\,
            in2 => \N__12011\,
            in3 => \N__13708\,
            lcout => \uu2.un15_w_data_displaying_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__11445\,
            in1 => \N__11412\,
            in2 => \N__11370\,
            in3 => \N__11325\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__22475\
        );

    \uu2.bitmap_RNI1PH82_40_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__10524\,
            in1 => \N__13740\,
            in2 => \N__11496\,
            in3 => \N__13710\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNI1PH82Z0Z_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI208E6_40_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12033\,
            in2 => \N__10518\,
            in3 => \N__12024\,
            lcout => OPEN,
            ltout => \uu2.N_401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIKE7JD_4_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11622\,
            in2 => \N__10515\,
            in3 => \N__12039\,
            lcout => \uu2.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__15988\,
            in1 => \N__12520\,
            in2 => \N__10710\,
            in3 => \N__12141\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__12519\,
            in1 => \N__10704\,
            in2 => \_gnd_net_\,
            in3 => \N__15989\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNII08G4_1_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111111"
        )
    port map (
            in0 => \N__10506\,
            in1 => \N__13442\,
            in2 => \N__10497\,
            in3 => \N__11580\,
            lcout => \uu2.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11707\,
            in1 => \N__11825\,
            in2 => \_gnd_net_\,
            in3 => \N__13172\,
            lcout => \uu2.mem0.N_81_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11754\,
            in1 => \N__11706\,
            in2 => \_gnd_net_\,
            in3 => \N__12018\,
            lcout => \uu2.mem0.N_80_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__12518\,
            in1 => \N__10708\,
            in2 => \N__16007\,
            in3 => \N__12102\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22803\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10737\,
            in1 => \N__12620\,
            in2 => \N__10596\,
            in3 => \N__10767\,
            lcout => \uu2.mem0.N_72_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_data_0_o2_0_4_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__12618\,
            in1 => \N__12119\,
            in2 => \_gnd_net_\,
            in3 => \N__12726\,
            lcout => \uu2.N_111\,
            ltout => \uu2.N_111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110110011"
        )
    port map (
            in0 => \N__10736\,
            in1 => \N__22860\,
            in2 => \N__10638\,
            in3 => \N__10766\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10765\,
            in1 => \N__12621\,
            in2 => \_gnd_net_\,
            in3 => \N__12124\,
            lcout => OPEN,
            ltout => \uu2.mem0.w_data_i_a2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010111011"
        )
    port map (
            in0 => \N__12729\,
            in1 => \N__10738\,
            in2 => \N__10611\,
            in3 => \N__10837\,
            lcout => \uu2.mem0.N_82_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12123\,
            in2 => \_gnd_net_\,
            in3 => \N__12728\,
            lcout => \uu2.mem0.N_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_a2_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011000"
        )
    port map (
            in0 => \N__12727\,
            in1 => \N__12619\,
            in2 => \N__12128\,
            in3 => \N__10764\,
            lcout => \uu2.N_144\,
            ltout => \uu2.N_144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIU0804_6_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__10587\,
            in1 => \N__10554\,
            in2 => \N__10527\,
            in3 => \N__10735\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110111011"
        )
    port map (
            in0 => \N__12596\,
            in1 => \N__10875\,
            in2 => \N__12517\,
            in3 => \N__13913\,
            lcout => \Lab_UT.dispString.dOut_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10752\,
            in1 => \N__10802\,
            in2 => \N__11543\,
            in3 => \N__10652\,
            lcout => OPEN,
            ltout => \uu2.mem0.w_data_0_a2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000110011"
        )
    port map (
            in0 => \N__10779\,
            in1 => \N__10844\,
            in2 => \N__10818\,
            in3 => \N__10740\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_o2_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10801\,
            in1 => \N__10778\,
            in2 => \N__11542\,
            in3 => \N__10651\,
            lcout => \uu2.N_109\,
            ltout => \uu2.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_i_0_tz_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10751\,
            in2 => \N__10743\,
            in3 => \N__10739\,
            lcout => \uu2.w_addr_i_0_tzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIOG7L_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12569\,
            in1 => \N__12667\,
            in2 => \N__12521\,
            in3 => \N__12712\,
            lcout => \Lab_UT.dispString.dOutP_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12713\,
            in1 => \N__12697\,
            in2 => \N__12507\,
            in3 => \N__12571\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__15994\,
            in1 => \N__14805\,
            in2 => \N__12505\,
            in3 => \N__14033\,
            lcout => \Lab_UT.dispString.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12666\,
            lcout => \Lab_UT.dispString.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111101111"
        )
    port map (
            in0 => \N__12668\,
            in1 => \N__13947\,
            in2 => \N__12506\,
            in3 => \N__12570\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__10866\,
            in1 => \N__10680\,
            in2 => \N__10668\,
            in3 => \N__10665\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__15993\,
            in1 => \N__14841\,
            in2 => \N__12504\,
            in3 => \N__13589\,
            lcout => \Lab_UT.dispString.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_2_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__12574\,
            in1 => \_gnd_net_\,
            in2 => \N__12492\,
            in3 => \N__12687\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22787\,
            ce => 'H',
            sr => \N__22499\
        );

    \Lab_UT.dispString.dOut_RNO_3_3_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12441\,
            in2 => \_gnd_net_\,
            in3 => \N__12572\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110001111"
        )
    port map (
            in0 => \N__12681\,
            in1 => \N__14643\,
            in2 => \N__10869\,
            in3 => \N__14507\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__12685\,
            in1 => \N__12442\,
            in2 => \N__16013\,
            in3 => \N__12575\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22787\,
            ce => 'H',
            sr => \N__22499\
        );

    \Lab_UT.dispString.cnt_1_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12573\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12686\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22787\,
            ce => 'H',
            sr => \N__22499\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__10910\,
            in1 => \N__11081\,
            in2 => \N__10941\,
            in3 => \N__11056\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__11027\,
            in1 => \N__11065\,
            in2 => \N__10860\,
            in3 => \N__10857\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22783\,
            ce => 'H',
            sr => \N__22522\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10856\,
            in2 => \_gnd_net_\,
            in3 => \N__10935\,
            lcout => OPEN,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__11080\,
            in1 => \N__10908\,
            in2 => \N__11091\,
            in3 => \N__12798\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__10909\,
            in1 => \_gnd_net_\,
            in2 => \N__11088\,
            in3 => \N__10936\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__11026\,
            in1 => \N__11064\,
            in2 => \N__11085\,
            in3 => \N__11082\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22783\,
            ce => 'H',
            sr => \N__22522\
        );

    \buart.Z_tx.bitcount_1_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110110"
        )
    port map (
            in0 => \N__11057\,
            in1 => \N__10911\,
            in2 => \N__11031\,
            in3 => \N__10940\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22783\,
            ce => 'H',
            sr => \N__22522\
        );

    \uu2.bitmap_314_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011011"
        )
    port map (
            in0 => \N__11214\,
            in1 => \N__11247\,
            in2 => \N__11290\,
            in3 => \N__13035\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__22485\
        );

    \uu2.bitmap_218_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000101"
        )
    port map (
            in0 => \N__13034\,
            in1 => \N__11277\,
            in2 => \N__11252\,
            in3 => \N__11213\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__22485\
        );

    \uu2.bitmap_90_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000011101"
        )
    port map (
            in0 => \N__11216\,
            in1 => \N__11251\,
            in2 => \N__11291\,
            in3 => \N__13037\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__22485\
        );

    \uu2.bitmap_RNILGG61_90_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__10896\,
            in1 => \N__13170\,
            in2 => \N__10890\,
            in3 => \N__13337\,
            lcout => \uu2.bitmap_pmux_25_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__11212\,
            in1 => \N__11243\,
            in2 => \N__11289\,
            in3 => \N__13033\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__22485\
        );

    \uu2.bitmap_58_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101101101"
        )
    port map (
            in0 => \N__13036\,
            in1 => \N__11281\,
            in2 => \N__11253\,
            in3 => \N__11215\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__22485\
        );

    \uu2.bitmap_RNI7GKQ_58_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13336\,
            in1 => \N__11184\,
            in2 => \_gnd_net_\,
            in3 => \N__11178\,
            lcout => OPEN,
            ltout => \uu2.N_216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIS4UH1_314_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12095\,
            in2 => \N__11172\,
            in3 => \N__13823\,
            lcout => \uu2.bitmap_RNIS4UH1Z0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI41KT3_1_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14948\,
            in1 => \N__17928\,
            in2 => \N__15572\,
            in3 => \N__15024\,
            lcout => \Lab_UT.sec1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI63KT3_2_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15026\,
            in1 => \N__17515\,
            in2 => \N__15524\,
            in3 => \N__14950\,
            lcout => \Lab_UT.sec1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNI49824_0_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__13912\,
            in1 => \N__15025\,
            in2 => \N__14962\,
            in3 => \N__15860\,
            lcout => \Lab_UT.min2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNI6B824_1_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15021\,
            in1 => \N__15903\,
            in2 => \N__14603\,
            in3 => \N__14949\,
            lcout => \Lab_UT.min2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNI8D824_2_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14951\,
            in1 => \N__15824\,
            in2 => \N__14388\,
            in3 => \N__15023\,
            lcout => \Lab_UT.min2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNIAF824_3_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__15022\,
            in1 => \N__15726\,
            in2 => \N__14508\,
            in3 => \N__14952\,
            lcout => \Lab_UT.min2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__11316\,
            in1 => \N__11353\,
            in2 => \N__11407\,
            in3 => \N__11436\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_200_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__11434\,
            in1 => \N__11392\,
            in2 => \N__11362\,
            in3 => \N__11314\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_72_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__11317\,
            in1 => \N__11354\,
            in2 => \N__11408\,
            in3 => \N__11437\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_RNIC4D61_72_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__13119\,
            in2 => \N__11475\,
            in3 => \N__13322\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_24_i_m2_bm_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI1UT12_75_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__13120\,
            in1 => \N__11451\,
            in2 => \N__11466\,
            in3 => \N__11457\,
            lcout => \uu2.bitmap_RNI1UT12Z0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__11438\,
            in1 => \N__11402\,
            in2 => \N__11363\,
            in3 => \N__11318\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_203_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__11315\,
            in1 => \N__11352\,
            in2 => \N__11406\,
            in3 => \N__11435\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_168_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__11433\,
            in1 => \N__11391\,
            in2 => \N__11361\,
            in3 => \N__11313\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__22483\
        );

    \uu2.bitmap_69_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011110011111"
        )
    port map (
            in0 => \N__14567\,
            in1 => \N__14538\,
            in2 => \N__13870\,
            in3 => \N__14875\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.bitmap_197_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__14537\,
            in1 => \N__13857\,
            in2 => \N__14887\,
            in3 => \N__14568\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.bitmap_RNI10J51_69_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000111111"
        )
    port map (
            in0 => \N__11562\,
            in1 => \N__13113\,
            in2 => \N__11556\,
            in3 => \N__13319\,
            lcout => \uu2.bitmap_pmux_25_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un437_ci_0_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__13477\,
            in2 => \_gnd_net_\,
            in3 => \N__13384\,
            lcout => OPEN,
            ltout => \uu2.un437_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12962\,
            in1 => \N__11920\,
            in2 => \N__11547\,
            in3 => \N__13320\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.w_addr_displaying_4_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__11924\,
            in1 => \N__12960\,
            in2 => \_gnd_net_\,
            in3 => \N__13478\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.w_addr_displaying_5_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12961\,
            in1 => \N__13385\,
            in2 => \N__13493\,
            in3 => \N__11925\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.w_addr_displaying_0_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__13114\,
            in1 => \_gnd_net_\,
            in2 => \N__11930\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_69C_net\,
            ce => 'H',
            sr => \N__22480\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__11705\,
            in1 => \N__11544\,
            in2 => \_gnd_net_\,
            in3 => \N__11732\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_8_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13812\,
            in1 => \N__13420\,
            in2 => \N__11931\,
            in3 => \N__12941\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_8C_net\,
            ce => 'H',
            sr => \N__22478\
        );

    \uu2.w_addr_displaying_RNIQN495_8_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100111111"
        )
    port map (
            in0 => \N__12939\,
            in1 => \N__11502\,
            in2 => \N__13431\,
            in3 => \N__13810\,
            lcout => \uu2.un33_w_data_displaying\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0ES07_8_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__13811\,
            in1 => \N__12940\,
            in2 => \N__13443\,
            in3 => \N__11704\,
            lcout => \uu2.un21_w_addr_displaying_i\,
            ltout => \uu2.un21_w_addr_displaying_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI47N27_8_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11625\,
            in3 => \N__22557\,
            lcout => \uu2.un21_w_addr_displaying_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIS6T61_1_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__11987\,
            in1 => \N__13702\,
            in2 => \_gnd_net_\,
            in3 => \N__13809\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_3_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13168\,
            in1 => \N__11887\,
            in2 => \N__12013\,
            in3 => \N__13706\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__13548\,
            sr => \N__22476\
        );

    \uu2.w_addr_displaying_nesr_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12000\,
            in2 => \_gnd_net_\,
            in3 => \N__13169\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__13548\,
            sr => \N__22476\
        );

    \uu2.w_addr_displaying_RNIGEPH1_4_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011000000"
        )
    port map (
            in0 => \N__13704\,
            in1 => \N__13498\,
            in2 => \N__11894\,
            in3 => \N__11998\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIUNPV1_2_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001101101100"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__11886\,
            in2 => \N__11604\,
            in3 => \N__13705\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIOM1S6_2_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010100000"
        )
    port map (
            in0 => \N__13212\,
            in1 => \N__11616\,
            in2 => \N__11607\,
            in3 => \N__11603\,
            lcout => \uu2.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI8NSO_2_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11882\,
            in2 => \_gnd_net_\,
            in3 => \N__13703\,
            lcout => \uu2.un15_w_data_displaying_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIVKR41_180_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13696\,
            in1 => \N__12096\,
            in2 => \_gnd_net_\,
            in3 => \N__12081\,
            lcout => OPEN,
            ltout => \uu2.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIAKAQ2_7_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__13701\,
            in1 => \N__13338\,
            in2 => \N__12072\,
            in3 => \N__12069\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI206J5_7_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12060\,
            in2 => \N__12051\,
            in3 => \N__12048\,
            lcout => \uu2.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIJHPH1_2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001110"
        )
    port map (
            in0 => \N__11860\,
            in1 => \N__13698\,
            in2 => \N__13346\,
            in3 => \N__11986\,
            lcout => \uu2.bitmap_pmux_sn_N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIM0T61_2_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000101"
        )
    port map (
            in0 => \N__13697\,
            in1 => \_gnd_net_\,
            in2 => \N__12010\,
            in3 => \N__11859\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIELSJ2_111_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__13614\,
            in1 => \_gnd_net_\,
            in2 => \N__12027\,
            in3 => \N__12213\,
            lcout => \uu2.bitmap_RNIELSJ2Z0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__11881\,
            in1 => \N__12017\,
            in2 => \N__13176\,
            in3 => \N__11929\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \uu2.w_addr_user_1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001011110000"
        )
    port map (
            in0 => \N__11826\,
            in1 => \N__12315\,
            in2 => \N__11768\,
            in3 => \N__12376\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \uu2.w_addr_user_4_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011010010"
        )
    port map (
            in0 => \N__12377\,
            in1 => \N__12360\,
            in2 => \N__12280\,
            in3 => \N__12316\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \uu2.bitmap_111_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12243\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \uu2.vram_rd_clk_det_0_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \uu2.vram_rd_clk_det_1_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12170\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2C_net\,
            ce => 'H',
            sr => \N__22474\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010111"
        )
    port map (
            in0 => \N__12511\,
            in1 => \N__12600\,
            in2 => \N__12698\,
            in3 => \N__14047\,
            lcout => \Lab_UT.dispString.dOutP_1_iv_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101000101"
        )
    port map (
            in0 => \N__12603\,
            in1 => \N__12714\,
            in2 => \N__12525\,
            in3 => \N__15573\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12694\,
            in2 => \N__12135\,
            in3 => \N__12384\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22795\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_5_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101111111"
        )
    port map (
            in0 => \N__12512\,
            in1 => \N__12601\,
            in2 => \N__12699\,
            in3 => \N__14048\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__16008\,
            in1 => \N__14732\,
            in2 => \N__12524\,
            in3 => \N__13991\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001111"
        )
    port map (
            in0 => \N__14379\,
            in1 => \N__12513\,
            in2 => \N__12741\,
            in3 => \N__12602\,
            lcout => \Lab_UT.dispString.dOut_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100011111"
        )
    port map (
            in0 => \N__12598\,
            in1 => \N__14159\,
            in2 => \N__12523\,
            in3 => \N__14682\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__12695\,
            in1 => \_gnd_net_\,
            in2 => \N__12738\,
            in3 => \N__12735\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI_1_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14221\,
            in2 => \_gnd_net_\,
            in3 => \N__14189\,
            lcout => \Lab_UT.alarmchar_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000111111"
        )
    port map (
            in0 => \N__14160\,
            in1 => \N__12599\,
            in2 => \N__15528\,
            in3 => \N__12502\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12696\,
            in2 => \N__12630\,
            in3 => \N__12627\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100010001"
        )
    port map (
            in0 => \N__12597\,
            in1 => \N__12531\,
            in2 => \N__12522\,
            in3 => \N__14607\,
            lcout => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18666\,
            in2 => \_gnd_net_\,
            in3 => \N__17563\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m1_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18667\,
            in2 => \_gnd_net_\,
            in3 => \N__17564\,
            lcout => \Lab_UT.dictrl.alarmstate8_2_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18669\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22788\,
            ce => \N__15606\,
            sr => \N__22520\
        );

    \Lab_UT.dictrl.shifter_ret_1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18668\,
            in2 => \_gnd_net_\,
            in3 => \N__17565\,
            lcout => \Lab_UT.dictrl.alarmstate8_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22788\,
            ce => \N__15606\,
            sr => \N__22520\
        );

    \buart.Z_rx.shifter_0_3_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21063\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22788\,
            ce => \N__15606\,
            sr => \N__22520\
        );

    \buart.Z_rx.shifter_ret_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17566\,
            lcout => bu_rx_data_i_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22788\,
            ce => \N__15606\,
            sr => \N__22520\
        );

    \buart.Z_rx.shifter_ret_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20799\,
            lcout => bu_rx_data_i_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22784\,
            ce => \N__15604\,
            sr => \N__22523\
        );

    \resetGen.escKey_4_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21069\,
            in1 => \N__18154\,
            in2 => \N__20833\,
            in3 => \N__18695\,
            lcout => \resetGen.escKeyZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_6_rep1_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21072\,
            lcout => bu_rx_data_i_4_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__15602\,
            sr => \N__22525\
        );

    \buart.Z_rx.shifter_ret_6_fast_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21071\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_4_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__15602\,
            sr => \N__22525\
        );

    \buart.Z_rx.shifter_0_fast_3_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21073\,
            lcout => \buart__rx_shifter_0_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__15602\,
            sr => \N__22525\
        );

    \buart.Z_rx.shifter_ret_6_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__21070\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__15602\,
            sr => \N__22525\
        );

    \buart.Z_rx.shifter_0_1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17596\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22779\,
            ce => \N__15602\,
            sr => \N__22525\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12887\,
            in1 => \N__12821\,
            in2 => \N__12860\,
            in3 => \N__12912\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12891\,
            in2 => \N__12864\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12924\,
            in3 => \N__12825\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__22776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12800\,
            in1 => \N__12822\,
            in2 => \_gnd_net_\,
            in3 => \N__12810\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__22776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12768\,
            in3 => \N__12807\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__22776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__12801\,
            in1 => \_gnd_net_\,
            in2 => \N__12780\,
            in3 => \N__12804\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__22776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__12755\,
            in1 => \N__12799\,
            in2 => \_gnd_net_\,
            in3 => \N__12783\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22776\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12776\,
            in1 => \N__12764\,
            in2 => \N__12756\,
            in3 => \N__12920\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNICJDT_1_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__15377\,
            in1 => \N__14023\,
            in2 => \N__13987\,
            in3 => \N__15457\,
            lcout => \Lab_UT.didp.did_alarmMatch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14459\,
            in3 => \N__15378\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17834\,
            in1 => \N__18729\,
            in2 => \N__12906\,
            in3 => \N__15428\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__15930\,
            in1 => \N__15429\,
            in2 => \N__12903\,
            in3 => \N__14445\,
            lcout => \Lab_UT.didp.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__15394\,
            in1 => \N__17833\,
            in2 => \N__14460\,
            in3 => \N__17634\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__14444\,
            in1 => \N__15929\,
            in2 => \N__12900\,
            in3 => \N__15395\,
            lcout => \Lab_UT.didp.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22835\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000001"
        )
    port map (
            in0 => \N__15776\,
            in1 => \N__16248\,
            in2 => \N__16281\,
            in3 => \N__12897\,
            lcout => \Lab_UT.didp.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__15858\,
            in1 => \N__15772\,
            in2 => \_gnd_net_\,
            in3 => \N__18214\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNINAVN_0_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13911\,
            in2 => \_gnd_net_\,
            in3 => \N__15857\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.un2_did_alarmMatch_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNIOMK62_0_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__15227\,
            in1 => \N__14834\,
            in2 => \N__13047\,
            in3 => \N__12969\,
            lcout => \Lab_UT.didp.regrce4.did_alarmMatch_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_1_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20886\,
            in1 => \N__15902\,
            in2 => \N__15786\,
            in3 => \N__15859\,
            lcout => \Lab_UT.didp.countrce3.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNI0LVO3_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14944\,
            in1 => \N__17795\,
            in2 => \N__15048\,
            in3 => \N__13588\,
            lcout => \Lab_UT.sec2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNIR0LH1_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__16764\,
            in1 => \N__20345\,
            in2 => \N__18024\,
            in3 => \N__16547\,
            lcout => \Lab_UT.loadalarm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_RNIITJO1_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110111"
        )
    port map (
            in0 => \N__22242\,
            in1 => \N__14770\,
            in2 => \N__20368\,
            in3 => \N__16765\,
            lcout => \Lab_UT.loadalarm_0_0\,
            ltout => \Lab_UT.loadalarm_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_RNI2VJT3_0_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__14664\,
            in1 => \N__17472\,
            in2 => \N__13008\,
            in3 => \N__15030\,
            lcout => \Lab_UT.sec1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_RNI8N121_0_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__13587\,
            in1 => \N__17471\,
            in2 => \N__14671\,
            in3 => \N__17794\,
            lcout => \Lab_UT.didp.did_alarmMatch_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNIANSM3_2_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14960\,
            in1 => \N__14423\,
            in2 => \N__14733\,
            in3 => \N__15031\,
            lcout => \Lab_UT.min1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_6_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__13380\,
            in1 => \N__13246\,
            in2 => \N__12963\,
            in3 => \N__13476\,
            lcout => OPEN,
            ltout => \uu2.o_adder_vbuf_w_addr_displaying_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_6_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011110000"
        )
    port map (
            in0 => \N__13815\,
            in1 => \_gnd_net_\,
            in2 => \N__13551\,
            in3 => \N__13424\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_ness_6C_net\,
            ce => \N__13547\,
            sr => \N__22484\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__13377\,
            in1 => \N__13311\,
            in2 => \N__13251\,
            in3 => \N__13813\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13312\,
            in1 => \N__13475\,
            in2 => \N__13253\,
            in3 => \N__13378\,
            lcout => \uu2.un15_w_data_displaying_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__13379\,
            in1 => \N__13313\,
            in2 => \N__13252\,
            in3 => \N__13814\,
            lcout => \uu2.bitmap_pmux_sn_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_290_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011011"
        )
    port map (
            in0 => \N__14533\,
            in1 => \N__13862\,
            in2 => \N__14900\,
            in3 => \N__14565\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__22481\
        );

    \uu2.bitmap_194_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000101"
        )
    port map (
            in0 => \N__14562\,
            in1 => \N__14888\,
            in2 => \N__13871\,
            in3 => \N__14535\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__22481\
        );

    \uu2.bitmap_66_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000011101"
        )
    port map (
            in0 => \N__14534\,
            in1 => \N__13863\,
            in2 => \N__14901\,
            in3 => \N__14566\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__22481\
        );

    \uu2.bitmap_RNIV8902_66_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111100010"
        )
    port map (
            in0 => \N__13200\,
            in1 => \N__13194\,
            in2 => \N__13188\,
            in3 => \N__13150\,
            lcout => \uu2.bitmap_RNIV8902Z0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__14532\,
            in1 => \N__13861\,
            in2 => \N__14899\,
            in3 => \N__14564\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__22481\
        );

    \uu2.bitmap_34_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011101101101"
        )
    port map (
            in0 => \N__14563\,
            in1 => \N__14889\,
            in2 => \N__13872\,
            in3 => \N__14536\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__22481\
        );

    \uu2.bitmap_RNIEJM91_34_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__13833\,
            in1 => \N__13805\,
            in2 => \N__13749\,
            in3 => \N__13700\,
            lcout => \uu2.bitmap_pmux_26_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI6RO21_162_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__13699\,
            in1 => \N__13629\,
            in2 => \_gnd_net_\,
            in3 => \N__13620\,
            lcout => \uu2.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14690\,
            in2 => \_gnd_net_\,
            in3 => \N__14413\,
            lcout => \Lab_UT.didp.countrce4.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNIOF7P_1_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__16159\,
            in1 => \N__14715\,
            in2 => \N__14422\,
            in3 => \N__14793\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNIGCKQ8_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15099\,
            in1 => \N__14343\,
            in2 => \N__13605\,
            in3 => \N__13602\,
            lcout => \Lab_UT.alarmMatch\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__14414\,
            in1 => \N__15173\,
            in2 => \N__14694\,
            in3 => \N__17620\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__16086\,
            in1 => \N__15141\,
            in2 => \N__13593\,
            in3 => \N__14415\,
            lcout => \Lab_UT.didp.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22800\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_0_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__18200\,
            in1 => \N__16548\,
            in2 => \N__13590\,
            in3 => \N__16436\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce1.q_1_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16549\,
            in1 => \N__20878\,
            in2 => \N__16450\,
            in3 => \N__14022\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce1.q_2_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17615\,
            in1 => \N__16550\,
            in2 => \N__13986\,
            in3 => \N__16440\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce1.q_3_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16551\,
            in1 => \N__18718\,
            in2 => \N__16451\,
            in3 => \N__13936\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce3.q_0_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__18201\,
            in1 => \N__16762\,
            in2 => \N__13914\,
            in3 => \N__16444\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce3.q_3_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16761\,
            in1 => \N__18719\,
            in2 => \N__16452\,
            in3 => \N__14493\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.didp.regrce3.q_2_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17616\,
            in1 => \N__16763\,
            in2 => \N__14387\,
            in3 => \N__16445\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22796\,
            ce => 'H',
            sr => \N__22498\
        );

    \Lab_UT.dictrl.g0_9_1_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18707\,
            in2 => \_gnd_net_\,
            in3 => \N__17600\,
            lcout => \Lab_UT.dictrl.g0_9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIR2IE1_2_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20175\,
            in1 => \N__16993\,
            in2 => \_gnd_net_\,
            in3 => \N__21386\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19645\,
            in1 => \N__14185\,
            in2 => \_gnd_net_\,
            in3 => \N__14214\,
            lcout => \Lab_UT.dictrl.alarmstate_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNIMIM09_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000100110"
        )
    port map (
            in0 => \N__14186\,
            in1 => \N__14112\,
            in2 => \N__14223\,
            in3 => \N__14148\,
            lcout => \Lab_UT.dictrl.alarmstate_1_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNIGCKQ8_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111000001100"
        )
    port map (
            in0 => \N__14147\,
            in1 => \N__14219\,
            in2 => \N__14058\,
            in3 => \N__14188\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNIK5FS8_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__14220\,
            in1 => \N__14085\,
            in2 => \N__14097\,
            in3 => \N__14091\,
            lcout => \Lab_UT.shifter_ret_3_RNIK5FS8_0\,
            ltout => \Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111111"
        )
    port map (
            in0 => \N__19644\,
            in1 => \_gnd_net_\,
            in2 => \N__14094\,
            in3 => \N__14184\,
            lcout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i\,
            ltout => \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNIQBH29_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__14187\,
            in1 => \N__14084\,
            in2 => \N__14076\,
            in3 => \N__14073\,
            lcout => \Lab_UT.shifter_ret_3_RNIQBH29_0\,
            ltout => \Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI_2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14067\,
            in3 => \N__14218\,
            lcout => \Lab_UT.trig\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI6H8A1_2_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21387\,
            in1 => \N__16449\,
            in2 => \_gnd_net_\,
            in3 => \N__20176\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__20359\,
            in1 => \N__14256\,
            in2 => \N__14247\,
            in3 => \N__14064\,
            lcout => \Lab_UT.dictrl.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI6626_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14108\,
            in2 => \_gnd_net_\,
            in3 => \N__14231\,
            lcout => \Lab_UT.dictrl.N_127_0_0\,
            ltout => \Lab_UT.dictrl.N_127_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNI_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100010"
        )
    port map (
            in0 => \N__14232\,
            in1 => \N__14049\,
            in2 => \N__14235\,
            in3 => \N__14127\,
            lcout => \Lab_UT.dictrl.justentered_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m9_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14222\,
            in2 => \_gnd_net_\,
            in3 => \N__14190\,
            lcout => \Lab_UT.armed\,
            ltout => \Lab_UT.armed_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14151\,
            in3 => \N__14146\,
            lcout => \G_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_5_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21532\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \buart.Z_rx.shifter_0_7_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19473\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \buart.Z_rx.shifter_0_6_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14271\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \Lab_UT.dictrl.shifter_ret_3_RNO_0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20967\,
            in1 => \N__21062\,
            in2 => \N__14274\,
            in3 => \N__20851\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.alarmstate8_10_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14121\,
            in1 => \N__19472\,
            in2 => \N__14115\,
            in3 => \N__21531\,
            lcout => \Lab_UT.dictrl.alarmstate8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \buart.Z_rx.shifter_0_4_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20968\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \buart.Z_rx.shifter_0_fast_6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14273\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \buart.Z_rx.shifter_0_6_rep1_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22781\,
            ce => \N__15605\,
            sr => \N__22524\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__21530\,
            in1 => \N__20962\,
            in2 => \N__22269\,
            in3 => \N__21385\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_5_fast_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20964\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_ret_5_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22778\,
            ce => \N__15603\,
            sr => \N__22526\
        );

    \buart.Z_rx.shifter_0_fast_4_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20966\,
            lcout => bu_rx_data_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22778\,
            ce => \N__15603\,
            sr => \N__22526\
        );

    \buart.Z_rx.shifter_ret_5_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20963\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22778\,
            ce => \N__15603\,
            sr => \N__22526\
        );

    \buart.Z_rx.shifter_0_4_rep1_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20965\,
            lcout => bu_rx_data_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22778\,
            ce => \N__15603\,
            sr => \N__22526\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21656\,
            in1 => \N__21430\,
            in2 => \N__17078\,
            in3 => \N__21698\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_0_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20800\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22778\,
            ce => \N__15603\,
            sr => \N__22526\
        );

    \Lab_UT.dictrl.g0_31_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__17380\,
            in1 => \N__17192\,
            in2 => \N__17277\,
            in3 => \N__17342\,
            lcout => \Lab_UT.dictrl.N_98_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m40_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17379\,
            in1 => \N__17275\,
            in2 => \N__14313\,
            in3 => \N__17193\,
            lcout => \Lab_UT.dictrl.N_99_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_1_4_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__14319\,
            in1 => \N__17271\,
            in2 => \N__14312\,
            in3 => \N__17378\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_1_RNICGMV1_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__17147\,
            in1 => \N__21544\,
            in2 => \N__14295\,
            in3 => \N__18137\,
            lcout => \Lab_UT.dictrl.g1_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_5_rep1_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21545\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22775\,
            ce => \N__15601\,
            sr => \N__22527\
        );

    \buart.Z_rx.shifter_0_fast_5_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21546\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22775\,
            ce => \N__15601\,
            sr => \N__22527\
        );

    \Lab_UT.dictrl.g0_43_x_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17311\,
            in1 => \N__17270\,
            in2 => \_gnd_net_\,
            in3 => \N__15344\,
            lcout => \Lab_UT.dictrl.g0_43_xZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_15_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15351\,
            in1 => \N__17234\,
            in2 => \N__15642\,
            in3 => \N__17307\,
            lcout => \Lab_UT.dictrl.N_98_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_20_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15677\,
            in1 => \N__15318\,
            in2 => \N__14292\,
            in3 => \N__20779\,
            lcout => \Lab_UT.dictrl.N_88_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_14_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17306\,
            in1 => \N__15350\,
            in2 => \_gnd_net_\,
            in3 => \N__20641\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_11_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20780\,
            in1 => \N__14283\,
            in2 => \N__14277\,
            in3 => \N__15678\,
            lcout => \Lab_UT.dictrl.N_88_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20887\,
            in1 => \N__15462\,
            in2 => \N__17835\,
            in3 => \N__17791\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15463\,
            in1 => \N__15923\,
            in2 => \N__14463\,
            in3 => \N__14443\,
            lcout => \Lab_UT.didp.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNIVHJJ_1_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15461\,
            in2 => \_gnd_net_\,
            in3 => \N__17790\,
            lcout => \Lab_UT.didp.countrce1.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI65GA_0_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14853\,
            in2 => \_gnd_net_\,
            in3 => \N__17709\,
            lcout => \Lab_UT.didp.un1_dicLdSones_0\,
            ltout => \Lab_UT.didp.un1_dicLdSones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__17792\,
            in1 => \N__15922\,
            in2 => \N__14430\,
            in3 => \N__17760\,
            lcout => \Lab_UT.didp.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14427\,
            lcout => \Lab_UT.didp.reset_12_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__15895\,
            in1 => \N__14383\,
            in2 => \N__15823\,
            in3 => \N__14584\,
            lcout => \Lab_UT.didp.did_alarmMatch_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI14UL1_2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__16241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15789\,
            lcout => \Lab_UT.didp.un1_dicLdMones_0\,
            ltout => \Lab_UT.didp.un1_dicLdMones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__15896\,
            in1 => \N__16270\,
            in2 => \N__14331\,
            in3 => \N__14328\,
            lcout => \Lab_UT.didp.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22839\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_0_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__18215\,
            in1 => \N__16768\,
            in2 => \N__14681\,
            in3 => \N__17026\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce2.q_1_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16766\,
            in1 => \N__20876\,
            in2 => \N__17036\,
            in3 => \N__15558\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce2.q_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17635\,
            in1 => \N__16769\,
            in2 => \N__15516\,
            in3 => \N__17030\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce2.q_3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__16767\,
            in1 => \N__18740\,
            in2 => \N__17037\,
            in3 => \N__14626\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce3.q_1_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__20875\,
            in1 => \N__16770\,
            in2 => \N__16417\,
            in3 => \N__14590\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce4.q_3_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__17025\,
            in1 => \N__14771\,
            in2 => \N__15089\,
            in3 => \N__18741\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22504\
        );

    \Lab_UT.didp.regrce4.q_RNI6JSM3_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__15225\,
            in1 => \N__14953\,
            in2 => \N__15049\,
            in3 => \N__14829\,
            lcout => \Lab_UT.min1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNI8LSM3_1_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14954\,
            in1 => \N__16171\,
            in2 => \N__15050\,
            in3 => \N__14794\,
            lcout => \Lab_UT.min1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNISBJ41_3_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__14503\,
            in1 => \N__15725\,
            in2 => \N__16129\,
            in3 => \N__15078\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNICAPA4_3_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15477\,
            in1 => \N__15126\,
            in2 => \N__15114\,
            in3 => \N__15111\,
            lcout => \Lab_UT.didp.regrce4.did_alarmMatch_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_RNICPSM3_3_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15079\,
            in1 => \N__15035\,
            in2 => \N__16130\,
            in3 => \N__14961\,
            lcout => \Lab_UT.min1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__14763\,
            in1 => \N__17722\,
            in2 => \N__22596\,
            in3 => \N__19947\,
            lcout => \Lab_UT.dicRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22819\,
            ce => 'H',
            sr => \N__22501\
        );

    \Lab_UT.didp.ce_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16012\,
            in1 => \N__14766\,
            in2 => \_gnd_net_\,
            in3 => \N__16407\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22819\,
            ce => 'H',
            sr => \N__22501\
        );

    \Lab_UT.didp.regrce4.q_0_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14764\,
            in1 => \N__18226\,
            in2 => \N__17034\,
            in3 => \N__14833\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22819\,
            ce => 'H',
            sr => \N__22501\
        );

    \Lab_UT.didp.regrce4.q_1_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__14798\,
            in1 => \N__20877\,
            in2 => \N__14772\,
            in3 => \N__17021\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22819\,
            ce => 'H',
            sr => \N__22501\
        );

    \Lab_UT.didp.regrce4.q_2_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14765\,
            in1 => \N__17633\,
            in2 => \N__17035\,
            in3 => \N__14722\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22819\,
            ce => 'H',
            sr => \N__22501\
        );

    \Lab_UT.didp.countrce4.q_RNI5GGH_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15214\,
            in2 => \_gnd_net_\,
            in3 => \N__16163\,
            lcout => \Lab_UT.didp.countrce4.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__15215\,
            in1 => \N__15170\,
            in2 => \_gnd_net_\,
            in3 => \N__18225\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100001"
        )
    port map (
            in0 => \N__15696\,
            in1 => \N__15174\,
            in2 => \N__15231\,
            in3 => \N__16080\,
            lcout => \Lab_UT.didp.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__16164\,
            in1 => \N__15171\,
            in2 => \N__15226\,
            in3 => \N__20888\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__16175\,
            in1 => \N__15139\,
            in2 => \N__15186\,
            in3 => \N__16081\,
            lcout => \Lab_UT.didp.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__18720\,
            in2 => \N__16128\,
            in3 => \N__15172\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__16118\,
            in1 => \N__16082\,
            in2 => \N__15177\,
            in3 => \N__15140\,
            lcout => \Lab_UT.didp.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22812\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNIDJKH1_3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15695\,
            in2 => \_gnd_net_\,
            in3 => \N__15169\,
            lcout => \Lab_UT.didp.un1_dicLdMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16481\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22804\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIE8RP4_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19889\,
            in1 => \N__16881\,
            in2 => \_gnd_net_\,
            in3 => \N__22093\,
            lcout => \Lab_UT.dictrl.N_121_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_0_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18882\,
            in1 => \N__19888\,
            in2 => \_gnd_net_\,
            in3 => \N__21120\,
            lcout => \Lab_UT.dictrl.g1_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__21121\,
            in1 => \_gnd_net_\,
            in2 => \N__19901\,
            in3 => \N__18883\,
            lcout => \Lab_UT.dictrl.g3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_27_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18536\,
            in1 => \N__16837\,
            in2 => \N__18223\,
            in3 => \N__18076\,
            lcout => \Lab_UT.dictrl.N_116_mux_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18077\,
            in1 => \N__16848\,
            in2 => \N__18224\,
            in3 => \N__18537\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_116_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI4N0L4_3_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011101"
        )
    port map (
            in0 => \N__20352\,
            in1 => \N__22201\,
            in2 => \N__15249\,
            in3 => \N__21359\,
            lcout => \Lab_UT.dictrl.N_1304_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNI24TF4_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101110011"
        )
    port map (
            in0 => \N__21357\,
            in1 => \N__20351\,
            in2 => \N__21146\,
            in3 => \N__15246\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1304_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIQ1339_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__22199\,
            in1 => \N__22095\,
            in2 => \N__15240\,
            in3 => \N__21358\,
            lcout => \Lab_UT.dictrl.N_94_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNISK689_0_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__22096\,
            in1 => \N__15237\,
            in2 => \N__21383\,
            in3 => \N__22200\,
            lcout => \Lab_UT.dictrl.N_94_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0_3_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101001111"
        )
    port map (
            in0 => \N__21366\,
            in1 => \N__22262\,
            in2 => \N__20370\,
            in3 => \N__20469\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__20879\,
            in1 => \N__21363\,
            in2 => \N__22268\,
            in3 => \N__20656\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNICSUJ_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19883\,
            in2 => \_gnd_net_\,
            in3 => \N__21149\,
            lcout => \Lab_UT.dicLdMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_7_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010011"
        )
    port map (
            in0 => \N__20468\,
            in1 => \N__18288\,
            in2 => \N__21158\,
            in3 => \N__21364\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1304_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_5_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__21365\,
            in1 => \N__21153\,
            in2 => \N__15273\,
            in3 => \N__22094\,
            lcout => \Lab_UT.dictrl.N_94_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIBHFL_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21355\,
            lcout => \Lab_UT.dictrl.m36_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIAUDM_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18286\,
            in2 => \_gnd_net_\,
            in3 => \N__21722\,
            lcout => \Lab_UT.dictrl.m45_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__17112\,
            in1 => \N__18854\,
            in2 => \_gnd_net_\,
            in3 => \N__18287\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_8_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__15270\,
            in1 => \N__15255\,
            in2 => \N__15258\,
            in3 => \N__21356\,
            lcout => \Lab_UT.dictrl.i9_mux_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_9_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17049\,
            in1 => \N__15651\,
            in2 => \_gnd_net_\,
            in3 => \N__16828\,
            lcout => \Lab_UT.dictrl.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m25_4_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__21699\,
            in1 => \N__17176\,
            in2 => \N__21431\,
            in3 => \N__15640\,
            lcout => \Lab_UT.dictrl.m25Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m25_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16943\,
            in1 => \_gnd_net_\,
            in2 => \N__17428\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.m25Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_fast_RNI13PI1_2_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__18136\,
            in1 => \N__17420\,
            in2 => \N__18544\,
            in3 => \N__16944\,
            lcout => g0_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m25_x1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16942\,
            in1 => \N__18532\,
            in2 => \N__17427\,
            in3 => \N__18135\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m25_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m25_ns_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15294\,
            in3 => \N__18067\,
            lcout => \Lab_UT.dictrl.N_116_mux\,
            ltout => \Lab_UT.dictrl.N_116_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNIB8OC4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__19882\,
            in1 => \N__17973\,
            in2 => \N__15291\,
            in3 => \N__21354\,
            lcout => \Lab_UT.dictrl.N_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_11_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20946\,
            in1 => \N__21037\,
            in2 => \N__21540\,
            in3 => \N__21630\,
            lcout => \Lab_UT.dictrl.N_98_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_1_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20637\,
            in1 => \N__20945\,
            in2 => \_gnd_net_\,
            in3 => \N__21038\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_35_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__20856\,
            in1 => \N__15680\,
            in2 => \N__15288\,
            in3 => \N__18561\,
            lcout => \Lab_UT.dictrl.g1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15285\,
            in1 => \N__20371\,
            in2 => \N__18576\,
            in3 => \N__21502\,
            lcout => \Lab_UT.dictrl.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_46_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20944\,
            in1 => \N__21036\,
            in2 => \N__21539\,
            in3 => \N__21629\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_98_mux_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_42_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__15357\,
            in1 => \N__15681\,
            in2 => \N__15276\,
            in3 => \N__20857\,
            lcout => \Lab_UT.dictrl.g1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_1_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20943\,
            in1 => \N__21035\,
            in2 => \_gnd_net_\,
            in3 => \N__20636\,
            lcout => \Lab_UT.dictrl.g1_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_2_1_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21631\,
            in1 => \N__20947\,
            in2 => \N__21560\,
            in3 => \N__21039\,
            lcout => \Lab_UT.dictrl.g1_2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_28_1_0_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100110011"
        )
    port map (
            in0 => \N__17336\,
            in1 => \N__15343\,
            in2 => \N__15312\,
            in3 => \N__20801\,
            lcout => \Lab_UT.dictrl.g0_28_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_3_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15311\,
            in1 => \N__17377\,
            in2 => \_gnd_net_\,
            in3 => \N__17338\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__15327\,
            in1 => \N__15679\,
            in2 => \N__15321\,
            in3 => \N__20802\,
            lcout => \Lab_UT.dictrl.N_88_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_4_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15310\,
            in1 => \N__17376\,
            in2 => \_gnd_net_\,
            in3 => \N__17337\,
            lcout => \Lab_UT.dictrl.g0_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_1_fast_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18716\,
            lcout => \buart__rx_shifter_ret_1_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22780\,
            ce => \N__15600\,
            sr => \N__22529\
        );

    \buart.Z_rx.shifter_0_fast_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart__rx_shifter_0_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22780\,
            ce => \N__15600\,
            sr => \N__22529\
        );

    \buart.Z_rx.shifter_ret_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18715\,
            lcout => bu_rx_data_i_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22780\,
            ce => \N__15600\,
            sr => \N__22529\
        );

    \Lab_UT.dictrl.m31_x0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20632\,
            in1 => \N__17375\,
            in2 => \N__15641\,
            in3 => \N__17335\,
            lcout => \Lab_UT.dictrl.m31_xZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m19_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17232\,
            in2 => \_gnd_net_\,
            in3 => \N__15635\,
            lcout => \Lab_UT.dictrl.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_12_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15636\,
            in1 => \N__17233\,
            in2 => \N__17312\,
            in3 => \N__21436\,
            lcout => \Lab_UT.dictrl.g0_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_3_fast_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19470\,
            lcout => bu_rx_data_i_4_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22777\,
            ce => \N__15599\,
            sr => \N__22531\
        );

    \buart.Z_rx.shifter_ret_3_rep1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19471\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_i_4_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22777\,
            ce => \N__15599\,
            sr => \N__22531\
        );

    \buart.Z_rx.shifter_ret_3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19469\,
            lcout => bu_rx_data_i_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22777\,
            ce => \N__15599\,
            sr => \N__22531\
        );

    \buart.Z_rx.shifter_ret_4_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21571\,
            lcout => bu_rx_data_i_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22774\,
            ce => \N__15598\,
            sr => \N__22533\
        );

    \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__17503\,
            in1 => \N__15559\,
            in2 => \N__15517\,
            in3 => \N__17920\,
            lcout => \Lab_UT.didp.did_alarmMatch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15464\,
            in1 => \N__15432\,
            in2 => \N__15396\,
            in3 => \N__17793\,
            lcout => \Lab_UT.didp.un18_ce\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__17921\,
            in1 => \N__17675\,
            in2 => \N__17516\,
            in3 => \N__17470\,
            lcout => \Lab_UT.didp.un24_ce_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__15867\,
            in1 => \N__15901\,
            in2 => \N__15825\,
            in3 => \N__15722\,
            lcout => \Lab_UT.didp.countrce3.ce_12_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNI36SS_0_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15900\,
            in2 => \_gnd_net_\,
            in3 => \N__15866\,
            lcout => \Lab_UT.didp.countrce3.un13_qPone\,
            ltout => \Lab_UT.didp.countrce3.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__15821\,
            in1 => \N__15787\,
            in2 => \N__15837\,
            in3 => \N__17636\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__16280\,
            in1 => \N__15734\,
            in2 => \N__15834\,
            in3 => \N__15822\,
            lcout => \Lab_UT.didp.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15831\,
            in2 => \_gnd_net_\,
            in3 => \N__15820\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__15788\,
            in1 => \N__18739\,
            in2 => \N__15741\,
            in3 => \N__15723\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__15724\,
            in1 => \N__16269\,
            in2 => \N__15738\,
            in3 => \N__15735\,
            lcout => \Lab_UT.didp.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_1_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16057\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.ce_3_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16061\,
            in1 => \N__16229\,
            in2 => \N__16214\,
            in3 => \N__16035\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.reset_2_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16032\,
            in1 => \N__16062\,
            in2 => \N__16215\,
            in3 => \N__16230\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.ce_2_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16058\,
            in1 => \N__16209\,
            in2 => \_gnd_net_\,
            in3 => \N__16034\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.reset_1_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16031\,
            in1 => \N__16205\,
            in2 => \_gnd_net_\,
            in3 => \N__16060\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16056\,
            in1 => \N__16228\,
            in2 => \N__16213\,
            in3 => \N__16029\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__16182\,
            in1 => \N__16176\,
            in2 => \N__16134\,
            in3 => \N__16131\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \Lab_UT.didp.reset_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16033\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22840\,
            ce => 'H',
            sr => \N__22505\
        );

    \resetGen.reset_count_1_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010100"
        )
    port map (
            in0 => \N__18480\,
            in1 => \N__16383\,
            in2 => \N__16368\,
            in3 => \N__16480\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100101"
        )
    port map (
            in0 => \N__16363\,
            in1 => \_gnd_net_\,
            in2 => \N__16482\,
            in3 => \N__18479\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16382\,
            in2 => \_gnd_net_\,
            in3 => \N__16362\,
            lcout => \resetGen.un241_ci\,
            ltout => \resetGen.un241_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011100"
        )
    port map (
            in0 => \N__16478\,
            in1 => \N__16340\,
            in2 => \N__16506\,
            in3 => \N__18481\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__18482\,
            in1 => \N__16479\,
            in2 => \N__16503\,
            in3 => \N__16326\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16499\,
            in2 => \_gnd_net_\,
            in3 => \N__16339\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001000100"
        )
    port map (
            in0 => \N__18483\,
            in1 => \N__16474\,
            in2 => \N__16491\,
            in3 => \N__16488\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNINALF_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20347\,
            lcout => \Lab_UT.dicRun_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__22988\,
            in1 => \N__19404\,
            in2 => \N__19166\,
            in3 => \N__18048\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22823\,
            ce => \N__19349\,
            sr => \N__22528\
        );

    \buart.Z_rx.bitcount_es_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__19403\,
            in1 => \N__22989\,
            in2 => \N__19200\,
            in3 => \N__18039\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22823\,
            ce => \N__19349\,
            sr => \N__22528\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16381\,
            in1 => \N__16367\,
            in2 => \_gnd_net_\,
            in3 => \N__16341\,
            lcout => \resetGen.un252_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_RNILLLG7_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__16320\,
            in1 => \N__16296\,
            in2 => \_gnd_net_\,
            in3 => \N__16644\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIQ3CG_2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__21951\,
            in3 => \N__20129\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIJT2J_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20095\,
            lcout => \Lab_UT.dicLdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUQEL8_1_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__16698\,
            in1 => \N__16683\,
            in2 => \N__16521\,
            in3 => \N__21298\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.i9_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIU0079_2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21937\,
            in1 => \_gnd_net_\,
            in2 => \N__16512\,
            in3 => \N__19547\,
            lcout => \Lab_UT.dictrl.N_2000_0\,
            ltout => \Lab_UT.dictrl.N_2000_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKPIVI_2_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__16722\,
            in2 => \N__16509\,
            in3 => \N__21941\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIGJHP81_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18453\,
            in1 => \N__18432\,
            in2 => \N__21943\,
            in3 => \N__20130\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__20132\,
            in1 => \N__21912\,
            in2 => \N__18441\,
            in3 => \N__18456\,
            lcout => \Lab_UT.dictrl.state_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22813\,
            ce => \N__18249\,
            sr => \N__22500\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__18454\,
            in1 => \N__18433\,
            in2 => \N__21944\,
            in3 => \N__20133\,
            lcout => \Lab_UT.dictrl.state_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22813\,
            ce => \N__18249\,
            sr => \N__22500\
        );

    \Lab_UT.dictrl.state_0_esr_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__20131\,
            in1 => \N__21910\,
            in2 => \N__18440\,
            in3 => \N__18455\,
            lcout => \Lab_UT.dictrl.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22813\,
            ce => \N__18249\,
            sr => \N__22500\
        );

    \Lab_UT.dictrl.state_ret_1_ess_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001101100001111"
        )
    port map (
            in0 => \N__21913\,
            in1 => \N__19572\,
            in2 => \N__16788\,
            in3 => \N__20134\,
            lcout => \Lab_UT.dictrl.state_i_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22813\,
            ce => \N__18249\,
            sr => \N__22500\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNIHOSE_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16776\,
            in2 => \_gnd_net_\,
            in3 => \N__21254\,
            lcout => \Lab_UT.dicLdAMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_2_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__21911\,
            in1 => \N__16718\,
            in2 => \N__20174\,
            in3 => \N__16704\,
            lcout => \Lab_UT.dictrl.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22813\,
            ce => \N__18249\,
            sr => \N__22500\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__16847\,
            in1 => \_gnd_net_\,
            in2 => \N__20034\,
            in3 => \N__16866\,
            lcout => \Lab_UT.dictrl.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16865\,
            in1 => \N__20030\,
            in2 => \_gnd_net_\,
            in3 => \N__16846\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUQEL8_0_1_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__16689\,
            in1 => \N__16682\,
            in2 => \N__16659\,
            in3 => \N__21295\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.i9_mux_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIU0079_0_2_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19546\,
            in2 => \N__16656\,
            in3 => \N__21929\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_2000_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNII6FQI_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__21930\,
            in1 => \N__16653\,
            in2 => \N__16647\,
            in3 => \N__20118\,
            lcout => \Lab_UT_dictrl_next_state_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU5J2B_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16994\,
            in1 => \N__16899\,
            in2 => \_gnd_net_\,
            in3 => \N__19026\,
            lcout => \Lab_UT.dictrl.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TO6_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21157\,
            in1 => \N__19586\,
            in2 => \_gnd_net_\,
            in3 => \N__22091\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6\,
            ltout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIHF8LB_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__18786\,
            in1 => \N__17006\,
            in2 => \N__16893\,
            in3 => \N__18893\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_96_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNICE00K_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18374\,
            in2 => \N__16890\,
            in3 => \N__21343\,
            lcout => \Lab_UT.dictrl.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIQ1339_3_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__22092\,
            in1 => \N__16887\,
            in2 => \_gnd_net_\,
            in3 => \N__16880\,
            lcout => \Lab_UT.dictrl.N_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIFKL21_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__21724\,
            in1 => \N__17082\,
            in2 => \N__17111\,
            in3 => \N__18282\,
            lcout => \Lab_UT.dictrl.g1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIS94O2_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18981\,
            in1 => \N__16854\,
            in2 => \N__17088\,
            in3 => \N__16827\,
            lcout => \Lab_UT.dictrl.N_119_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__16806\,
            in1 => \N__16797\,
            in2 => \N__19554\,
            in3 => \N__21945\,
            lcout => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNI0DI21_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__17086\,
            in1 => \N__18281\,
            in2 => \N__21579\,
            in3 => \N__17391\,
            lcout => \Lab_UT.dictrl.g0_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_13_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18300\,
            in1 => \N__17104\,
            in2 => \N__17087\,
            in3 => \N__21723\,
            lcout => \Lab_UT.dictrl.g1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIEIOO8_0_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__21949\,
            in1 => \N__16905\,
            in2 => \N__21975\,
            in3 => \N__16917\,
            lcout => \Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIPHQ67_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000001000"
        )
    port map (
            in0 => \N__17043\,
            in1 => \N__16923\,
            in2 => \N__21147\,
            in3 => \N__22056\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1300_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOH1FC_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__16998\,
            in1 => \N__18889\,
            in2 => \N__16956\,
            in3 => \N__16953\,
            lcout => \Lab_UT.dictrl.N_96_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOJ371_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__21125\,
            in1 => \N__20855\,
            in2 => \N__21946\,
            in3 => \N__20652\,
            lcout => \Lab_UT.dictrl.g0_4_a4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_5_x1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21432\,
            in1 => \N__17429\,
            in2 => \N__21648\,
            in3 => \N__21720\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_5_ns_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16947\,
            in3 => \N__16941\,
            lcout => \Lab_UT.dictrl.g0_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIP5KF4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21947\,
            in1 => \N__21145\,
            in2 => \N__19902\,
            in3 => \N__22040\,
            lcout => \Lab_UT.dictrl.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIN8JN3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__19899\,
            in1 => \N__17121\,
            in2 => \N__18888\,
            in3 => \N__16911\,
            lcout => \Lab_UT.dictrl.N_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_3_RNI9ARR_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__21628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21561\,
            lcout => \N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m33_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__17430\,
            in1 => \N__21721\,
            in2 => \N__19077\,
            in3 => \N__19044\,
            lcout => \Lab_UT.dictrl.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m30_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__17194\,
            in1 => \N__17387\,
            in2 => \N__17276\,
            in3 => \N__17346\,
            lcout => \Lab_UT.dictrl.N_98_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_28_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__17313\,
            in1 => \N__17269\,
            in2 => \N__17244\,
            in3 => \N__17196\,
            lcout => \Lab_UT.dictrl.g1_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m31_ns_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17235\,
            in2 => \_gnd_net_\,
            in3 => \N__17202\,
            lcout => \Lab_UT.dictrl.N_84\,
            ltout => \Lab_UT.dictrl.N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__17195\,
            in1 => \N__17163\,
            in2 => \N__17154\,
            in3 => \N__20853\,
            lcout => \Lab_UT.dictrl.g1_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.shifter_ret_1_RNI1OGT_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20702\,
            in1 => \N__17151\,
            in2 => \_gnd_net_\,
            in3 => \N__18191\,
            lcout => \Lab_UT.dictrl.m68_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIG3207_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__19900\,
            in1 => \N__20703\,
            in2 => \N__17130\,
            in3 => \N__22020\,
            lcout => \Lab_UT.dictrl.N_95_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_4_a4_5_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20984\,
            in1 => \N__21077\,
            in2 => \N__21580\,
            in3 => \N__21621\,
            lcout => \Lab_UT.dictrl.g0_4_a4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__17461\,
            in1 => \N__17858\,
            in2 => \N__17958\,
            in3 => \N__17643\,
            lcout => \Lab_UT.didp.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17460\,
            in2 => \_gnd_net_\,
            in3 => \N__17925\,
            lcout => \Lab_UT.didp.countrce2.un13_qPone\,
            ltout => \Lab_UT.didp.countrce2.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_3_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17697\,
            in3 => \N__17510\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__17895\,
            in1 => \N__18738\,
            in2 => \N__17694\,
            in3 => \N__17676\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__17957\,
            in1 => \N__17677\,
            in2 => \N__17691\,
            in3 => \N__17859\,
            lcout => \Lab_UT.didp.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22855\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__17886\,
            in1 => \N__18231\,
            in2 => \_gnd_net_\,
            in3 => \N__17462\,
            lcout => \Lab_UT.didp.countrce2.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000111100"
        )
    port map (
            in0 => \N__17637\,
            in1 => \N__17526\,
            in2 => \N__17517\,
            in3 => \N__17890\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__17948\,
            in2 => \N__17520\,
            in3 => \N__17852\,
            lcout => \Lab_UT.didp.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_1_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__20892\,
            in1 => \N__17463\,
            in2 => \N__17894\,
            in3 => \N__17926\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__17927\,
            in1 => \N__17947\,
            in2 => \N__17931\,
            in3 => \N__17851\,
            lcout => \Lab_UT.didp.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__19702\,
            in1 => \N__19981\,
            in2 => \N__17748\,
            in3 => \N__19944\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22849\,
            ce => \N__18252\,
            sr => \N__22507\
        );

    \Lab_UT.dictrl.state_ret_8_ess_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__19946\,
            in1 => \N__17746\,
            in2 => \N__19989\,
            in3 => \N__19704\,
            lcout => \Lab_UT.LdStens_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22849\,
            ce => \N__18252\,
            sr => \N__22507\
        );

    \Lab_UT.dictrl.state_ret_7_esr_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19945\,
            in1 => \N__17745\,
            in2 => \N__19988\,
            in3 => \N__19703\,
            lcout => \Lab_UT.LdStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22849\,
            ce => \N__18252\,
            sr => \N__22507\
        );

    \Lab_UT.didp.ce_RNI62AM_1_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17865\,
            lcout => \Lab_UT.didp.un1_dicLdStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__18227\,
            in1 => \N__17815\,
            in2 => \_gnd_net_\,
            in3 => \N__17799\,
            lcout => \Lab_UT.didp.countrce1.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_ess_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__19701\,
            in1 => \N__19973\,
            in2 => \N__17747\,
            in3 => \N__19943\,
            lcout => \Lab_UT.LdSones_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22841\,
            ce => \N__18251\,
            sr => \N__22506\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19377\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19147\,
            in2 => \_gnd_net_\,
            in3 => \N__18042\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19186\,
            in2 => \_gnd_net_\,
            in3 => \N__18033\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19799\,
            in2 => \_gnd_net_\,
            in3 => \N__18030\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__19402\,
            in1 => \N__22981\,
            in2 => \N__19122\,
            in3 => \N__18027\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22834\,
            ce => \N__19350\,
            sr => \N__22530\
        );

    \Lab_UT.dictrl.state_ret_5_ess_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__17989\,
            in1 => \N__18401\,
            in2 => \_gnd_net_\,
            in3 => \N__20509\,
            lcout => \Lab_UT.dictrl.state_i_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__18250\,
            sr => \N__22503\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17988\,
            in1 => \N__18363\,
            in2 => \_gnd_net_\,
            in3 => \N__20414\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010011100001111"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__18378\,
            in2 => \N__18003\,
            in3 => \N__21299\,
            lcout => \Lab_UT.dictrl.state_i_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__18250\,
            sr => \N__22503\
        );

    \Lab_UT.dictrl.state_ret_6_esr_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011010100000000"
        )
    port map (
            in0 => \N__18402\,
            in1 => \N__20510\,
            in2 => \N__17994\,
            in3 => \N__19700\,
            lcout => \Lab_UT.dictrl.dicLdStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__18250\,
            sr => \N__22503\
        );

    \Lab_UT.dictrl.state_0_esr_RNI9CU3Q_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101100"
        )
    port map (
            in0 => \N__20413\,
            in1 => \N__18317\,
            in2 => \N__20177\,
            in3 => \N__21880\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI4L025_3_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__22198\,
            in1 => \N__18609\,
            in2 => \N__20332\,
            in3 => \N__21294\,
            lcout => \Lab_UT.dictrl.N_101\,
            ltout => \Lab_UT.dictrl.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI3QHJ5_1_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18333\,
            in2 => \N__18321\,
            in3 => \N__21879\,
            lcout => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1\,
            ltout => \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_1_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__21885\,
            in1 => \N__18318\,
            in2 => \N__18303\,
            in3 => \N__20151\,
            lcout => \Lab_UT.dictrl.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22820\,
            ce => \N__18248\,
            sr => \N__22502\
        );

    \Lab_UT.dictrl.state_0_esr_3_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__19259\,
            in1 => \N__19291\,
            in2 => \N__20179\,
            in3 => \N__21886\,
            lcout => \Lab_UT.dictrl.stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22820\,
            ce => \N__18248\,
            sr => \N__22502\
        );

    \Lab_UT.dictrl.state_0_fast_esr_3_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__20159\,
            in1 => \N__19293\,
            in2 => \N__21936\,
            in3 => \N__19260\,
            lcout => \Lab_UT.dictrl.state_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22820\,
            ce => \N__18248\,
            sr => \N__22502\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__19257\,
            in1 => \N__19290\,
            in2 => \N__20178\,
            in3 => \N__21881\,
            lcout => \Lab_UT.dictrl.state_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22820\,
            ce => \N__18248\,
            sr => \N__22502\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__20158\,
            in1 => \N__19292\,
            in2 => \N__21935\,
            in3 => \N__19258\,
            lcout => \Lab_UT.dictrl.state_3_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22820\,
            ce => \N__18248\,
            sr => \N__22502\
        );

    \Lab_UT.dictrl.g0_30_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18549\,
            in1 => \N__18216\,
            in2 => \N__18093\,
            in3 => \N__18081\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_116_mux_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIU2C38_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011110011"
        )
    port map (
            in0 => \N__20337\,
            in1 => \N__22202\,
            in2 => \N__18051\,
            in3 => \N__22104\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_120_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNI5OGCH_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000001"
        )
    port map (
            in0 => \N__21296\,
            in1 => \N__21931\,
            in2 => \N__18459\,
            in3 => \N__18420\,
            lcout => \Lab_UT.dictrl.N_1302_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIHNKSM_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001010101"
        )
    port map (
            in0 => \N__18807\,
            in1 => \N__18585\,
            in2 => \N__20367\,
            in3 => \N__21297\,
            lcout => \Lab_UT.dictrl.N_119_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNIVIE9H_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000101"
        )
    port map (
            in0 => \N__18387\,
            in1 => \N__18419\,
            in2 => \N__21950\,
            in3 => \N__21344\,
            lcout => \Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIOT908_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101111"
        )
    port map (
            in0 => \N__20486\,
            in1 => \N__20336\,
            in2 => \N__22249\,
            in3 => \N__22105\,
            lcout => \Lab_UT.dictrl.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI4CET7_3_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100011111"
        )
    port map (
            in0 => \N__22220\,
            in1 => \N__20485\,
            in2 => \N__20366\,
            in3 => \N__19024\,
            lcout => \Lab_UT.dictrl.N_99\,
            ltout => \Lab_UT.dictrl.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__21345\,
            in1 => \N__18359\,
            in2 => \N__18348\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18345\,
            in2 => \N__18336\,
            in3 => \N__20168\,
            lcout => \Lab_UT.dictrl.next_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22805\,
            ce => \N__22295\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIH7T88_3_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100100010"
        )
    port map (
            in0 => \N__22090\,
            in1 => \N__20305\,
            in2 => \N__19025\,
            in3 => \N__22219\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI51E3N_1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__21342\,
            in1 => \_gnd_net_\,
            in2 => \N__18324\,
            in3 => \N__18750\,
            lcout => \Lab_UT.dictrl.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI48008_3_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__22089\,
            in1 => \N__20304\,
            in2 => \N__18899\,
            in3 => \N__18777\,
            lcout => \Lab_UT.dictrl.N_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI89VA1_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20300\,
            in1 => \N__22216\,
            in2 => \N__21948\,
            in3 => \N__21340\,
            lcout => \Lab_UT.dictrl.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI4CET7_0_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100011111"
        )
    port map (
            in0 => \N__22217\,
            in1 => \N__20481\,
            in2 => \N__20346\,
            in3 => \N__19016\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_99_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIJGPPK_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21341\,
            in2 => \N__18594\,
            in3 => \N__18591\,
            lcout => \Lab_UT.dictrl.N_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIOIJR7_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__22218\,
            in1 => \N__19017\,
            in2 => \_gnd_net_\,
            in3 => \N__22088\,
            lcout => \Lab_UT.dictrl.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIPED74_3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20341\,
            in1 => \N__18897\,
            in2 => \_gnd_net_\,
            in3 => \N__18776\,
            lcout => \Lab_UT.dictrl.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__20970\,
            in1 => \N__21065\,
            in2 => \N__18900\,
            in3 => \N__21650\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_37_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__20969\,
            in1 => \N__21064\,
            in2 => \N__21572\,
            in3 => \N__21649\,
            lcout => \Lab_UT.dictrl.N_98_mux_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_5_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21651\,
            in1 => \N__18548\,
            in2 => \N__20664\,
            in3 => \N__21556\,
            lcout => OPEN,
            ltout => \resetGen.escKeyZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18498\,
            in1 => \N__19800\,
            in2 => \N__18486\,
            in3 => \N__19740\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKE4Q8_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011111010"
        )
    port map (
            in0 => \N__22039\,
            in1 => \N__18887\,
            in2 => \N__22263\,
            in3 => \N__18921\,
            lcout => \Lab_UT.dictrl.g2_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIGU6P7_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__19894\,
            in1 => \N__18912\,
            in2 => \N__18898\,
            in3 => \N__22038\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_95_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI9TD6E_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__22247\,
            in1 => \_gnd_net_\,
            in2 => \N__18810\,
            in3 => \N__18959\,
            lcout => \Lab_UT.dictrl.N_103_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__20865\,
            in1 => \N__19080\,
            in2 => \N__18798\,
            in3 => \N__20660\,
            lcout => \Lab_UT.dictrl.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m47_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19079\,
            in1 => \N__20864\,
            in2 => \_gnd_net_\,
            in3 => \N__19047\,
            lcout => \Lab_UT.dictrl.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIT67DE_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__18960\,
            in1 => \_gnd_net_\,
            in2 => \N__18762\,
            in3 => \N__22248\,
            lcout => \Lab_UT.dictrl.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m63_0_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011111001111"
        )
    port map (
            in0 => \N__19046\,
            in1 => \N__18714\,
            in2 => \N__19078\,
            in3 => \N__21728\,
            lcout => \Lab_UT.dictrl.m63_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIVHJND_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22243\,
            in1 => \N__18933\,
            in2 => \_gnd_net_\,
            in3 => \N__18600\,
            lcout => \Lab_UT.dictrl.N_103_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m48_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000001000000"
        )
    port map (
            in0 => \N__20854\,
            in1 => \N__19068\,
            in2 => \N__20706\,
            in3 => \N__19045\,
            lcout => \Lab_UT.dictrl.N_89\,
            ltout => \Lab_UT.dictrl.N_89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNI3DTV5_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__18990\,
            in2 => \N__18984\,
            in3 => \N__18980\,
            lcout => \Lab_UT.dictrl.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIPS7A6_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101011111010"
        )
    port map (
            in0 => \N__18951\,
            in1 => \N__20704\,
            in2 => \N__19893\,
            in3 => \N__18939\,
            lcout => \Lab_UT.dictrl.N_102_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23063\,
            in1 => \N__20545\,
            in2 => \N__22929\,
            in3 => \N__20581\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23047\,
            in2 => \N__18927\,
            in3 => \N__20562\,
            lcout => \buart__rx_ser_clk\,
            ltout => \buart__rx_ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__23073\,
            in1 => \N__22983\,
            in2 => \N__18924\,
            in3 => \N__20546\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__20582\,
            in1 => \_gnd_net_\,
            in2 => \N__22994\,
            in3 => \N__20564\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__23048\,
            in1 => \N__23021\,
            in2 => \N__23034\,
            in3 => \N__22987\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__22982\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20563\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNICF9U4_3_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__22869\,
            in1 => \N__21897\,
            in2 => \_gnd_net_\,
            in3 => \N__19236\,
            lcout => \Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m91_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__19371\,
            in1 => \N__19126\,
            in2 => \N__19167\,
            in3 => \N__19198\,
            lcout => \Lab_UT.dictrl.N_102_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m81_e_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__19127\,
            in1 => \N__19165\,
            in2 => \_gnd_net_\,
            in3 => \N__19774\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m82_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001000"
        )
    port map (
            in0 => \N__19372\,
            in1 => \N__23016\,
            in2 => \N__19221\,
            in3 => \N__19199\,
            lcout => \buart__rx_sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__19197\,
            in1 => \N__19161\,
            in2 => \N__19128\,
            in3 => \N__19370\,
            lcout => \buart__rx_valid_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__19098\,
            in1 => \N__23022\,
            in2 => \_gnd_net_\,
            in3 => \N__19509\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m89_bm_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__19417\,
            in1 => \N__19452\,
            in2 => \N__19503\,
            in3 => \N__19776\,
            lcout => m89_bm,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.N_27_0_i_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__19726\,
            in1 => \_gnd_net_\,
            in2 => \N__19789\,
            in3 => \N__19418\,
            lcout => \buart__rx_N_27_0_i\,
            ltout => \buart__rx_N_27_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011010100111010"
        )
    port map (
            in0 => \N__19092\,
            in1 => \N__22980\,
            in2 => \N__19083\,
            in3 => \N__19781\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22842\,
            ce => \N__19345\,
            sr => \N__22532\
        );

    \Lab_UT.dictrl.m9_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19451\,
            in1 => \N__19498\,
            in2 => \_gnd_net_\,
            in3 => \N__19416\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_107_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m89_am_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19775\,
            in2 => \N__19512\,
            in3 => \N__19725\,
            lcout => m89_am,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m10_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19777\,
            in1 => \N__19502\,
            in2 => \N__19468\,
            in3 => \N__19419\,
            lcout => \buart__rx_startbit\,
            ltout => \buart__rx_startbit_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001110100101110"
        )
    port map (
            in0 => \N__22899\,
            in1 => \N__19401\,
            in2 => \N__19380\,
            in3 => \N__19376\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22842\,
            ce => \N__19345\,
            sr => \N__22532\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_6_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__21837\,
            in2 => \_gnd_net_\,
            in3 => \N__19320\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_2000_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__21838\,
            in1 => \N__19308\,
            in2 => \N__19296\,
            in3 => \N__20182\,
            lcout => \Lab_UT.dictrl.next_state_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_3_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__22580\,
            in1 => \N__21835\,
            in2 => \_gnd_net_\,
            in3 => \N__19638\,
            lcout => \Lab_UT.dictrl.state_ret_12_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22582\,
            in1 => \N__19677\,
            in2 => \_gnd_net_\,
            in3 => \N__19640\,
            lcout => \Lab_UT.dictrl.state_ret_12and_a0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIKRG8A_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__19279\,
            in1 => \N__19256\,
            in2 => \N__21903\,
            in3 => \N__20141\,
            lcout => \Lab_UT_dictrl_next_state_3\,
            ltout => \Lab_UT_dictrl_next_state_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__22581\,
            in1 => \N__21836\,
            in2 => \N__20016\,
            in3 => \N__19639\,
            lcout => \Lab_UT.dictrl.state_ret_12_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20013\,
            in1 => \N__20007\,
            in2 => \_gnd_net_\,
            in3 => \N__20001\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_12and_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__19995\,
            in1 => \N__19972\,
            in2 => \N__19950\,
            in3 => \N__19942\,
            lcout => \Lab_UT_dictrl_un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22826\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNIH05S_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__21367\,
            in1 => \N__19887\,
            in2 => \_gnd_net_\,
            in3 => \N__21820\,
            lcout => \Lab_UT.dictrl.m46_i_0_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19788\,
            in2 => \_gnd_net_\,
            in3 => \N__19736\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_RNIMHUCC_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__21839\,
            in1 => \N__19676\,
            in2 => \N__19650\,
            in3 => \N__19646\,
            lcout => \resetGen.r_m3_i_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_2_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010110000000"
        )
    port map (
            in0 => \N__21369\,
            in1 => \N__20532\,
            in2 => \N__22264\,
            in3 => \N__19593\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.i9_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20183\,
            in2 => \N__19575\,
            in3 => \N__19571\,
            lcout => \Lab_UT.dictrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22815\,
            ce => \N__22282\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__22252\,
            in1 => \N__20531\,
            in2 => \N__20373\,
            in3 => \N__22107\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21370\,
            in2 => \N__20517\,
            in3 => \N__20439\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__20184\,
            in1 => \N__20514\,
            in2 => \N__20490\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.next_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22815\,
            ce => \N__22282\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_1_0_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011001110"
        )
    port map (
            in0 => \N__22106\,
            in1 => \N__22251\,
            in2 => \N__20372\,
            in3 => \N__20487\,
            lcout => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIL2ATH_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__21735\,
            in1 => \N__21981\,
            in2 => \N__20433\,
            in3 => \N__22097\,
            lcout => \Lab_UT.dictrl.N_1302_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIGENTQ_2_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__20418\,
            in1 => \N__20180\,
            in2 => \N__21942\,
            in3 => \N__20394\,
            lcout => \N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI38BCN_3_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000111011"
        )
    port map (
            in0 => \N__20385\,
            in1 => \N__21368\,
            in2 => \N__20369\,
            in3 => \N__20205\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_119_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIIE1Q91_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__21899\,
            in1 => \N__20193\,
            in2 => \N__20187\,
            in3 => \N__20181\,
            lcout => \Lab_UT_dictrl_next_state_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_4_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21652\,
            in1 => \N__20980\,
            in2 => \N__21581\,
            in3 => \N__21441\,
            lcout => \Lab_UT.dictrl.g1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI6KC68_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__22250\,
            in1 => \N__20991\,
            in2 => \N__22119\,
            in3 => \N__22103\,
            lcout => \Lab_UT.dictrl.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNISBBJ4_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21968\,
            in1 => \N__21898\,
            in2 => \_gnd_net_\,
            in3 => \N__21183\,
            lcout => \Lab_UT.dictrl.m46_i_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_5_RNIIJHP1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__21729\,
            in1 => \N__21657\,
            in2 => \N__21582\,
            in3 => \N__21440\,
            lcout => OPEN,
            ltout => \g0_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU7Q14_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100000"
        )
    port map (
            in0 => \N__21167\,
            in1 => \N__21384\,
            in2 => \N__21198\,
            in3 => \N__21195\,
            lcout => \Lab_UT.dictrl.g1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIK8B43_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20589\,
            in1 => \N__21177\,
            in2 => \N__21168\,
            in3 => \N__21081\,
            lcout => \Lab_UT.dictrl.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_ret_6_rep1_RNI4S9J1_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__20985\,
            in1 => \N__20852\,
            in2 => \N__20705\,
            in3 => \N__20651\,
            lcout => m46_i_0_a3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20583\,
            in2 => \N__20568\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_3_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20547\,
            in2 => \_gnd_net_\,
            in3 => \N__23067\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22990\,
            in1 => \N__23064\,
            in2 => \_gnd_net_\,
            in3 => \N__23052\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__22856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23049\,
            in2 => \_gnd_net_\,
            in3 => \N__23025\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__22928\,
            in1 => \N__23020\,
            in2 => \N__22995\,
            in3 => \N__22932\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22856\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22900\,
            lcout => \Lab_UT.dictrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22850\,
            ce => \N__22299\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_ctle_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22583\,
            in2 => \_gnd_net_\,
            in3 => \N__22558\,
            lcout => bu_rx_data_rdy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_RNIAL6V33_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__22332\,
            in1 => \N__22326\,
            in2 => \N__22320\,
            in3 => \N__22305\,
            lcout => \rst_RNIAL6V33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
