-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 19 2019 22:38:35

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23320\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23267\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23222\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23210\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23198\ : std_logic;
signal \N__23197\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23195\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23170\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23150\ : std_logic;
signal \N__23147\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23141\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23072\ : std_logic;
signal \N__23069\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23047\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23045\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23033\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22970\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22959\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22953\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22925\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22831\ : std_logic;
signal \N__22828\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22769\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22760\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22749\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22736\ : std_logic;
signal \N__22733\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22727\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22336\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22318\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22301\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22288\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22285\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22274\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22271\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22068\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22039\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22014\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22011\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22005\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22002\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21996\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21974\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21954\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21945\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21942\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21939\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21792\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21717\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21708\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21699\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21648\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21642\ : std_logic;
signal \N__21623\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21466\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21435\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21369\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21274\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21244\ : std_logic;
signal \N__21241\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21174\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21130\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21123\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21067\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21064\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21061\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20954\ : std_logic;
signal \N__20953\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20951\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20899\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20858\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20848\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20741\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20726\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20708\ : std_logic;
signal \N__20705\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20681\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20657\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20654\ : std_logic;
signal \N__20651\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20646\ : std_logic;
signal \N__20645\ : std_logic;
signal \N__20642\ : std_logic;
signal \N__20639\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20609\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20516\ : std_logic;
signal \N__20513\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20486\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20478\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20460\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20441\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20420\ : std_logic;
signal \N__20417\ : std_logic;
signal \N__20414\ : std_logic;
signal \N__20411\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20405\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20378\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20363\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20339\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20272\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20204\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20184\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20111\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20108\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20080\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20030\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20024\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20021\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19908\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19879\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19846\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19797\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19781\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19673\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19634\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19628\ : std_logic;
signal \N__19625\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19601\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19565\ : std_logic;
signal \N__19556\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19503\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19475\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19419\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19413\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19406\ : std_logic;
signal \N__19403\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19052\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18899\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18722\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18671\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18647\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18629\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18623\ : std_logic;
signal \N__18620\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18608\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18554\ : std_logic;
signal \N__18551\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18524\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18398\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18383\ : std_logic;
signal \N__18380\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18289\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18209\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18176\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18116\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18113\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18005\ : std_logic;
signal \N__18002\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17957\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17836\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17699\ : std_logic;
signal \N__17696\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17648\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17636\ : std_logic;
signal \N__17633\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17600\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17516\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17429\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17403\ : std_logic;
signal \N__17400\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17321\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17255\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17237\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17174\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17171\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17000\ : std_logic;
signal \N__16997\ : std_logic;
signal \N__16994\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16814\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16766\ : std_logic;
signal \N__16763\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16754\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16745\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16547\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16403\ : std_logic;
signal \N__16400\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16390\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16349\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16334\ : std_logic;
signal \N__16331\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16301\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16274\ : std_logic;
signal \N__16271\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16259\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16208\ : std_logic;
signal \N__16205\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16151\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16127\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16106\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16076\ : std_logic;
signal \N__16073\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16055\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16046\ : std_logic;
signal \N__16043\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16040\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15854\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15797\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15741\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15722\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15383\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15217\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15214\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14891\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14810\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14506\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14272\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14090\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14048\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13994\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13988\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13889\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13793\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13691\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13519\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12904\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu0.un88_ci_3_cascade_\ : std_logic;
signal \uu0.un55_ci_cascade_\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \INVuu2.r_data_reg_2C_net\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_14\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.un4_l_count_18_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un4_l_count_11\ : std_logic;
signal \uu0.un4_l_count_16\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det_cascade_\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.un404_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.mem0.w_data_0\ : std_logic;
signal \uu2.mem0.N_30_i_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \Lab_UT.dispString.m32_ns_1_cascade_\ : std_logic;
signal \Lab_UT.sec1Z0Z_3\ : std_logic;
signal \Lab_UT.sec2Z0Z_1\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_5\ : std_logic;
signal \Lab_UT.dispString.m35_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOut_RNO_0Z0Z_1\ : std_logic;
signal \Lab_UT.sec2Z0Z_0\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.N_46\ : std_logic;
signal \Lab_UT.min2Z0Z_1\ : std_logic;
signal \Lab_UT.min2Z0Z_2\ : std_logic;
signal \Lab_UT.sec1Z0Z_2\ : std_logic;
signal \Lab_UT.dicLdAStens_0_cascade_\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \resetGen.reset_count_2_0_4\ : std_logic;
signal \Lab_UT.three_2_1_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_fastZ0Z_2\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_6_cascade_\ : std_logic;
signal \Lab_UT.min2Z0Z_3\ : std_logic;
signal \Lab_UT.min1Z0Z_1\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.didp.regrce1.LdASones_0\ : std_logic;
signal \buart.Z_rx.valid_0_cascade_\ : std_logic;
signal \buart.Z_rx.idle_0_cascade_\ : std_logic;
signal \buart.Z_rx.idle_cascade_\ : std_logic;
signal \buart.Z_rx.N_27_0_i_cascade_\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal clk : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_0_1_3\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_33_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_\ : std_logic;
signal \uu2.mem0.N_409\ : std_logic;
signal \uu2.N_34_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_4C_net\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_1\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \Lab_UT.dispString.m40_ns_1\ : std_logic;
signal \Lab_UT.min1Z0Z_3\ : std_logic;
signal \Lab_UT.dispString.N_77_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_80\ : std_logic;
signal \Lab_UT.sec2Z0Z_3\ : std_logic;
signal \Lab_UT.dispString.N_86_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_89\ : std_logic;
signal \Lab_UT.min2Z0Z_0\ : std_logic;
signal \Lab_UT.dispString.m49_ns_1\ : std_logic;
signal \Lab_UT.sec1Z0Z_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \Lab_UT.min1Z0Z_0\ : std_logic;
signal \Lab_UT.dispString.m25_ns_1\ : std_logic;
signal \Lab_UT.min1Z0Z_2\ : std_logic;
signal \Lab_UT.dispString.N_65\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_6\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_2\ : std_logic;
signal \Lab_UT.sec2Z0Z_2\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.N_68\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_5\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_11\ : std_logic;
signal \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\ : std_logic;
signal \Lab_UT.didp.q_fast_0\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_fastZ0Z_3\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_3\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_2\ : std_logic;
signal \Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_12\ : std_logic;
signal \Lab_UT.three_2_0_cascade_\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_fastZ0Z_1\ : std_logic;
signal \Lab_UT.didp.countrce3.q_fastZ0Z_1\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_fastZ0Z_3\ : std_logic;
signal \Lab_UT.didp.q_fast_3\ : std_logic;
signal \Lab_UT.didp.countrce3.did_alarmMatch_0\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.dicLdAMones_0_cascade_\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.dicLdAMones_0\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \resetGen.escKeyZ0Z_5\ : std_logic;
signal \resetGen.escKeyZ0Z_4_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.ser_clk_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.startbit_cascade_\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \bfn_6_2_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \uu2.un3_w_addr_user_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_44\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_33_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_43\ : std_logic;
signal \uu2.N_34\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_42\ : std_logic;
signal \uu2.N_49\ : std_logic;
signal \uu2.N_57_cascade_\ : std_logic;
signal \uu2.w_data_i_a3_0_5\ : std_logic;
signal \uu2.mem0.w_data_0_a3_0_6_cascade_\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.w_data_displaying_2_i_a2_i_a2_0_0\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_4\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \uu2.un1_w_user_crZ0Z_4\ : std_logic;
signal \uu2_un1_w_user_cr_0_cascade_\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.dictrl.G_64\ : std_logic;
signal \Lab_UT.alarmMatch\ : std_logic;
signal \Lab_UT.dictrl.idle_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\ : std_logic;
signal \Lab_UT.alarmchar9\ : std_logic;
signal \Lab_UT.alarmchar10\ : std_logic;
signal \Lab_UT.alarmchar10_i_2\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_1\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_i_3_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z_1\ : std_logic;
signal \Lab_UT.alarmchar_2_1_1\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_1\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3\ : std_logic;
signal \Lab_UT.didp.q_fast_1\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.three_2_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.reset_12_3_3_cascade_\ : std_logic;
signal \Lab_UT.didp.reset_12_1_3_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0\ : std_logic;
signal \uu0_sec_clkD\ : std_logic;
signal \Lab_UT.didp.regrce4.LdAMtens_0\ : std_logic;
signal \Lab_UT.didp.ce_11_0_2\ : std_logic;
signal \Lab_UT.didp.un26_ce_0_cascade_\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.ce_12_0_3_cascade_\ : std_logic;
signal \Lab_UT.didp.un26_ce_0\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.nine_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.nine\ : std_logic;
signal \Lab_UT.five\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.ser_clk\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.g2_0_1_0_cascade_\ : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g2_1_0_0\ : std_logic;
signal \INVuu2.w_addr_user_5C_net\ : std_logic;
signal \uu2.un1_w_user_lf_0_0\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4\ : std_logic;
signal \uu2.un20_w_addr_userZ0Z_1\ : std_logic;
signal \uu2.un3_w_addr_user\ : std_logic;
signal \uu2.un20_w_addr_userZ0Z_1_cascade_\ : std_logic;
signal \uu2.w_addr_user_RNI43E87Z0Z_2_cascade_\ : std_logic;
signal \uu2.un28_w_addr_user_i\ : std_logic;
signal \INVuu2.w_addr_user_0C_net\ : std_logic;
signal \uu2.un3_w_addr_user_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.un426_ci_3_cascade_\ : std_logic;
signal \uu2.un426_ci_3\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.w_addr_user_RNI43E87Z0Z_2\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_42\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_8C_net\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.vbuf_w_addr_user.un448_ci_0\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_0\ : std_logic;
signal \INVuu2.bitmap_40C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.N_97_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_0_0\ : std_logic;
signal \Lab_UT.dictrl.un1_next_alarmstate21_0\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.sec1Z0Z_1\ : std_logic;
signal rst : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_6\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_0Z0Z_0\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.three_2\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_\ : std_logic;
signal \Lab_UT.dicLdSones_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_2\ : std_logic;
signal \Lab_UT.dictrl.g3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_2\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.dictrl.g0_1_2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_29_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_30_0\ : std_logic;
signal \Lab_UT.dictrl.N_30_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.i6_mux_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.dicLdAMones_0_sx_cascade_\ : std_logic;
signal \Lab_UT.dicLdAMones_1\ : std_logic;
signal \Lab_UT.dictrl.g0_1_3\ : std_logic;
signal \Lab_UT.dictrl.g2_1_0_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_7_1_0\ : std_logic;
signal bu_rx_data_fast_4 : std_logic;
signal \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state18_1_0\ : std_logic;
signal \Lab_UT.dictrl.g1_0_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1\ : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal \uu2.mem0.N_98_0_cascade_\ : std_logic;
signal \uu2.mem0.G_11_0_0_a3_0_2\ : std_logic;
signal \uu2.mem0.N_62_cascade_\ : std_logic;
signal \uu2.mem0.N_36\ : std_logic;
signal \uu2.mem0.N_9_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_26_bm_1\ : std_logic;
signal \uu2.bitmap_RNI31F32Z0Z_34_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNIBICU6_0Z0Z_2\ : std_logic;
signal \uu2.N_401_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_RNIBICU6Z0Z_2\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.N_99_cascade_\ : std_logic;
signal \uu2.bitmap_RNI2Q8F1Z0Z_111\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_nesr_3C_net\ : std_logic;
signal \uu2.N_31_0\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.N_98_cascade_\ : std_logic;
signal \uu2.bitmap_RNI04AD1Z0Z_314\ : std_logic;
signal \INVuu2.bitmap_90C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.N_383\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal uu2_un1_w_user_cr_0 : std_logic;
signal \uu2.N_57\ : std_logic;
signal \uu2.N_38\ : std_logic;
signal \uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_7C_net\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_0Z0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_4\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_6\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_0Z0Z_1\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_5\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \INVuu2.bitmap_203C_net\ : std_logic;
signal \Lab_UT.LdASones\ : std_logic;
signal \Lab_UT.LdASones_cascade_\ : std_logic;
signal \Lab_UT.LdSones_i_3\ : std_logic;
signal \Lab_UT.dicRun_2\ : std_logic;
signal \Lab_UT.didp.ce_9_0_0\ : std_logic;
signal \Lab_UT.dicRun_2_cascade_\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_11_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_3_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_3_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_4\ : std_logic;
signal \Lab_UT.dictrl.N_9_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z4\ : std_logic;
signal \Lab_UT.dictrl.N_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_10_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_o4_0\ : std_logic;
signal \Lab_UT.dictrl.N_3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_2_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_o4_0\ : std_logic;
signal \Lab_UT.dictrl.g0_1Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state18_0\ : std_logic;
signal \Lab_UT.dictrl.next_state18_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_7_0\ : std_logic;
signal \Lab_UT.dictrl.N_11\ : std_logic;
signal \Lab_UT.dictrl.g2_2_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g2_1_2\ : std_logic;
signal \Lab_UT.dictrl.g1_5_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_3\ : std_logic;
signal \Lab_UT.dictrl.g0Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_3_cascade_\ : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal \Lab_UT.dictrl.next_state12_0\ : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal \Lab_UT.dictrl.g0_8Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1_3\ : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_28\ : std_logic;
signal \uu2.mem0.N_44\ : std_logic;
signal \uu2.mem0.N_41_cascade_\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_36\ : std_logic;
signal \uu2.mem0.N_24_i_cascade_\ : std_logic;
signal \uu2.N_406\ : std_logic;
signal \uu2.mem0.N_45\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.mem0.G_11_0_0_a2_3_4\ : std_logic;
signal \N_272_mux\ : std_logic;
signal \uu2.mem0.G_11_0_0_a2_3_5_cascade_\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \uu2.mem0.G_11_0_0_0\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_1\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_5\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_4\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_2\ : std_logic;
signal \INVuu2.bitmap_87C_net\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmap_pmux_17_ns_1_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.N_104_cascade_\ : std_logic;
signal \uu2.mem0.G_11_0_0_a3_5_0_cascade_\ : std_logic;
signal \uu2.mem0.N_40\ : std_logic;
signal \uu2.mem0.N_30\ : std_logic;
signal \uu2.w_addr_displaying_2_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_41\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_RNIVAPV6Z0Z_5\ : std_logic;
signal \INVuu2.w_addr_displaying_2_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.bitmap_pmux_20_ns_1_cascade_\ : std_logic;
signal \uu2.mem0.N_108\ : std_logic;
signal \INVuu2.bitmap_194C_net\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.bitmap_pmux_20_ns_1\ : std_logic;
signal \uu2.mem0.N_108_0_cascade_\ : std_logic;
signal \uu2.mem0.N_404_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_16_ns_1_cascade_\ : std_logic;
signal \uu2.N_30_i\ : std_logic;
signal \uu2.mem0.N_22_cascade_\ : std_logic;
signal \uu2.mem0.G_11_0_0_a3_6_0\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.N_30_i_1\ : std_logic;
signal \uu2.mem0.N_22_0_cascade_\ : std_logic;
signal \uu2.N_104\ : std_logic;
signal \uu2.mem0.bitmap_pmux_27_ns_1_0\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.mem0.N_109\ : std_logic;
signal \uu2.bitmap_pmux_19_ns_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.mem0.N_109_0\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_3\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_5\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_6\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_0\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_1\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \INVuu2.bitmap_218C_net\ : std_logic;
signal \Lab_UT.dictrl.N_14_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_0_3\ : std_logic;
signal \Lab_UT.dictrl.N_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_13_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_6_cascade_\ : std_logic;
signal \Lab_UT.LdStens\ : std_logic;
signal \Lab_UT.state_i_3_2\ : std_logic;
signal \Lab_UT.LdStens_i_3\ : std_logic;
signal \Lab_UT.didp.ce_10_0_1\ : std_logic;
signal \Lab_UT.dictrl.m27_1\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_19_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_19\ : std_logic;
signal \Lab_UT.dictrl.N_11_0_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_5_RNOZ0Z_1\ : std_logic;
signal \Lab_UT.dicRun_1\ : std_logic;
signal \Lab_UT.dictrl.N_10\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_2\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_0_3\ : std_logic;
signal \Lab_UT.dictrl.i6_mux\ : std_logic;
signal \Lab_UT.dictrl.N_15_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_i_3Z0Z_0\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.dictrl.g0_6_o3_2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_5_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_3_0\ : std_logic;
signal \Lab_UT.dictrl.g2_2\ : std_logic;
signal \Lab_UT.dictrl.N_16_0_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a3_0_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a3_0_6_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a3_0_5\ : std_logic;
signal \Lab_UT.dictrl.N_3\ : std_logic;
signal \Lab_UT.dictrl.g1_4\ : std_logic;
signal \Lab_UT.dictrl.gZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.next_state12_1\ : std_logic;
signal \Lab_UT.dictrl.next_state32Z0Z_4\ : std_logic;
signal \Lab_UT.dictrl.g1Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_13_0_0\ : std_logic;
signal \Lab_UT.dictrl.g1_2_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1_1\ : std_logic;
signal \Lab_UT.dictrl.g2_0\ : std_logic;
signal \Lab_UT.dictrl.g1_2_3\ : std_logic;
signal \Lab_UT.dictrl.g0_1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a3_4\ : std_logic;
signal bu_rx_data_4_rep1 : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \Lab_UT.dictrl.g1_4_0\ : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_2 : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \INVuu2.bitmap_34C_net\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_0Z0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment4.segmentUQ_0_4\ : std_logic;
signal \Lab_UT.bcd2segment4.segmentUQ_0_5\ : std_logic;
signal \Lab_UT.bcd2segment4.segmentUQ_0_6\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_0Z0Z_0\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_0Z0Z_1\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_\ : std_logic;
signal \Lab_UT.Run\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \Lab_UT.dictrl.N_39_mux\ : std_logic;
signal \Lab_UT.dictrl.g0_0_a3_2\ : std_logic;
signal \Lab_UT.dictrl.g0_0_0_a3_1\ : std_logic;
signal \Lab_UT.dictrl.un1_next_state66_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_i_a3_1\ : std_logic;
signal \Lab_UT.dicLdAStens_0\ : std_logic;
signal \Lab_UT.dictrl.N_40_mux\ : std_logic;
signal \Lab_UT.state_3\ : std_logic;
signal \Lab_UT.dictrl.N_13_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_16\ : std_logic;
signal \Lab_UT.dictrl.state_fast_3\ : std_logic;
signal bu_rx_data_2_rep2 : std_logic;
signal \Lab_UT.dictrl.N_15\ : std_logic;
signal \Lab_UT.dictrl.next_state12\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.N_21_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_0_1\ : std_logic;
signal \Lab_UT.dictrl.next_state18\ : std_logic;
signal bu_rx_data_1_rep2 : std_logic;
signal \Lab_UT.dictrl.g1_5_0\ : std_logic;
signal \Lab_UT.state_1\ : std_logic;
signal \Lab_UT.dictrl.N_23\ : std_logic;
signal \Lab_UT.dictrl.N_30\ : std_logic;
signal \Lab_UT.dictrl.next_state5_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state32Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_18\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep1\ : std_logic;
signal \Lab_UT.dictrl.m17_1\ : std_logic;
signal \Lab_UT.state_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z32\ : std_logic;
signal \Lab_UT.dictrl.N_29_0\ : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal \Lab_UT.dictrl.g1_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_6\ : std_logic;
signal \Lab_UT.dictrl.g1_0_0\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep2\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a3_3\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_3_rep2 : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_4 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_g : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal rst_g : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__10175\&\N__10151\&\N__10046\&\N__10079\&\N__10112\&\N__9923\&\N__10022\&\N__9989\&\N__9959\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__12251\&\N__14003\&\N__14021\&\N__11153\&\N__10931\&\N__11207\&\N__12398\&\N__10985\&\N__12236\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__12542\&'0'&\N__10226\&'0'&\N__10238\&'0'&\N__10217\&'0'&\N__12416\&'0'&\N__16823\&'0'&\N__10232\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__8588\,
            RESETB => \N__12671\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22354\,
            RE => \N__12664\,
            WCLKE => \N__10952\,
            WCLK => \N__22353\,
            WE => \N__10948\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23331\,
            DIN => \N__23330\,
            DOUT => \N__23329\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23331\,
            PADOUT => \N__23330\,
            PADIN => \N__23329\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23322\,
            DIN => \N__23321\,
            DOUT => \N__23320\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23322\,
            PADOUT => \N__23321\,
            PADIN => \N__23320\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23313\,
            DIN => \N__23312\,
            DOUT => \N__23311\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23313\,
            PADOUT => \N__23312\,
            PADIN => \N__23311\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__22321\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23304\,
            DIN => \N__23303\,
            DOUT => \N__23302\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__23304\,
            PADOUT => \N__23303\,
            PADIN => \N__23302\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23295\,
            DIN => \N__23294\,
            DOUT => \N__23293\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23295\,
            PADOUT => \N__23294\,
            PADIN => \N__23293\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23286\,
            DIN => \N__23285\,
            DOUT => \N__23284\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23286\,
            PADOUT => \N__23285\,
            PADIN => \N__23284\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23277\,
            DIN => \N__23276\,
            DOUT => \N__23275\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23277\,
            PADOUT => \N__23276\,
            PADIN => \N__23275\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23268\,
            DIN => \N__23267\,
            DOUT => \N__23266\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23268\,
            PADOUT => \N__23267\,
            PADIN => \N__23266\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9314\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23259\,
            DIN => \N__23258\,
            DOUT => \N__23257\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__23259\,
            PADOUT => \N__23258\,
            PADIN => \N__23257\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23250\,
            DIN => \N__23249\,
            DOUT => \N__23248\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__23250\,
            PADOUT => \N__23249\,
            PADIN => \N__23248\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__23231\,
            I => \Lab_UT.dictrl.g1_5_cascade_\
        );

    \I__5611\ : InMux
    port map (
            O => \N__23228\,
            I => \N__23225\
        );

    \I__5610\ : LocalMux
    port map (
            O => \N__23225\,
            I => \Lab_UT.dictrl.g1_6\
        );

    \I__5609\ : InMux
    port map (
            O => \N__23222\,
            I => \N__23219\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__23219\,
            I => \N__23216\
        );

    \I__5607\ : Span4Mux_h
    port map (
            O => \N__23216\,
            I => \N__23213\
        );

    \I__5606\ : Odrv4
    port map (
            O => \N__23213\,
            I => \Lab_UT.dictrl.g1_0_0\
        );

    \I__5605\ : InMux
    port map (
            O => \N__23210\,
            I => \N__23206\
        );

    \I__5604\ : InMux
    port map (
            O => \N__23209\,
            I => \N__23199\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23206\,
            I => \N__23189\
        );

    \I__5602\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23182\
        );

    \I__5601\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23182\
        );

    \I__5600\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23182\
        );

    \I__5599\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23178\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23175\
        );

    \I__5597\ : CascadeMux
    port map (
            O => \N__23198\,
            I => \N__23171\
        );

    \I__5596\ : CascadeMux
    port map (
            O => \N__23197\,
            I => \N__23167\
        );

    \I__5595\ : InMux
    port map (
            O => \N__23196\,
            I => \N__23160\
        );

    \I__5594\ : InMux
    port map (
            O => \N__23195\,
            I => \N__23160\
        );

    \I__5593\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23160\
        );

    \I__5592\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23155\
        );

    \I__5591\ : InMux
    port map (
            O => \N__23192\,
            I => \N__23155\
        );

    \I__5590\ : Span4Mux_h
    port map (
            O => \N__23189\,
            I => \N__23150\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__23182\,
            I => \N__23150\
        );

    \I__5588\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23147\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__23178\,
            I => \N__23144\
        );

    \I__5586\ : Span4Mux_v
    port map (
            O => \N__23175\,
            I => \N__23141\
        );

    \I__5585\ : InMux
    port map (
            O => \N__23174\,
            I => \N__23138\
        );

    \I__5584\ : InMux
    port map (
            O => \N__23171\,
            I => \N__23135\
        );

    \I__5583\ : InMux
    port map (
            O => \N__23170\,
            I => \N__23130\
        );

    \I__5582\ : InMux
    port map (
            O => \N__23167\,
            I => \N__23130\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23160\,
            I => \N__23125\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23125\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__23150\,
            I => \N__23122\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23147\,
            I => \N__23117\
        );

    \I__5577\ : Span4Mux_h
    port map (
            O => \N__23144\,
            I => \N__23117\
        );

    \I__5576\ : Span4Mux_h
    port map (
            O => \N__23141\,
            I => \N__23108\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__23138\,
            I => \N__23108\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23108\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__23130\,
            I => \N__23108\
        );

    \I__5572\ : Span12Mux_s10_h
    port map (
            O => \N__23125\,
            I => \N__23105\
        );

    \I__5571\ : Odrv4
    port map (
            O => \N__23122\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__5570\ : Odrv4
    port map (
            O => \N__23117\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__5569\ : Odrv4
    port map (
            O => \N__23108\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__5568\ : Odrv12
    port map (
            O => \N__23105\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__5567\ : InMux
    port map (
            O => \N__23096\,
            I => \N__23093\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__23093\,
            I => \N__23090\
        );

    \I__5565\ : Odrv4
    port map (
            O => \N__23090\,
            I => \Lab_UT.dictrl.g0_i_a3_3\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__23087\,
            I => \N__23080\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__23086\,
            I => \N__23074\
        );

    \I__5562\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23069\
        );

    \I__5561\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23066\
        );

    \I__5560\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23061\
        );

    \I__5559\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23061\
        );

    \I__5558\ : InMux
    port map (
            O => \N__23079\,
            I => \N__23058\
        );

    \I__5557\ : InMux
    port map (
            O => \N__23078\,
            I => \N__23055\
        );

    \I__5556\ : InMux
    port map (
            O => \N__23077\,
            I => \N__23052\
        );

    \I__5555\ : InMux
    port map (
            O => \N__23074\,
            I => \N__23047\
        );

    \I__5554\ : InMux
    port map (
            O => \N__23073\,
            I => \N__23047\
        );

    \I__5553\ : InMux
    port map (
            O => \N__23072\,
            I => \N__23042\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__23069\,
            I => \N__23035\
        );

    \I__5551\ : LocalMux
    port map (
            O => \N__23066\,
            I => \N__23035\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23035\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__23058\,
            I => \N__23030\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__23055\,
            I => \N__23025\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23025\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__23047\,
            I => \N__23022\
        );

    \I__5545\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23017\
        );

    \I__5544\ : InMux
    port map (
            O => \N__23045\,
            I => \N__23017\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__23042\,
            I => \N__23014\
        );

    \I__5542\ : Span4Mux_v
    port map (
            O => \N__23035\,
            I => \N__23011\
        );

    \I__5541\ : InMux
    port map (
            O => \N__23034\,
            I => \N__23008\
        );

    \I__5540\ : InMux
    port map (
            O => \N__23033\,
            I => \N__23005\
        );

    \I__5539\ : Span4Mux_v
    port map (
            O => \N__23030\,
            I => \N__23002\
        );

    \I__5538\ : Span4Mux_h
    port map (
            O => \N__23025\,
            I => \N__22999\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__23022\,
            I => \N__22994\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__22994\
        );

    \I__5535\ : Span4Mux_s2_v
    port map (
            O => \N__23014\,
            I => \N__22989\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__23011\,
            I => \N__22989\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23008\,
            I => bu_rx_data_7
        );

    \I__5532\ : LocalMux
    port map (
            O => \N__23005\,
            I => bu_rx_data_7
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__23002\,
            I => bu_rx_data_7
        );

    \I__5530\ : Odrv4
    port map (
            O => \N__22999\,
            I => bu_rx_data_7
        );

    \I__5529\ : Odrv4
    port map (
            O => \N__22994\,
            I => bu_rx_data_7
        );

    \I__5528\ : Odrv4
    port map (
            O => \N__22989\,
            I => bu_rx_data_7
        );

    \I__5527\ : InMux
    port map (
            O => \N__22976\,
            I => \N__22966\
        );

    \I__5526\ : CascadeMux
    port map (
            O => \N__22975\,
            I => \N__22962\
        );

    \I__5525\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22956\
        );

    \I__5524\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22953\
        );

    \I__5523\ : CascadeMux
    port map (
            O => \N__22972\,
            I => \N__22949\
        );

    \I__5522\ : CascadeMux
    port map (
            O => \N__22971\,
            I => \N__22946\
        );

    \I__5521\ : InMux
    port map (
            O => \N__22970\,
            I => \N__22941\
        );

    \I__5520\ : InMux
    port map (
            O => \N__22969\,
            I => \N__22941\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__22966\,
            I => \N__22938\
        );

    \I__5518\ : InMux
    port map (
            O => \N__22965\,
            I => \N__22933\
        );

    \I__5517\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22933\
        );

    \I__5516\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22930\
        );

    \I__5515\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22925\
        );

    \I__5514\ : InMux
    port map (
            O => \N__22959\,
            I => \N__22925\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__22956\,
            I => \N__22920\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__22953\,
            I => \N__22920\
        );

    \I__5511\ : InMux
    port map (
            O => \N__22952\,
            I => \N__22917\
        );

    \I__5510\ : InMux
    port map (
            O => \N__22949\,
            I => \N__22914\
        );

    \I__5509\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22911\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__22941\,
            I => \N__22904\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__22938\,
            I => \N__22904\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__22933\,
            I => \N__22904\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22901\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__22925\,
            I => \N__22898\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__22920\,
            I => \N__22895\
        );

    \I__5502\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22886\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22886\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__22911\,
            I => \N__22886\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__22904\,
            I => \N__22886\
        );

    \I__5498\ : Odrv4
    port map (
            O => \N__22901\,
            I => bu_rx_data_3_rep2
        );

    \I__5497\ : Odrv4
    port map (
            O => \N__22898\,
            I => bu_rx_data_3_rep2
        );

    \I__5496\ : Odrv4
    port map (
            O => \N__22895\,
            I => bu_rx_data_3_rep2
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__22886\,
            I => bu_rx_data_3_rep2
        );

    \I__5494\ : InMux
    port map (
            O => \N__22877\,
            I => \N__22872\
        );

    \I__5493\ : InMux
    port map (
            O => \N__22876\,
            I => \N__22866\
        );

    \I__5492\ : CascadeMux
    port map (
            O => \N__22875\,
            I => \N__22859\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__22872\,
            I => \N__22856\
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__22871\,
            I => \N__22853\
        );

    \I__5489\ : InMux
    port map (
            O => \N__22870\,
            I => \N__22848\
        );

    \I__5488\ : InMux
    port map (
            O => \N__22869\,
            I => \N__22848\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22845\
        );

    \I__5486\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22842\
        );

    \I__5485\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22839\
        );

    \I__5484\ : InMux
    port map (
            O => \N__22863\,
            I => \N__22834\
        );

    \I__5483\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22834\
        );

    \I__5482\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22831\
        );

    \I__5481\ : Span4Mux_s2_h
    port map (
            O => \N__22856\,
            I => \N__22828\
        );

    \I__5480\ : InMux
    port map (
            O => \N__22853\,
            I => \N__22821\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__22848\,
            I => \N__22814\
        );

    \I__5478\ : Span4Mux_h
    port map (
            O => \N__22845\,
            I => \N__22814\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N__22814\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__22839\,
            I => \N__22809\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__22834\,
            I => \N__22809\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__22831\,
            I => \N__22804\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__22828\,
            I => \N__22804\
        );

    \I__5472\ : InMux
    port map (
            O => \N__22827\,
            I => \N__22801\
        );

    \I__5471\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22798\
        );

    \I__5470\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22793\
        );

    \I__5469\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22793\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__22821\,
            I => \N__22788\
        );

    \I__5467\ : Span4Mux_h
    port map (
            O => \N__22814\,
            I => \N__22788\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__22809\,
            I => \N__22785\
        );

    \I__5465\ : Span4Mux_h
    port map (
            O => \N__22804\,
            I => \N__22782\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__22801\,
            I => bu_rx_data_6
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__22798\,
            I => bu_rx_data_6
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__22793\,
            I => bu_rx_data_6
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__22788\,
            I => bu_rx_data_6
        );

    \I__5460\ : Odrv4
    port map (
            O => \N__22785\,
            I => bu_rx_data_6
        );

    \I__5459\ : Odrv4
    port map (
            O => \N__22782\,
            I => bu_rx_data_6
        );

    \I__5458\ : InMux
    port map (
            O => \N__22769\,
            I => \N__22761\
        );

    \I__5457\ : InMux
    port map (
            O => \N__22768\,
            I => \N__22756\
        );

    \I__5456\ : InMux
    port map (
            O => \N__22767\,
            I => \N__22752\
        );

    \I__5455\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22749\
        );

    \I__5454\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22744\
        );

    \I__5453\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22738\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__22761\,
            I => \N__22733\
        );

    \I__5451\ : InMux
    port map (
            O => \N__22760\,
            I => \N__22728\
        );

    \I__5450\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22728\
        );

    \I__5449\ : LocalMux
    port map (
            O => \N__22756\,
            I => \N__22724\
        );

    \I__5448\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22721\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__22752\,
            I => \N__22716\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__22749\,
            I => \N__22716\
        );

    \I__5445\ : InMux
    port map (
            O => \N__22748\,
            I => \N__22713\
        );

    \I__5444\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22710\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__22744\,
            I => \N__22707\
        );

    \I__5442\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22702\
        );

    \I__5441\ : InMux
    port map (
            O => \N__22742\,
            I => \N__22697\
        );

    \I__5440\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22697\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__22738\,
            I => \N__22694\
        );

    \I__5438\ : InMux
    port map (
            O => \N__22737\,
            I => \N__22691\
        );

    \I__5437\ : InMux
    port map (
            O => \N__22736\,
            I => \N__22688\
        );

    \I__5436\ : Span4Mux_s3_v
    port map (
            O => \N__22733\,
            I => \N__22685\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__22728\,
            I => \N__22682\
        );

    \I__5434\ : InMux
    port map (
            O => \N__22727\,
            I => \N__22679\
        );

    \I__5433\ : Span4Mux_v
    port map (
            O => \N__22724\,
            I => \N__22672\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__22721\,
            I => \N__22672\
        );

    \I__5431\ : Span4Mux_v
    port map (
            O => \N__22716\,
            I => \N__22672\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22713\,
            I => \N__22665\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__22710\,
            I => \N__22665\
        );

    \I__5428\ : Span4Mux_v
    port map (
            O => \N__22707\,
            I => \N__22665\
        );

    \I__5427\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22660\
        );

    \I__5426\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22660\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__22702\,
            I => \N__22655\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__22697\,
            I => \N__22655\
        );

    \I__5423\ : Span4Mux_s2_h
    port map (
            O => \N__22694\,
            I => \N__22652\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22647\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__22688\,
            I => \N__22647\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__22685\,
            I => \N__22642\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__22682\,
            I => \N__22642\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22635\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__22672\,
            I => \N__22635\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__22665\,
            I => \N__22635\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__22660\,
            I => \N__22630\
        );

    \I__5414\ : Span4Mux_h
    port map (
            O => \N__22655\,
            I => \N__22630\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__22652\,
            I => \N__22627\
        );

    \I__5412\ : Odrv12
    port map (
            O => \N__22647\,
            I => bu_rx_data_1
        );

    \I__5411\ : Odrv4
    port map (
            O => \N__22642\,
            I => bu_rx_data_1
        );

    \I__5410\ : Odrv4
    port map (
            O => \N__22635\,
            I => bu_rx_data_1
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__22630\,
            I => bu_rx_data_1
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__22627\,
            I => bu_rx_data_1
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__22616\,
            I => \N__22612\
        );

    \I__5406\ : CascadeMux
    port map (
            O => \N__22615\,
            I => \N__22606\
        );

    \I__5405\ : InMux
    port map (
            O => \N__22612\,
            I => \N__22603\
        );

    \I__5404\ : CascadeMux
    port map (
            O => \N__22611\,
            I => \N__22600\
        );

    \I__5403\ : InMux
    port map (
            O => \N__22610\,
            I => \N__22592\
        );

    \I__5402\ : InMux
    port map (
            O => \N__22609\,
            I => \N__22592\
        );

    \I__5401\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22592\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22603\,
            I => \N__22589\
        );

    \I__5399\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22586\
        );

    \I__5398\ : InMux
    port map (
            O => \N__22599\,
            I => \N__22583\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__22592\,
            I => \N__22580\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__22589\,
            I => \N__22577\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22574\
        );

    \I__5394\ : LocalMux
    port map (
            O => \N__22583\,
            I => \N__22571\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__22580\,
            I => \N__22568\
        );

    \I__5392\ : Odrv4
    port map (
            O => \N__22577\,
            I => bu_rx_data_0_rep1
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__22574\,
            I => bu_rx_data_0_rep1
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__22571\,
            I => bu_rx_data_0_rep1
        );

    \I__5389\ : Odrv4
    port map (
            O => \N__22568\,
            I => bu_rx_data_0_rep1
        );

    \I__5388\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22553\
        );

    \I__5387\ : InMux
    port map (
            O => \N__22558\,
            I => \N__22550\
        );

    \I__5386\ : CascadeMux
    port map (
            O => \N__22557\,
            I => \N__22547\
        );

    \I__5385\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22541\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22536\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__22550\,
            I => \N__22536\
        );

    \I__5382\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22533\
        );

    \I__5381\ : InMux
    port map (
            O => \N__22546\,
            I => \N__22528\
        );

    \I__5380\ : InMux
    port map (
            O => \N__22545\,
            I => \N__22524\
        );

    \I__5379\ : InMux
    port map (
            O => \N__22544\,
            I => \N__22521\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__22541\,
            I => \N__22513\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__22536\,
            I => \N__22513\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22513\
        );

    \I__5375\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22508\
        );

    \I__5374\ : InMux
    port map (
            O => \N__22531\,
            I => \N__22508\
        );

    \I__5373\ : LocalMux
    port map (
            O => \N__22528\,
            I => \N__22505\
        );

    \I__5372\ : InMux
    port map (
            O => \N__22527\,
            I => \N__22499\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__22524\,
            I => \N__22494\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__22521\,
            I => \N__22494\
        );

    \I__5369\ : InMux
    port map (
            O => \N__22520\,
            I => \N__22491\
        );

    \I__5368\ : Span4Mux_h
    port map (
            O => \N__22513\,
            I => \N__22488\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22483\
        );

    \I__5366\ : Span12Mux_v
    port map (
            O => \N__22505\,
            I => \N__22483\
        );

    \I__5365\ : InMux
    port map (
            O => \N__22504\,
            I => \N__22476\
        );

    \I__5364\ : InMux
    port map (
            O => \N__22503\,
            I => \N__22476\
        );

    \I__5363\ : InMux
    port map (
            O => \N__22502\,
            I => \N__22476\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__22499\,
            I => \N__22471\
        );

    \I__5361\ : Span4Mux_s3_v
    port map (
            O => \N__22494\,
            I => \N__22471\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22491\,
            I => bu_rx_data_5
        );

    \I__5359\ : Odrv4
    port map (
            O => \N__22488\,
            I => bu_rx_data_5
        );

    \I__5358\ : Odrv12
    port map (
            O => \N__22483\,
            I => bu_rx_data_5
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__22476\,
            I => bu_rx_data_5
        );

    \I__5356\ : Odrv4
    port map (
            O => \N__22471\,
            I => bu_rx_data_5
        );

    \I__5355\ : InMux
    port map (
            O => \N__22460\,
            I => \N__22452\
        );

    \I__5354\ : InMux
    port map (
            O => \N__22459\,
            I => \N__22446\
        );

    \I__5353\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22443\
        );

    \I__5352\ : InMux
    port map (
            O => \N__22457\,
            I => \N__22440\
        );

    \I__5351\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22437\
        );

    \I__5350\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22431\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__22452\,
            I => \N__22427\
        );

    \I__5348\ : InMux
    port map (
            O => \N__22451\,
            I => \N__22420\
        );

    \I__5347\ : InMux
    port map (
            O => \N__22450\,
            I => \N__22420\
        );

    \I__5346\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22420\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__22446\,
            I => \N__22416\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22443\,
            I => \N__22409\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22440\,
            I => \N__22409\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__22437\,
            I => \N__22409\
        );

    \I__5341\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22402\
        );

    \I__5340\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22402\
        );

    \I__5339\ : InMux
    port map (
            O => \N__22434\,
            I => \N__22402\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__22431\,
            I => \N__22399\
        );

    \I__5337\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22396\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__22427\,
            I => \N__22391\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22420\,
            I => \N__22391\
        );

    \I__5334\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22388\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__22416\,
            I => \N__22385\
        );

    \I__5332\ : Span4Mux_h
    port map (
            O => \N__22409\,
            I => \N__22380\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__22402\,
            I => \N__22380\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__22399\,
            I => \N__22375\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22396\,
            I => \N__22375\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__22391\,
            I => \N__22372\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__22388\,
            I => bu_rx_data_4
        );

    \I__5326\ : Odrv4
    port map (
            O => \N__22385\,
            I => bu_rx_data_4
        );

    \I__5325\ : Odrv4
    port map (
            O => \N__22380\,
            I => bu_rx_data_4
        );

    \I__5324\ : Odrv4
    port map (
            O => \N__22375\,
            I => bu_rx_data_4
        );

    \I__5323\ : Odrv4
    port map (
            O => \N__22372\,
            I => bu_rx_data_4
        );

    \I__5322\ : ClkMux
    port map (
            O => \N__22361\,
            I => \N__22082\
        );

    \I__5321\ : ClkMux
    port map (
            O => \N__22360\,
            I => \N__22082\
        );

    \I__5320\ : ClkMux
    port map (
            O => \N__22359\,
            I => \N__22082\
        );

    \I__5319\ : ClkMux
    port map (
            O => \N__22358\,
            I => \N__22082\
        );

    \I__5318\ : ClkMux
    port map (
            O => \N__22357\,
            I => \N__22082\
        );

    \I__5317\ : ClkMux
    port map (
            O => \N__22356\,
            I => \N__22082\
        );

    \I__5316\ : ClkMux
    port map (
            O => \N__22355\,
            I => \N__22082\
        );

    \I__5315\ : ClkMux
    port map (
            O => \N__22354\,
            I => \N__22082\
        );

    \I__5314\ : ClkMux
    port map (
            O => \N__22353\,
            I => \N__22082\
        );

    \I__5313\ : ClkMux
    port map (
            O => \N__22352\,
            I => \N__22082\
        );

    \I__5312\ : ClkMux
    port map (
            O => \N__22351\,
            I => \N__22082\
        );

    \I__5311\ : ClkMux
    port map (
            O => \N__22350\,
            I => \N__22082\
        );

    \I__5310\ : ClkMux
    port map (
            O => \N__22349\,
            I => \N__22082\
        );

    \I__5309\ : ClkMux
    port map (
            O => \N__22348\,
            I => \N__22082\
        );

    \I__5308\ : ClkMux
    port map (
            O => \N__22347\,
            I => \N__22082\
        );

    \I__5307\ : ClkMux
    port map (
            O => \N__22346\,
            I => \N__22082\
        );

    \I__5306\ : ClkMux
    port map (
            O => \N__22345\,
            I => \N__22082\
        );

    \I__5305\ : ClkMux
    port map (
            O => \N__22344\,
            I => \N__22082\
        );

    \I__5304\ : ClkMux
    port map (
            O => \N__22343\,
            I => \N__22082\
        );

    \I__5303\ : ClkMux
    port map (
            O => \N__22342\,
            I => \N__22082\
        );

    \I__5302\ : ClkMux
    port map (
            O => \N__22341\,
            I => \N__22082\
        );

    \I__5301\ : ClkMux
    port map (
            O => \N__22340\,
            I => \N__22082\
        );

    \I__5300\ : ClkMux
    port map (
            O => \N__22339\,
            I => \N__22082\
        );

    \I__5299\ : ClkMux
    port map (
            O => \N__22338\,
            I => \N__22082\
        );

    \I__5298\ : ClkMux
    port map (
            O => \N__22337\,
            I => \N__22082\
        );

    \I__5297\ : ClkMux
    port map (
            O => \N__22336\,
            I => \N__22082\
        );

    \I__5296\ : ClkMux
    port map (
            O => \N__22335\,
            I => \N__22082\
        );

    \I__5295\ : ClkMux
    port map (
            O => \N__22334\,
            I => \N__22082\
        );

    \I__5294\ : ClkMux
    port map (
            O => \N__22333\,
            I => \N__22082\
        );

    \I__5293\ : ClkMux
    port map (
            O => \N__22332\,
            I => \N__22082\
        );

    \I__5292\ : ClkMux
    port map (
            O => \N__22331\,
            I => \N__22082\
        );

    \I__5291\ : ClkMux
    port map (
            O => \N__22330\,
            I => \N__22082\
        );

    \I__5290\ : ClkMux
    port map (
            O => \N__22329\,
            I => \N__22082\
        );

    \I__5289\ : ClkMux
    port map (
            O => \N__22328\,
            I => \N__22082\
        );

    \I__5288\ : ClkMux
    port map (
            O => \N__22327\,
            I => \N__22082\
        );

    \I__5287\ : ClkMux
    port map (
            O => \N__22326\,
            I => \N__22082\
        );

    \I__5286\ : ClkMux
    port map (
            O => \N__22325\,
            I => \N__22082\
        );

    \I__5285\ : ClkMux
    port map (
            O => \N__22324\,
            I => \N__22082\
        );

    \I__5284\ : ClkMux
    port map (
            O => \N__22323\,
            I => \N__22082\
        );

    \I__5283\ : ClkMux
    port map (
            O => \N__22322\,
            I => \N__22082\
        );

    \I__5282\ : ClkMux
    port map (
            O => \N__22321\,
            I => \N__22082\
        );

    \I__5281\ : ClkMux
    port map (
            O => \N__22320\,
            I => \N__22082\
        );

    \I__5280\ : ClkMux
    port map (
            O => \N__22319\,
            I => \N__22082\
        );

    \I__5279\ : ClkMux
    port map (
            O => \N__22318\,
            I => \N__22082\
        );

    \I__5278\ : ClkMux
    port map (
            O => \N__22317\,
            I => \N__22082\
        );

    \I__5277\ : ClkMux
    port map (
            O => \N__22316\,
            I => \N__22082\
        );

    \I__5276\ : ClkMux
    port map (
            O => \N__22315\,
            I => \N__22082\
        );

    \I__5275\ : ClkMux
    port map (
            O => \N__22314\,
            I => \N__22082\
        );

    \I__5274\ : ClkMux
    port map (
            O => \N__22313\,
            I => \N__22082\
        );

    \I__5273\ : ClkMux
    port map (
            O => \N__22312\,
            I => \N__22082\
        );

    \I__5272\ : ClkMux
    port map (
            O => \N__22311\,
            I => \N__22082\
        );

    \I__5271\ : ClkMux
    port map (
            O => \N__22310\,
            I => \N__22082\
        );

    \I__5270\ : ClkMux
    port map (
            O => \N__22309\,
            I => \N__22082\
        );

    \I__5269\ : ClkMux
    port map (
            O => \N__22308\,
            I => \N__22082\
        );

    \I__5268\ : ClkMux
    port map (
            O => \N__22307\,
            I => \N__22082\
        );

    \I__5267\ : ClkMux
    port map (
            O => \N__22306\,
            I => \N__22082\
        );

    \I__5266\ : ClkMux
    port map (
            O => \N__22305\,
            I => \N__22082\
        );

    \I__5265\ : ClkMux
    port map (
            O => \N__22304\,
            I => \N__22082\
        );

    \I__5264\ : ClkMux
    port map (
            O => \N__22303\,
            I => \N__22082\
        );

    \I__5263\ : ClkMux
    port map (
            O => \N__22302\,
            I => \N__22082\
        );

    \I__5262\ : ClkMux
    port map (
            O => \N__22301\,
            I => \N__22082\
        );

    \I__5261\ : ClkMux
    port map (
            O => \N__22300\,
            I => \N__22082\
        );

    \I__5260\ : ClkMux
    port map (
            O => \N__22299\,
            I => \N__22082\
        );

    \I__5259\ : ClkMux
    port map (
            O => \N__22298\,
            I => \N__22082\
        );

    \I__5258\ : ClkMux
    port map (
            O => \N__22297\,
            I => \N__22082\
        );

    \I__5257\ : ClkMux
    port map (
            O => \N__22296\,
            I => \N__22082\
        );

    \I__5256\ : ClkMux
    port map (
            O => \N__22295\,
            I => \N__22082\
        );

    \I__5255\ : ClkMux
    port map (
            O => \N__22294\,
            I => \N__22082\
        );

    \I__5254\ : ClkMux
    port map (
            O => \N__22293\,
            I => \N__22082\
        );

    \I__5253\ : ClkMux
    port map (
            O => \N__22292\,
            I => \N__22082\
        );

    \I__5252\ : ClkMux
    port map (
            O => \N__22291\,
            I => \N__22082\
        );

    \I__5251\ : ClkMux
    port map (
            O => \N__22290\,
            I => \N__22082\
        );

    \I__5250\ : ClkMux
    port map (
            O => \N__22289\,
            I => \N__22082\
        );

    \I__5249\ : ClkMux
    port map (
            O => \N__22288\,
            I => \N__22082\
        );

    \I__5248\ : ClkMux
    port map (
            O => \N__22287\,
            I => \N__22082\
        );

    \I__5247\ : ClkMux
    port map (
            O => \N__22286\,
            I => \N__22082\
        );

    \I__5246\ : ClkMux
    port map (
            O => \N__22285\,
            I => \N__22082\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__22284\,
            I => \N__22082\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__22283\,
            I => \N__22082\
        );

    \I__5243\ : ClkMux
    port map (
            O => \N__22282\,
            I => \N__22082\
        );

    \I__5242\ : ClkMux
    port map (
            O => \N__22281\,
            I => \N__22082\
        );

    \I__5241\ : ClkMux
    port map (
            O => \N__22280\,
            I => \N__22082\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__22279\,
            I => \N__22082\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__22278\,
            I => \N__22082\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__22277\,
            I => \N__22082\
        );

    \I__5237\ : ClkMux
    port map (
            O => \N__22276\,
            I => \N__22082\
        );

    \I__5236\ : ClkMux
    port map (
            O => \N__22275\,
            I => \N__22082\
        );

    \I__5235\ : ClkMux
    port map (
            O => \N__22274\,
            I => \N__22082\
        );

    \I__5234\ : ClkMux
    port map (
            O => \N__22273\,
            I => \N__22082\
        );

    \I__5233\ : ClkMux
    port map (
            O => \N__22272\,
            I => \N__22082\
        );

    \I__5232\ : ClkMux
    port map (
            O => \N__22271\,
            I => \N__22082\
        );

    \I__5231\ : ClkMux
    port map (
            O => \N__22270\,
            I => \N__22082\
        );

    \I__5230\ : ClkMux
    port map (
            O => \N__22269\,
            I => \N__22082\
        );

    \I__5229\ : GlobalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__5228\ : gio2CtrlBuf
    port map (
            O => \N__22079\,
            I => clk_g
        );

    \I__5227\ : CEMux
    port map (
            O => \N__22076\,
            I => \N__22046\
        );

    \I__5226\ : CEMux
    port map (
            O => \N__22075\,
            I => \N__22046\
        );

    \I__5225\ : CEMux
    port map (
            O => \N__22074\,
            I => \N__22046\
        );

    \I__5224\ : CEMux
    port map (
            O => \N__22073\,
            I => \N__22046\
        );

    \I__5223\ : CEMux
    port map (
            O => \N__22072\,
            I => \N__22046\
        );

    \I__5222\ : CEMux
    port map (
            O => \N__22071\,
            I => \N__22046\
        );

    \I__5221\ : CEMux
    port map (
            O => \N__22070\,
            I => \N__22046\
        );

    \I__5220\ : CEMux
    port map (
            O => \N__22069\,
            I => \N__22046\
        );

    \I__5219\ : CEMux
    port map (
            O => \N__22068\,
            I => \N__22046\
        );

    \I__5218\ : CEMux
    port map (
            O => \N__22067\,
            I => \N__22046\
        );

    \I__5217\ : GlobalMux
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__5216\ : gio2CtrlBuf
    port map (
            O => \N__22043\,
            I => \buart.Z_rx.sample_g\
        );

    \I__5215\ : InMux
    port map (
            O => \N__22040\,
            I => \N__22031\
        );

    \I__5214\ : InMux
    port map (
            O => \N__22039\,
            I => \N__22028\
        );

    \I__5213\ : InMux
    port map (
            O => \N__22038\,
            I => \N__22025\
        );

    \I__5212\ : InMux
    port map (
            O => \N__22037\,
            I => \N__22022\
        );

    \I__5211\ : InMux
    port map (
            O => \N__22036\,
            I => \N__22019\
        );

    \I__5210\ : SRMux
    port map (
            O => \N__22035\,
            I => \N__22014\
        );

    \I__5209\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22014\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__22031\,
            I => \N__21966\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__21963\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__22025\,
            I => \N__21960\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22022\,
            I => \N__21957\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__22019\,
            I => \N__21954\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__22014\,
            I => \N__21935\
        );

    \I__5202\ : SRMux
    port map (
            O => \N__22013\,
            I => \N__21800\
        );

    \I__5201\ : SRMux
    port map (
            O => \N__22012\,
            I => \N__21800\
        );

    \I__5200\ : SRMux
    port map (
            O => \N__22011\,
            I => \N__21800\
        );

    \I__5199\ : SRMux
    port map (
            O => \N__22010\,
            I => \N__21800\
        );

    \I__5198\ : SRMux
    port map (
            O => \N__22009\,
            I => \N__21800\
        );

    \I__5197\ : SRMux
    port map (
            O => \N__22008\,
            I => \N__21800\
        );

    \I__5196\ : SRMux
    port map (
            O => \N__22007\,
            I => \N__21800\
        );

    \I__5195\ : SRMux
    port map (
            O => \N__22006\,
            I => \N__21800\
        );

    \I__5194\ : SRMux
    port map (
            O => \N__22005\,
            I => \N__21800\
        );

    \I__5193\ : SRMux
    port map (
            O => \N__22004\,
            I => \N__21800\
        );

    \I__5192\ : SRMux
    port map (
            O => \N__22003\,
            I => \N__21800\
        );

    \I__5191\ : SRMux
    port map (
            O => \N__22002\,
            I => \N__21800\
        );

    \I__5190\ : SRMux
    port map (
            O => \N__22001\,
            I => \N__21800\
        );

    \I__5189\ : SRMux
    port map (
            O => \N__22000\,
            I => \N__21800\
        );

    \I__5188\ : SRMux
    port map (
            O => \N__21999\,
            I => \N__21800\
        );

    \I__5187\ : SRMux
    port map (
            O => \N__21998\,
            I => \N__21800\
        );

    \I__5186\ : SRMux
    port map (
            O => \N__21997\,
            I => \N__21800\
        );

    \I__5185\ : SRMux
    port map (
            O => \N__21996\,
            I => \N__21800\
        );

    \I__5184\ : SRMux
    port map (
            O => \N__21995\,
            I => \N__21800\
        );

    \I__5183\ : SRMux
    port map (
            O => \N__21994\,
            I => \N__21800\
        );

    \I__5182\ : SRMux
    port map (
            O => \N__21993\,
            I => \N__21800\
        );

    \I__5181\ : SRMux
    port map (
            O => \N__21992\,
            I => \N__21800\
        );

    \I__5180\ : SRMux
    port map (
            O => \N__21991\,
            I => \N__21800\
        );

    \I__5179\ : SRMux
    port map (
            O => \N__21990\,
            I => \N__21800\
        );

    \I__5178\ : SRMux
    port map (
            O => \N__21989\,
            I => \N__21800\
        );

    \I__5177\ : SRMux
    port map (
            O => \N__21988\,
            I => \N__21800\
        );

    \I__5176\ : SRMux
    port map (
            O => \N__21987\,
            I => \N__21800\
        );

    \I__5175\ : SRMux
    port map (
            O => \N__21986\,
            I => \N__21800\
        );

    \I__5174\ : SRMux
    port map (
            O => \N__21985\,
            I => \N__21800\
        );

    \I__5173\ : SRMux
    port map (
            O => \N__21984\,
            I => \N__21800\
        );

    \I__5172\ : SRMux
    port map (
            O => \N__21983\,
            I => \N__21800\
        );

    \I__5171\ : SRMux
    port map (
            O => \N__21982\,
            I => \N__21800\
        );

    \I__5170\ : SRMux
    port map (
            O => \N__21981\,
            I => \N__21800\
        );

    \I__5169\ : SRMux
    port map (
            O => \N__21980\,
            I => \N__21800\
        );

    \I__5168\ : SRMux
    port map (
            O => \N__21979\,
            I => \N__21800\
        );

    \I__5167\ : SRMux
    port map (
            O => \N__21978\,
            I => \N__21800\
        );

    \I__5166\ : SRMux
    port map (
            O => \N__21977\,
            I => \N__21800\
        );

    \I__5165\ : SRMux
    port map (
            O => \N__21976\,
            I => \N__21800\
        );

    \I__5164\ : SRMux
    port map (
            O => \N__21975\,
            I => \N__21800\
        );

    \I__5163\ : SRMux
    port map (
            O => \N__21974\,
            I => \N__21800\
        );

    \I__5162\ : SRMux
    port map (
            O => \N__21973\,
            I => \N__21800\
        );

    \I__5161\ : SRMux
    port map (
            O => \N__21972\,
            I => \N__21800\
        );

    \I__5160\ : SRMux
    port map (
            O => \N__21971\,
            I => \N__21800\
        );

    \I__5159\ : SRMux
    port map (
            O => \N__21970\,
            I => \N__21800\
        );

    \I__5158\ : SRMux
    port map (
            O => \N__21969\,
            I => \N__21800\
        );

    \I__5157\ : Glb2LocalMux
    port map (
            O => \N__21966\,
            I => \N__21800\
        );

    \I__5156\ : Glb2LocalMux
    port map (
            O => \N__21963\,
            I => \N__21800\
        );

    \I__5155\ : Glb2LocalMux
    port map (
            O => \N__21960\,
            I => \N__21800\
        );

    \I__5154\ : Glb2LocalMux
    port map (
            O => \N__21957\,
            I => \N__21800\
        );

    \I__5153\ : Glb2LocalMux
    port map (
            O => \N__21954\,
            I => \N__21800\
        );

    \I__5152\ : SRMux
    port map (
            O => \N__21953\,
            I => \N__21800\
        );

    \I__5151\ : SRMux
    port map (
            O => \N__21952\,
            I => \N__21800\
        );

    \I__5150\ : SRMux
    port map (
            O => \N__21951\,
            I => \N__21800\
        );

    \I__5149\ : SRMux
    port map (
            O => \N__21950\,
            I => \N__21800\
        );

    \I__5148\ : SRMux
    port map (
            O => \N__21949\,
            I => \N__21800\
        );

    \I__5147\ : SRMux
    port map (
            O => \N__21948\,
            I => \N__21800\
        );

    \I__5146\ : SRMux
    port map (
            O => \N__21947\,
            I => \N__21800\
        );

    \I__5145\ : SRMux
    port map (
            O => \N__21946\,
            I => \N__21800\
        );

    \I__5144\ : SRMux
    port map (
            O => \N__21945\,
            I => \N__21800\
        );

    \I__5143\ : SRMux
    port map (
            O => \N__21944\,
            I => \N__21800\
        );

    \I__5142\ : SRMux
    port map (
            O => \N__21943\,
            I => \N__21800\
        );

    \I__5141\ : SRMux
    port map (
            O => \N__21942\,
            I => \N__21800\
        );

    \I__5140\ : SRMux
    port map (
            O => \N__21941\,
            I => \N__21800\
        );

    \I__5139\ : SRMux
    port map (
            O => \N__21940\,
            I => \N__21800\
        );

    \I__5138\ : SRMux
    port map (
            O => \N__21939\,
            I => \N__21800\
        );

    \I__5137\ : SRMux
    port map (
            O => \N__21938\,
            I => \N__21800\
        );

    \I__5136\ : Glb2LocalMux
    port map (
            O => \N__21935\,
            I => \N__21800\
        );

    \I__5135\ : GlobalMux
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__5134\ : gio2CtrlBuf
    port map (
            O => \N__21797\,
            I => rst_g
        );

    \I__5133\ : CascadeMux
    port map (
            O => \N__21794\,
            I => \N__21787\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21793\,
            I => \N__21781\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__21792\,
            I => \N__21778\
        );

    \I__5130\ : CascadeMux
    port map (
            O => \N__21791\,
            I => \N__21769\
        );

    \I__5129\ : CascadeMux
    port map (
            O => \N__21790\,
            I => \N__21765\
        );

    \I__5128\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21754\
        );

    \I__5127\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21754\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21785\,
            I => \N__21754\
        );

    \I__5125\ : InMux
    port map (
            O => \N__21784\,
            I => \N__21754\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__21781\,
            I => \N__21749\
        );

    \I__5123\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21746\
        );

    \I__5122\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21741\
        );

    \I__5121\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21741\
        );

    \I__5120\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21729\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21729\
        );

    \I__5118\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21729\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21772\,
            I => \N__21729\
        );

    \I__5116\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21722\
        );

    \I__5115\ : InMux
    port map (
            O => \N__21768\,
            I => \N__21722\
        );

    \I__5114\ : InMux
    port map (
            O => \N__21765\,
            I => \N__21722\
        );

    \I__5113\ : InMux
    port map (
            O => \N__21764\,
            I => \N__21719\
        );

    \I__5112\ : CascadeMux
    port map (
            O => \N__21763\,
            I => \N__21714\
        );

    \I__5111\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21708\
        );

    \I__5110\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21705\
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__21752\,
            I => \N__21702\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__21749\,
            I => \N__21699\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__21746\,
            I => \N__21694\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21694\
        );

    \I__5105\ : InMux
    port map (
            O => \N__21740\,
            I => \N__21686\
        );

    \I__5104\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21686\
        );

    \I__5103\ : InMux
    port map (
            O => \N__21738\,
            I => \N__21686\
        );

    \I__5102\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21679\
        );

    \I__5101\ : LocalMux
    port map (
            O => \N__21722\,
            I => \N__21679\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21679\
        );

    \I__5099\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21674\
        );

    \I__5098\ : InMux
    port map (
            O => \N__21717\,
            I => \N__21674\
        );

    \I__5097\ : InMux
    port map (
            O => \N__21714\,
            I => \N__21665\
        );

    \I__5096\ : InMux
    port map (
            O => \N__21713\,
            I => \N__21665\
        );

    \I__5095\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21665\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21711\,
            I => \N__21665\
        );

    \I__5093\ : Span4Mux_h
    port map (
            O => \N__21708\,
            I => \N__21662\
        );

    \I__5092\ : LocalMux
    port map (
            O => \N__21705\,
            I => \N__21659\
        );

    \I__5091\ : InMux
    port map (
            O => \N__21702\,
            I => \N__21656\
        );

    \I__5090\ : Span4Mux_s3_h
    port map (
            O => \N__21699\,
            I => \N__21651\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__21694\,
            I => \N__21651\
        );

    \I__5088\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21648\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__21686\,
            I => \N__21645\
        );

    \I__5086\ : Span4Mux_v
    port map (
            O => \N__21679\,
            I => \N__21642\
        );

    \I__5085\ : LocalMux
    port map (
            O => \N__21674\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__21665\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5083\ : Odrv4
    port map (
            O => \N__21662\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5082\ : Odrv4
    port map (
            O => \N__21659\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5081\ : LocalMux
    port map (
            O => \N__21656\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__21651\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5079\ : LocalMux
    port map (
            O => \N__21648\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5078\ : Odrv4
    port map (
            O => \N__21645\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__21642\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__21623\,
            I => \Lab_UT.dictrl.N_21_cascade_\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21614\
        );

    \I__5074\ : InMux
    port map (
            O => \N__21619\,
            I => \N__21614\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__21611\,
            I => \N__21608\
        );

    \I__5071\ : Odrv4
    port map (
            O => \N__21608\,
            I => \Lab_UT.dictrl.next_state_latmux_0_1\
        );

    \I__5070\ : InMux
    port map (
            O => \N__21605\,
            I => \N__21598\
        );

    \I__5069\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21591\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21591\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21591\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21601\,
            I => \N__21588\
        );

    \I__5065\ : LocalMux
    port map (
            O => \N__21598\,
            I => \N__21583\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__21591\,
            I => \N__21583\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__21588\,
            I => \N__21580\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__21583\,
            I => \N__21577\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__21580\,
            I => \Lab_UT.dictrl.next_state18\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__21577\,
            I => \Lab_UT.dictrl.next_state18\
        );

    \I__5059\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21565\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__21571\,
            I => \N__21561\
        );

    \I__5057\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21556\
        );

    \I__5056\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21556\
        );

    \I__5055\ : InMux
    port map (
            O => \N__21568\,
            I => \N__21551\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21565\,
            I => \N__21548\
        );

    \I__5053\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21545\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21542\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__21556\,
            I => \N__21539\
        );

    \I__5050\ : InMux
    port map (
            O => \N__21555\,
            I => \N__21536\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__21554\,
            I => \N__21531\
        );

    \I__5048\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21527\
        );

    \I__5047\ : Span4Mux_h
    port map (
            O => \N__21548\,
            I => \N__21524\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__21545\,
            I => \N__21519\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__21542\,
            I => \N__21519\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__21539\,
            I => \N__21516\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21513\
        );

    \I__5042\ : InMux
    port map (
            O => \N__21535\,
            I => \N__21508\
        );

    \I__5041\ : InMux
    port map (
            O => \N__21534\,
            I => \N__21508\
        );

    \I__5040\ : InMux
    port map (
            O => \N__21531\,
            I => \N__21503\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21503\
        );

    \I__5038\ : Span4Mux_s2_h
    port map (
            O => \N__21527\,
            I => \N__21500\
        );

    \I__5037\ : Odrv4
    port map (
            O => \N__21524\,
            I => bu_rx_data_1_rep2
        );

    \I__5036\ : Odrv12
    port map (
            O => \N__21519\,
            I => bu_rx_data_1_rep2
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__21516\,
            I => bu_rx_data_1_rep2
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__21513\,
            I => bu_rx_data_1_rep2
        );

    \I__5033\ : LocalMux
    port map (
            O => \N__21508\,
            I => bu_rx_data_1_rep2
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21503\,
            I => bu_rx_data_1_rep2
        );

    \I__5031\ : Odrv4
    port map (
            O => \N__21500\,
            I => bu_rx_data_1_rep2
        );

    \I__5030\ : CascadeMux
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21476\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__21476\,
            I => \N__21473\
        );

    \I__5026\ : Odrv4
    port map (
            O => \N__21473\,
            I => \Lab_UT.dictrl.g1_5_0\
        );

    \I__5025\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21456\
        );

    \I__5024\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21456\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21456\
        );

    \I__5022\ : InMux
    port map (
            O => \N__21467\,
            I => \N__21456\
        );

    \I__5021\ : CascadeMux
    port map (
            O => \N__21466\,
            I => \N__21449\
        );

    \I__5020\ : InMux
    port map (
            O => \N__21465\,
            I => \N__21443\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__21456\,
            I => \N__21440\
        );

    \I__5018\ : InMux
    port map (
            O => \N__21455\,
            I => \N__21435\
        );

    \I__5017\ : InMux
    port map (
            O => \N__21454\,
            I => \N__21435\
        );

    \I__5016\ : InMux
    port map (
            O => \N__21453\,
            I => \N__21424\
        );

    \I__5015\ : InMux
    port map (
            O => \N__21452\,
            I => \N__21420\
        );

    \I__5014\ : InMux
    port map (
            O => \N__21449\,
            I => \N__21411\
        );

    \I__5013\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21411\
        );

    \I__5012\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21411\
        );

    \I__5011\ : InMux
    port map (
            O => \N__21446\,
            I => \N__21411\
        );

    \I__5010\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21406\
        );

    \I__5009\ : Span4Mux_v
    port map (
            O => \N__21440\,
            I => \N__21406\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__21435\,
            I => \N__21403\
        );

    \I__5007\ : InMux
    port map (
            O => \N__21434\,
            I => \N__21400\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__21433\,
            I => \N__21397\
        );

    \I__5005\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21392\
        );

    \I__5004\ : InMux
    port map (
            O => \N__21431\,
            I => \N__21392\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21430\,
            I => \N__21387\
        );

    \I__5002\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21387\
        );

    \I__5001\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21384\
        );

    \I__5000\ : InMux
    port map (
            O => \N__21427\,
            I => \N__21381\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21378\
        );

    \I__4998\ : CascadeMux
    port map (
            O => \N__21423\,
            I => \N__21370\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21366\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21356\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__21406\,
            I => \N__21356\
        );

    \I__4994\ : Span4Mux_v
    port map (
            O => \N__21403\,
            I => \N__21356\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21353\
        );

    \I__4992\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21350\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__21392\,
            I => \N__21347\
        );

    \I__4990\ : LocalMux
    port map (
            O => \N__21387\,
            I => \N__21340\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21384\,
            I => \N__21340\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21381\,
            I => \N__21340\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__21378\,
            I => \N__21337\
        );

    \I__4986\ : InMux
    port map (
            O => \N__21377\,
            I => \N__21334\
        );

    \I__4985\ : InMux
    port map (
            O => \N__21376\,
            I => \N__21323\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21323\
        );

    \I__4983\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21323\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21323\
        );

    \I__4981\ : InMux
    port map (
            O => \N__21370\,
            I => \N__21323\
        );

    \I__4980\ : InMux
    port map (
            O => \N__21369\,
            I => \N__21320\
        );

    \I__4979\ : Span4Mux_h
    port map (
            O => \N__21366\,
            I => \N__21317\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21365\,
            I => \N__21310\
        );

    \I__4977\ : InMux
    port map (
            O => \N__21364\,
            I => \N__21310\
        );

    \I__4976\ : InMux
    port map (
            O => \N__21363\,
            I => \N__21310\
        );

    \I__4975\ : Sp12to4
    port map (
            O => \N__21356\,
            I => \N__21307\
        );

    \I__4974\ : Span4Mux_s3_h
    port map (
            O => \N__21353\,
            I => \N__21296\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21350\,
            I => \N__21296\
        );

    \I__4972\ : Span4Mux_h
    port map (
            O => \N__21347\,
            I => \N__21296\
        );

    \I__4971\ : Span4Mux_h
    port map (
            O => \N__21340\,
            I => \N__21296\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__21337\,
            I => \N__21296\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21334\,
            I => \Lab_UT.state_1\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__21323\,
            I => \Lab_UT.state_1\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__21320\,
            I => \Lab_UT.state_1\
        );

    \I__4966\ : Odrv4
    port map (
            O => \N__21317\,
            I => \Lab_UT.state_1\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21310\,
            I => \Lab_UT.state_1\
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__21307\,
            I => \Lab_UT.state_1\
        );

    \I__4963\ : Odrv4
    port map (
            O => \N__21296\,
            I => \Lab_UT.state_1\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21281\,
            I => \N__21277\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21280\,
            I => \N__21274\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21277\,
            I => \Lab_UT.dictrl.N_23\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__21274\,
            I => \Lab_UT.dictrl.N_23\
        );

    \I__4958\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4957\ : LocalMux
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__4956\ : Span4Mux_h
    port map (
            O => \N__21263\,
            I => \N__21260\
        );

    \I__4955\ : Odrv4
    port map (
            O => \N__21260\,
            I => \Lab_UT.dictrl.N_30\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__21257\,
            I => \Lab_UT.dictrl.next_state5_3_cascade_\
        );

    \I__4953\ : InMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__4952\ : LocalMux
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__4951\ : Span4Mux_s2_h
    port map (
            O => \N__21248\,
            I => \N__21244\
        );

    \I__4950\ : InMux
    port map (
            O => \N__21247\,
            I => \N__21241\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__21244\,
            I => \Lab_UT.dictrl.next_state32Z0Z_1\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__21241\,
            I => \Lab_UT.dictrl.next_state32Z0Z_1\
        );

    \I__4947\ : CascadeMux
    port map (
            O => \N__21236\,
            I => \N__21232\
        );

    \I__4946\ : CascadeMux
    port map (
            O => \N__21235\,
            I => \N__21229\
        );

    \I__4945\ : InMux
    port map (
            O => \N__21232\,
            I => \N__21224\
        );

    \I__4944\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21224\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4941\ : Sp12to4
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4940\ : Odrv12
    port map (
            O => \N__21215\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__4939\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21203\
        );

    \I__4938\ : InMux
    port map (
            O => \N__21211\,
            I => \N__21203\
        );

    \I__4937\ : InMux
    port map (
            O => \N__21210\,
            I => \N__21199\
        );

    \I__4936\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21195\
        );

    \I__4935\ : InMux
    port map (
            O => \N__21208\,
            I => \N__21192\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__21203\,
            I => \N__21189\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21186\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21183\
        );

    \I__4931\ : CascadeMux
    port map (
            O => \N__21198\,
            I => \N__21179\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__21195\,
            I => \N__21174\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__21192\,
            I => \N__21174\
        );

    \I__4928\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21169\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__21186\,
            I => \N__21169\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__21183\,
            I => \N__21166\
        );

    \I__4925\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21163\
        );

    \I__4924\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21160\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__21174\,
            I => \N__21157\
        );

    \I__4922\ : Span4Mux_h
    port map (
            O => \N__21169\,
            I => \N__21154\
        );

    \I__4921\ : Sp12to4
    port map (
            O => \N__21166\,
            I => \N__21147\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21147\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__21160\,
            I => \N__21147\
        );

    \I__4918\ : Odrv4
    port map (
            O => \N__21157\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__21154\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__4916\ : Odrv12
    port map (
            O => \N__21147\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__4915\ : InMux
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__21137\,
            I => \Lab_UT.dictrl.m17_1\
        );

    \I__4913\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21118\
        );

    \I__4912\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21118\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__21132\,
            I => \N__21115\
        );

    \I__4910\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21105\
        );

    \I__4909\ : InMux
    port map (
            O => \N__21130\,
            I => \N__21100\
        );

    \I__4908\ : InMux
    port map (
            O => \N__21129\,
            I => \N__21100\
        );

    \I__4907\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21095\
        );

    \I__4906\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21095\
        );

    \I__4905\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21092\
        );

    \I__4904\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21087\
        );

    \I__4903\ : InMux
    port map (
            O => \N__21124\,
            I => \N__21087\
        );

    \I__4902\ : InMux
    port map (
            O => \N__21123\,
            I => \N__21084\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__21118\,
            I => \N__21081\
        );

    \I__4900\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21074\
        );

    \I__4899\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21074\
        );

    \I__4898\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21074\
        );

    \I__4897\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21068\
        );

    \I__4896\ : InMux
    port map (
            O => \N__21111\,
            I => \N__21056\
        );

    \I__4895\ : InMux
    port map (
            O => \N__21110\,
            I => \N__21051\
        );

    \I__4894\ : InMux
    port map (
            O => \N__21109\,
            I => \N__21051\
        );

    \I__4893\ : InMux
    port map (
            O => \N__21108\,
            I => \N__21048\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__21105\,
            I => \N__21043\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__21100\,
            I => \N__21043\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__21095\,
            I => \N__21036\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__21092\,
            I => \N__21036\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__21087\,
            I => \N__21036\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__21084\,
            I => \N__21033\
        );

    \I__4886\ : Span4Mux_v
    port map (
            O => \N__21081\,
            I => \N__21028\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__21074\,
            I => \N__21028\
        );

    \I__4884\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21023\
        );

    \I__4883\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21023\
        );

    \I__4882\ : InMux
    port map (
            O => \N__21071\,
            I => \N__21020\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__21068\,
            I => \N__21017\
        );

    \I__4880\ : InMux
    port map (
            O => \N__21067\,
            I => \N__21010\
        );

    \I__4879\ : InMux
    port map (
            O => \N__21066\,
            I => \N__21010\
        );

    \I__4878\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21010\
        );

    \I__4877\ : InMux
    port map (
            O => \N__21064\,
            I => \N__21007\
        );

    \I__4876\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21002\
        );

    \I__4875\ : InMux
    port map (
            O => \N__21062\,
            I => \N__21002\
        );

    \I__4874\ : InMux
    port map (
            O => \N__21061\,
            I => \N__20995\
        );

    \I__4873\ : InMux
    port map (
            O => \N__21060\,
            I => \N__20995\
        );

    \I__4872\ : InMux
    port map (
            O => \N__21059\,
            I => \N__20995\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__21056\,
            I => \N__20988\
        );

    \I__4870\ : LocalMux
    port map (
            O => \N__21051\,
            I => \N__20988\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__21048\,
            I => \N__20988\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__21043\,
            I => \N__20983\
        );

    \I__4867\ : Span4Mux_v
    port map (
            O => \N__21036\,
            I => \N__20983\
        );

    \I__4866\ : Span4Mux_v
    port map (
            O => \N__21033\,
            I => \N__20980\
        );

    \I__4865\ : Span4Mux_s3_h
    port map (
            O => \N__21028\,
            I => \N__20977\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__21023\,
            I => \Lab_UT.state_0\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__21020\,
            I => \Lab_UT.state_0\
        );

    \I__4862\ : Odrv12
    port map (
            O => \N__21017\,
            I => \Lab_UT.state_0\
        );

    \I__4861\ : LocalMux
    port map (
            O => \N__21010\,
            I => \Lab_UT.state_0\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__21007\,
            I => \Lab_UT.state_0\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__21002\,
            I => \Lab_UT.state_0\
        );

    \I__4858\ : LocalMux
    port map (
            O => \N__20995\,
            I => \Lab_UT.state_0\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__20988\,
            I => \Lab_UT.state_0\
        );

    \I__4856\ : Odrv4
    port map (
            O => \N__20983\,
            I => \Lab_UT.state_0\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__20980\,
            I => \Lab_UT.state_0\
        );

    \I__4854\ : Odrv4
    port map (
            O => \N__20977\,
            I => \Lab_UT.state_0\
        );

    \I__4853\ : InMux
    port map (
            O => \N__20954\,
            I => \N__20944\
        );

    \I__4852\ : InMux
    port map (
            O => \N__20953\,
            I => \N__20944\
        );

    \I__4851\ : InMux
    port map (
            O => \N__20952\,
            I => \N__20936\
        );

    \I__4850\ : InMux
    port map (
            O => \N__20951\,
            I => \N__20936\
        );

    \I__4849\ : InMux
    port map (
            O => \N__20950\,
            I => \N__20936\
        );

    \I__4848\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20933\
        );

    \I__4847\ : LocalMux
    port map (
            O => \N__20944\,
            I => \N__20930\
        );

    \I__4846\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20927\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__20936\,
            I => \N__20924\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__20933\,
            I => \N__20921\
        );

    \I__4843\ : Span4Mux_s2_h
    port map (
            O => \N__20930\,
            I => \N__20918\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__20927\,
            I => \Lab_UT.dictrl.next_stateZ0Z32\
        );

    \I__4841\ : Odrv12
    port map (
            O => \N__20924\,
            I => \Lab_UT.dictrl.next_stateZ0Z32\
        );

    \I__4840\ : Odrv4
    port map (
            O => \N__20921\,
            I => \Lab_UT.dictrl.next_stateZ0Z32\
        );

    \I__4839\ : Odrv4
    port map (
            O => \N__20918\,
            I => \Lab_UT.dictrl.next_stateZ0Z32\
        );

    \I__4838\ : InMux
    port map (
            O => \N__20909\,
            I => \N__20906\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__20906\,
            I => \Lab_UT.dictrl.N_29_0\
        );

    \I__4836\ : CascadeMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__4835\ : InMux
    port map (
            O => \N__20900\,
            I => \N__20896\
        );

    \I__4834\ : CascadeMux
    port map (
            O => \N__20899\,
            I => \N__20893\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__20896\,
            I => \N__20890\
        );

    \I__4832\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20887\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__20890\,
            I => \N__20882\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__20887\,
            I => \N__20882\
        );

    \I__4829\ : Span4Mux_s2_h
    port map (
            O => \N__20882\,
            I => \N__20879\
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__20879\,
            I => bu_rx_data_fast_0
        );

    \I__4827\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20873\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__20873\,
            I => \N__20870\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__20870\,
            I => \Lab_UT.dictrl.g0_0_0_a3_1\
        );

    \I__4824\ : CascadeMux
    port map (
            O => \N__20867\,
            I => \N__20862\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__20866\,
            I => \N__20859\
        );

    \I__4822\ : InMux
    port map (
            O => \N__20865\,
            I => \N__20833\
        );

    \I__4821\ : InMux
    port map (
            O => \N__20862\,
            I => \N__20833\
        );

    \I__4820\ : InMux
    port map (
            O => \N__20859\,
            I => \N__20833\
        );

    \I__4819\ : InMux
    port map (
            O => \N__20858\,
            I => \N__20833\
        );

    \I__4818\ : InMux
    port map (
            O => \N__20857\,
            I => \N__20833\
        );

    \I__4817\ : InMux
    port map (
            O => \N__20856\,
            I => \N__20833\
        );

    \I__4816\ : InMux
    port map (
            O => \N__20855\,
            I => \N__20833\
        );

    \I__4815\ : CascadeMux
    port map (
            O => \N__20854\,
            I => \N__20830\
        );

    \I__4814\ : InMux
    port map (
            O => \N__20853\,
            I => \N__20825\
        );

    \I__4813\ : InMux
    port map (
            O => \N__20852\,
            I => \N__20818\
        );

    \I__4812\ : InMux
    port map (
            O => \N__20851\,
            I => \N__20818\
        );

    \I__4811\ : InMux
    port map (
            O => \N__20850\,
            I => \N__20818\
        );

    \I__4810\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20812\
        );

    \I__4809\ : InMux
    port map (
            O => \N__20848\,
            I => \N__20812\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20808\
        );

    \I__4807\ : InMux
    port map (
            O => \N__20830\,
            I => \N__20801\
        );

    \I__4806\ : InMux
    port map (
            O => \N__20829\,
            I => \N__20801\
        );

    \I__4805\ : InMux
    port map (
            O => \N__20828\,
            I => \N__20801\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__20825\,
            I => \N__20790\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__20818\,
            I => \N__20790\
        );

    \I__4802\ : InMux
    port map (
            O => \N__20817\,
            I => \N__20787\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__20812\,
            I => \N__20784\
        );

    \I__4800\ : InMux
    port map (
            O => \N__20811\,
            I => \N__20781\
        );

    \I__4799\ : Span4Mux_v
    port map (
            O => \N__20808\,
            I => \N__20778\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20801\,
            I => \N__20775\
        );

    \I__4797\ : InMux
    port map (
            O => \N__20800\,
            I => \N__20764\
        );

    \I__4796\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20764\
        );

    \I__4795\ : InMux
    port map (
            O => \N__20798\,
            I => \N__20764\
        );

    \I__4794\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20764\
        );

    \I__4793\ : InMux
    port map (
            O => \N__20796\,
            I => \N__20764\
        );

    \I__4792\ : InMux
    port map (
            O => \N__20795\,
            I => \N__20761\
        );

    \I__4791\ : Span4Mux_h
    port map (
            O => \N__20790\,
            I => \N__20756\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20787\,
            I => \N__20756\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__20784\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__20781\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4787\ : Odrv4
    port map (
            O => \N__20778\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4786\ : Odrv4
    port map (
            O => \N__20775\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__20764\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__20761\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__20756\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20741\,
            I => \N__20738\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__20738\,
            I => \N__20735\
        );

    \I__4780\ : Odrv12
    port map (
            O => \N__20735\,
            I => \Lab_UT.dictrl.g0_0_i_a3_1\
        );

    \I__4779\ : InMux
    port map (
            O => \N__20732\,
            I => \N__20729\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20722\
        );

    \I__4777\ : InMux
    port map (
            O => \N__20728\,
            I => \N__20719\
        );

    \I__4776\ : InMux
    port map (
            O => \N__20727\,
            I => \N__20716\
        );

    \I__4775\ : InMux
    port map (
            O => \N__20726\,
            I => \N__20711\
        );

    \I__4774\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20711\
        );

    \I__4773\ : Span4Mux_v
    port map (
            O => \N__20722\,
            I => \N__20708\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__20719\,
            I => \N__20705\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20716\,
            I => \N__20698\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20711\,
            I => \N__20698\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__20708\,
            I => \N__20698\
        );

    \I__4768\ : Span12Mux_s8_v
    port map (
            O => \N__20705\,
            I => \N__20695\
        );

    \I__4767\ : Odrv4
    port map (
            O => \N__20698\,
            I => \Lab_UT.dicLdAStens_0\
        );

    \I__4766\ : Odrv12
    port map (
            O => \N__20695\,
            I => \Lab_UT.dicLdAStens_0\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__20690\,
            I => \N__20686\
        );

    \I__4764\ : CascadeMux
    port map (
            O => \N__20689\,
            I => \N__20683\
        );

    \I__4763\ : InMux
    port map (
            O => \N__20686\,
            I => \N__20672\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20672\
        );

    \I__4761\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20672\
        );

    \I__4760\ : InMux
    port map (
            O => \N__20681\,
            I => \N__20672\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20672\,
            I => \N__20669\
        );

    \I__4758\ : Odrv4
    port map (
            O => \N__20669\,
            I => \Lab_UT.dictrl.N_40_mux\
        );

    \I__4757\ : CascadeMux
    port map (
            O => \N__20666\,
            I => \N__20659\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__20665\,
            I => \N__20651\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__20664\,
            I => \N__20646\
        );

    \I__4754\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20642\
        );

    \I__4753\ : CascadeMux
    port map (
            O => \N__20662\,
            I => \N__20639\
        );

    \I__4752\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20628\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20658\,
            I => \N__20628\
        );

    \I__4750\ : InMux
    port map (
            O => \N__20657\,
            I => \N__20628\
        );

    \I__4749\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20628\
        );

    \I__4748\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20628\
        );

    \I__4747\ : InMux
    port map (
            O => \N__20654\,
            I => \N__20623\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20651\,
            I => \N__20623\
        );

    \I__4745\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20620\
        );

    \I__4744\ : InMux
    port map (
            O => \N__20649\,
            I => \N__20615\
        );

    \I__4743\ : InMux
    port map (
            O => \N__20646\,
            I => \N__20615\
        );

    \I__4742\ : InMux
    port map (
            O => \N__20645\,
            I => \N__20612\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__20642\,
            I => \N__20609\
        );

    \I__4740\ : InMux
    port map (
            O => \N__20639\,
            I => \N__20598\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__20628\,
            I => \N__20591\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__20623\,
            I => \N__20591\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__20620\,
            I => \N__20591\
        );

    \I__4736\ : LocalMux
    port map (
            O => \N__20615\,
            I => \N__20586\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__20612\,
            I => \N__20586\
        );

    \I__4734\ : Span4Mux_h
    port map (
            O => \N__20609\,
            I => \N__20583\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20608\,
            I => \N__20578\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20607\,
            I => \N__20578\
        );

    \I__4731\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20573\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20573\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20604\,
            I => \N__20570\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20603\,
            I => \N__20563\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20602\,
            I => \N__20563\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20601\,
            I => \N__20563\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__20598\,
            I => \N__20560\
        );

    \I__4724\ : Span12Mux_s10_h
    port map (
            O => \N__20591\,
            I => \N__20557\
        );

    \I__4723\ : Span4Mux_v
    port map (
            O => \N__20586\,
            I => \N__20548\
        );

    \I__4722\ : Span4Mux_v
    port map (
            O => \N__20583\,
            I => \N__20548\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20578\,
            I => \N__20548\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20573\,
            I => \N__20548\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__20570\,
            I => \Lab_UT.state_3\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__20563\,
            I => \Lab_UT.state_3\
        );

    \I__4717\ : Odrv12
    port map (
            O => \N__20560\,
            I => \Lab_UT.state_3\
        );

    \I__4716\ : Odrv12
    port map (
            O => \N__20557\,
            I => \Lab_UT.state_3\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__20548\,
            I => \Lab_UT.state_3\
        );

    \I__4714\ : CascadeMux
    port map (
            O => \N__20537\,
            I => \Lab_UT.dictrl.N_13_cascade_\
        );

    \I__4713\ : CascadeMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20531\,
            I => \N__20528\
        );

    \I__4711\ : LocalMux
    port map (
            O => \N__20528\,
            I => \N__20525\
        );

    \I__4710\ : Span4Mux_h
    port map (
            O => \N__20525\,
            I => \N__20522\
        );

    \I__4709\ : Odrv4
    port map (
            O => \N__20522\,
            I => \Lab_UT.dictrl.N_16\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20516\
        );

    \I__4707\ : LocalMux
    port map (
            O => \N__20516\,
            I => \N__20513\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__20513\,
            I => \N__20509\
        );

    \I__4705\ : InMux
    port map (
            O => \N__20512\,
            I => \N__20506\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__20509\,
            I => \N__20501\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20506\,
            I => \N__20501\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__20501\,
            I => \Lab_UT.dictrl.state_fast_3\
        );

    \I__4701\ : CascadeMux
    port map (
            O => \N__20498\,
            I => \N__20495\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20495\,
            I => \N__20486\
        );

    \I__4699\ : InMux
    port map (
            O => \N__20494\,
            I => \N__20486\
        );

    \I__4698\ : CascadeMux
    port map (
            O => \N__20493\,
            I => \N__20483\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20492\,
            I => \N__20478\
        );

    \I__4696\ : InMux
    port map (
            O => \N__20491\,
            I => \N__20475\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__20486\,
            I => \N__20472\
        );

    \I__4694\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20469\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20464\
        );

    \I__4692\ : InMux
    port map (
            O => \N__20481\,
            I => \N__20464\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20478\,
            I => \N__20457\
        );

    \I__4690\ : LocalMux
    port map (
            O => \N__20475\,
            I => \N__20454\
        );

    \I__4689\ : Span4Mux_h
    port map (
            O => \N__20472\,
            I => \N__20451\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__20469\,
            I => \N__20446\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__20464\,
            I => \N__20446\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20441\
        );

    \I__4685\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20441\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20436\
        );

    \I__4683\ : InMux
    port map (
            O => \N__20460\,
            I => \N__20436\
        );

    \I__4682\ : Span4Mux_s2_h
    port map (
            O => \N__20457\,
            I => \N__20433\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__20454\,
            I => bu_rx_data_2_rep2
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__20451\,
            I => bu_rx_data_2_rep2
        );

    \I__4679\ : Odrv4
    port map (
            O => \N__20446\,
            I => bu_rx_data_2_rep2
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20441\,
            I => bu_rx_data_2_rep2
        );

    \I__4677\ : LocalMux
    port map (
            O => \N__20436\,
            I => bu_rx_data_2_rep2
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__20433\,
            I => bu_rx_data_2_rep2
        );

    \I__4675\ : InMux
    port map (
            O => \N__20420\,
            I => \N__20417\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__20417\,
            I => \Lab_UT.dictrl.N_15\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20414\,
            I => \N__20411\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20411\,
            I => \N__20405\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20410\,
            I => \N__20402\
        );

    \I__4670\ : InMux
    port map (
            O => \N__20409\,
            I => \N__20399\
        );

    \I__4669\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20396\
        );

    \I__4668\ : Span4Mux_v
    port map (
            O => \N__20405\,
            I => \N__20391\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20402\,
            I => \N__20384\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__20399\,
            I => \N__20384\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__20396\,
            I => \N__20384\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20381\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20378\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__20391\,
            I => \N__20373\
        );

    \I__4661\ : Span4Mux_s3_h
    port map (
            O => \N__20384\,
            I => \N__20373\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20381\,
            I => \N__20368\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20378\,
            I => \N__20368\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__20373\,
            I => \Lab_UT.dictrl.next_state12\
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__20368\,
            I => \Lab_UT.dictrl.next_state12\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20363\,
            I => \N__20360\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__20360\,
            I => \N__20357\
        );

    \I__4654\ : Odrv4
    port map (
            O => \N__20357\,
            I => \Lab_UT.bcd2segment4.segment_0Z0Z_0\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20354\,
            I => \N__20351\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20351\,
            I => \N__20348\
        );

    \I__4651\ : Odrv4
    port map (
            O => \N__20348\,
            I => \Lab_UT.bcd2segment4.segment_0Z0Z_1\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__20345\,
            I => \N__20335\
        );

    \I__4649\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20320\
        );

    \I__4648\ : InMux
    port map (
            O => \N__20343\,
            I => \N__20320\
        );

    \I__4647\ : InMux
    port map (
            O => \N__20342\,
            I => \N__20320\
        );

    \I__4646\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20320\
        );

    \I__4645\ : InMux
    port map (
            O => \N__20340\,
            I => \N__20320\
        );

    \I__4644\ : InMux
    port map (
            O => \N__20339\,
            I => \N__20320\
        );

    \I__4643\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20320\
        );

    \I__4642\ : InMux
    port map (
            O => \N__20335\,
            I => \N__20317\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__20320\,
            I => \N__20313\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20307\
        );

    \I__4639\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20304\
        );

    \I__4638\ : Span4Mux_s3_h
    port map (
            O => \N__20313\,
            I => \N__20301\
        );

    \I__4637\ : InMux
    port map (
            O => \N__20312\,
            I => \N__20298\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20311\,
            I => \N__20293\
        );

    \I__4635\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20293\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__20307\,
            I => \N__20290\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20304\,
            I => \N__20285\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__20301\,
            I => \N__20285\
        );

    \I__4631\ : LocalMux
    port map (
            O => \N__20298\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__20293\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__20290\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__20285\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__20276\,
            I => \N__20269\
        );

    \I__4626\ : CascadeMux
    port map (
            O => \N__20275\,
            I => \N__20265\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__20274\,
            I => \N__20261\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20273\,
            I => \N__20246\
        );

    \I__4623\ : InMux
    port map (
            O => \N__20272\,
            I => \N__20246\
        );

    \I__4622\ : InMux
    port map (
            O => \N__20269\,
            I => \N__20246\
        );

    \I__4621\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20246\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20265\,
            I => \N__20246\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20246\
        );

    \I__4618\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20246\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20246\,
            I => \N__20243\
        );

    \I__4616\ : Span4Mux_s1_h
    port map (
            O => \N__20243\,
            I => \N__20237\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20234\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20229\
        );

    \I__4613\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20229\
        );

    \I__4612\ : Span4Mux_h
    port map (
            O => \N__20237\,
            I => \N__20226\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__20234\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__20229\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__4609\ : Odrv4
    port map (
            O => \N__20226\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__20219\,
            I => \N__20210\
        );

    \I__4607\ : CascadeMux
    port map (
            O => \N__20218\,
            I => \N__20207\
        );

    \I__4606\ : CascadeMux
    port map (
            O => \N__20217\,
            I => \N__20204\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__20216\,
            I => \N__20201\
        );

    \I__4604\ : InMux
    port map (
            O => \N__20215\,
            I => \N__20194\
        );

    \I__4603\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20194\
        );

    \I__4602\ : InMux
    port map (
            O => \N__20213\,
            I => \N__20194\
        );

    \I__4601\ : InMux
    port map (
            O => \N__20210\,
            I => \N__20185\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20185\
        );

    \I__4599\ : InMux
    port map (
            O => \N__20204\,
            I => \N__20185\
        );

    \I__4598\ : InMux
    port map (
            O => \N__20201\,
            I => \N__20185\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20194\,
            I => \N__20179\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__20185\,
            I => \N__20179\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__20184\,
            I => \N__20174\
        );

    \I__4594\ : Span4Mux_s1_h
    port map (
            O => \N__20179\,
            I => \N__20169\
        );

    \I__4593\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20162\
        );

    \I__4592\ : InMux
    port map (
            O => \N__20177\,
            I => \N__20162\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20174\,
            I => \N__20162\
        );

    \I__4590\ : InMux
    port map (
            O => \N__20173\,
            I => \N__20157\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20172\,
            I => \N__20157\
        );

    \I__4588\ : Span4Mux_h
    port map (
            O => \N__20169\,
            I => \N__20154\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__20162\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__20157\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__4585\ : Odrv4
    port map (
            O => \N__20154\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__4584\ : InMux
    port map (
            O => \N__20147\,
            I => \N__20131\
        );

    \I__4583\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20131\
        );

    \I__4582\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20131\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20131\
        );

    \I__4580\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20124\
        );

    \I__4579\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20124\
        );

    \I__4578\ : InMux
    port map (
            O => \N__20141\,
            I => \N__20124\
        );

    \I__4577\ : CascadeMux
    port map (
            O => \N__20140\,
            I => \N__20120\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__20131\,
            I => \N__20115\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__20124\,
            I => \N__20115\
        );

    \I__4574\ : CascadeMux
    port map (
            O => \N__20123\,
            I => \N__20112\
        );

    \I__4573\ : InMux
    port map (
            O => \N__20120\,
            I => \N__20104\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__20115\,
            I => \N__20101\
        );

    \I__4571\ : InMux
    port map (
            O => \N__20112\,
            I => \N__20098\
        );

    \I__4570\ : InMux
    port map (
            O => \N__20111\,
            I => \N__20093\
        );

    \I__4569\ : InMux
    port map (
            O => \N__20110\,
            I => \N__20093\
        );

    \I__4568\ : InMux
    port map (
            O => \N__20109\,
            I => \N__20086\
        );

    \I__4567\ : InMux
    port map (
            O => \N__20108\,
            I => \N__20086\
        );

    \I__4566\ : InMux
    port map (
            O => \N__20107\,
            I => \N__20086\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__20104\,
            I => \N__20083\
        );

    \I__4564\ : Span4Mux_v
    port map (
            O => \N__20101\,
            I => \N__20080\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__20098\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__20093\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__20086\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4560\ : Odrv12
    port map (
            O => \N__20083\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4559\ : Odrv4
    port map (
            O => \N__20080\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4558\ : CascadeMux
    port map (
            O => \N__20069\,
            I => \Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_\
        );

    \I__4557\ : InMux
    port map (
            O => \N__20066\,
            I => \N__20060\
        );

    \I__4556\ : InMux
    port map (
            O => \N__20065\,
            I => \N__20060\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__20060\,
            I => \N__20049\
        );

    \I__4554\ : InMux
    port map (
            O => \N__20059\,
            I => \N__20046\
        );

    \I__4553\ : InMux
    port map (
            O => \N__20058\,
            I => \N__20043\
        );

    \I__4552\ : InMux
    port map (
            O => \N__20057\,
            I => \N__20034\
        );

    \I__4551\ : InMux
    port map (
            O => \N__20056\,
            I => \N__20034\
        );

    \I__4550\ : InMux
    port map (
            O => \N__20055\,
            I => \N__20034\
        );

    \I__4549\ : InMux
    port map (
            O => \N__20054\,
            I => \N__20034\
        );

    \I__4548\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20025\
        );

    \I__4547\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20025\
        );

    \I__4546\ : Span4Mux_v
    port map (
            O => \N__20049\,
            I => \N__20014\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__20014\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__20043\,
            I => \N__20011\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__20034\,
            I => \N__20008\
        );

    \I__4542\ : InMux
    port map (
            O => \N__20033\,
            I => \N__19999\
        );

    \I__4541\ : InMux
    port map (
            O => \N__20032\,
            I => \N__19999\
        );

    \I__4540\ : InMux
    port map (
            O => \N__20031\,
            I => \N__19999\
        );

    \I__4539\ : InMux
    port map (
            O => \N__20030\,
            I => \N__19999\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__20025\,
            I => \N__19996\
        );

    \I__4537\ : InMux
    port map (
            O => \N__20024\,
            I => \N__19989\
        );

    \I__4536\ : InMux
    port map (
            O => \N__20023\,
            I => \N__19989\
        );

    \I__4535\ : InMux
    port map (
            O => \N__20022\,
            I => \N__19989\
        );

    \I__4534\ : InMux
    port map (
            O => \N__20021\,
            I => \N__19982\
        );

    \I__4533\ : InMux
    port map (
            O => \N__20020\,
            I => \N__19982\
        );

    \I__4532\ : InMux
    port map (
            O => \N__20019\,
            I => \N__19982\
        );

    \I__4531\ : Span4Mux_v
    port map (
            O => \N__20014\,
            I => \N__19971\
        );

    \I__4530\ : Span4Mux_v
    port map (
            O => \N__20011\,
            I => \N__19968\
        );

    \I__4529\ : Span4Mux_v
    port map (
            O => \N__20008\,
            I => \N__19963\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__19999\,
            I => \N__19963\
        );

    \I__4527\ : Span4Mux_v
    port map (
            O => \N__19996\,
            I => \N__19956\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__19989\,
            I => \N__19956\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19956\
        );

    \I__4524\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19953\
        );

    \I__4523\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19950\
        );

    \I__4522\ : InMux
    port map (
            O => \N__19979\,
            I => \N__19937\
        );

    \I__4521\ : InMux
    port map (
            O => \N__19978\,
            I => \N__19937\
        );

    \I__4520\ : InMux
    port map (
            O => \N__19977\,
            I => \N__19937\
        );

    \I__4519\ : InMux
    port map (
            O => \N__19976\,
            I => \N__19937\
        );

    \I__4518\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19937\
        );

    \I__4517\ : InMux
    port map (
            O => \N__19974\,
            I => \N__19937\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__19971\,
            I => \Lab_UT.Run\
        );

    \I__4515\ : Odrv4
    port map (
            O => \N__19968\,
            I => \Lab_UT.Run\
        );

    \I__4514\ : Odrv4
    port map (
            O => \N__19963\,
            I => \Lab_UT.Run\
        );

    \I__4513\ : Odrv4
    port map (
            O => \N__19956\,
            I => \Lab_UT.Run\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__19953\,
            I => \Lab_UT.Run\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__19950\,
            I => \Lab_UT.Run\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__19937\,
            I => \Lab_UT.Run\
        );

    \I__4509\ : InMux
    port map (
            O => \N__19922\,
            I => \N__19919\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19916\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__19916\,
            I => \N__19913\
        );

    \I__4506\ : Odrv4
    port map (
            O => \N__19913\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__4505\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19898\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19909\,
            I => \N__19898\
        );

    \I__4503\ : InMux
    port map (
            O => \N__19908\,
            I => \N__19898\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19898\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19898\,
            I => \N__19895\
        );

    \I__4500\ : Odrv4
    port map (
            O => \N__19895\,
            I => \Lab_UT.dictrl.N_39_mux\
        );

    \I__4499\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19889\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__19889\,
            I => \N__19886\
        );

    \I__4497\ : Span4Mux_h
    port map (
            O => \N__19886\,
            I => \N__19883\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__19883\,
            I => \Lab_UT.dictrl.g0_0_a3_2\
        );

    \I__4495\ : InMux
    port map (
            O => \N__19880\,
            I => \N__19867\
        );

    \I__4494\ : CascadeMux
    port map (
            O => \N__19879\,
            I => \N__19864\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__19878\,
            I => \N__19860\
        );

    \I__4492\ : InMux
    port map (
            O => \N__19877\,
            I => \N__19857\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19876\,
            I => \N__19852\
        );

    \I__4490\ : InMux
    port map (
            O => \N__19875\,
            I => \N__19849\
        );

    \I__4489\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19846\
        );

    \I__4488\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19843\
        );

    \I__4487\ : InMux
    port map (
            O => \N__19872\,
            I => \N__19840\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__19871\,
            I => \N__19837\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__19870\,
            I => \N__19834\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19829\
        );

    \I__4483\ : InMux
    port map (
            O => \N__19864\,
            I => \N__19826\
        );

    \I__4482\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19821\
        );

    \I__4481\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19821\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19818\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19856\,
            I => \N__19815\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__19855\,
            I => \N__19812\
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19805\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19849\,
            I => \N__19805\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__19846\,
            I => \N__19805\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__19843\,
            I => \N__19800\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19800\
        );

    \I__4472\ : InMux
    port map (
            O => \N__19837\,
            I => \N__19797\
        );

    \I__4471\ : InMux
    port map (
            O => \N__19834\,
            I => \N__19792\
        );

    \I__4470\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19792\
        );

    \I__4469\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19789\
        );

    \I__4468\ : Span4Mux_v
    port map (
            O => \N__19829\,
            I => \N__19784\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__19826\,
            I => \N__19784\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19821\,
            I => \N__19781\
        );

    \I__4465\ : Span4Mux_v
    port map (
            O => \N__19818\,
            I => \N__19775\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__19815\,
            I => \N__19772\
        );

    \I__4463\ : InMux
    port map (
            O => \N__19812\,
            I => \N__19769\
        );

    \I__4462\ : Span4Mux_v
    port map (
            O => \N__19805\,
            I => \N__19766\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__19800\,
            I => \N__19759\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__19797\,
            I => \N__19759\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__19792\,
            I => \N__19759\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__19789\,
            I => \N__19756\
        );

    \I__4457\ : Span4Mux_h
    port map (
            O => \N__19784\,
            I => \N__19753\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__19781\,
            I => \N__19750\
        );

    \I__4455\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19747\
        );

    \I__4454\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19742\
        );

    \I__4453\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19742\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__19775\,
            I => \N__19735\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__19772\,
            I => \N__19735\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__19769\,
            I => \N__19735\
        );

    \I__4449\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19730\
        );

    \I__4448\ : Span4Mux_v
    port map (
            O => \N__19759\,
            I => \N__19730\
        );

    \I__4447\ : Span4Mux_s2_v
    port map (
            O => \N__19756\,
            I => \N__19723\
        );

    \I__4446\ : Span4Mux_v
    port map (
            O => \N__19753\,
            I => \N__19723\
        );

    \I__4445\ : Span4Mux_h
    port map (
            O => \N__19750\,
            I => \N__19723\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__19747\,
            I => bu_rx_data_2
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__19742\,
            I => bu_rx_data_2
        );

    \I__4442\ : Odrv4
    port map (
            O => \N__19735\,
            I => bu_rx_data_2
        );

    \I__4441\ : Odrv4
    port map (
            O => \N__19730\,
            I => bu_rx_data_2
        );

    \I__4440\ : Odrv4
    port map (
            O => \N__19723\,
            I => bu_rx_data_2
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__19712\,
            I => \N__19709\
        );

    \I__4438\ : InMux
    port map (
            O => \N__19709\,
            I => \N__19700\
        );

    \I__4437\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19700\
        );

    \I__4436\ : InMux
    port map (
            O => \N__19707\,
            I => \N__19700\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__19700\,
            I => \N__19695\
        );

    \I__4434\ : CascadeMux
    port map (
            O => \N__19699\,
            I => \N__19691\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__19698\,
            I => \N__19688\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__19695\,
            I => \N__19685\
        );

    \I__4431\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19678\
        );

    \I__4430\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19678\
        );

    \I__4429\ : InMux
    port map (
            O => \N__19688\,
            I => \N__19678\
        );

    \I__4428\ : Odrv4
    port map (
            O => \N__19685\,
            I => bu_rx_data_3_rep1
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__19678\,
            I => bu_rx_data_3_rep1
        );

    \I__4426\ : InMux
    port map (
            O => \N__19673\,
            I => \N__19670\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19670\,
            I => \N__19667\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__19667\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__4423\ : InMux
    port map (
            O => \N__19664\,
            I => \N__19661\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19661\,
            I => \N__19658\
        );

    \I__4421\ : Odrv4
    port map (
            O => \N__19658\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__4420\ : InMux
    port map (
            O => \N__19655\,
            I => \N__19652\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19649\
        );

    \I__4418\ : Odrv4
    port map (
            O => \N__19649\,
            I => \Lab_UT.bcd2segment4.segment_0Z0Z_2\
        );

    \I__4417\ : InMux
    port map (
            O => \N__19646\,
            I => \N__19643\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19640\
        );

    \I__4415\ : Odrv4
    port map (
            O => \N__19640\,
            I => \Lab_UT.bcd2segment4.segmentUQ_0_4\
        );

    \I__4414\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19634\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__19634\,
            I => \N__19631\
        );

    \I__4412\ : Odrv4
    port map (
            O => \N__19631\,
            I => \Lab_UT.bcd2segment4.segmentUQ_0_5\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19628\,
            I => \N__19625\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19625\,
            I => \N__19622\
        );

    \I__4409\ : Odrv4
    port map (
            O => \N__19622\,
            I => \Lab_UT.bcd2segment4.segmentUQ_0_6\
        );

    \I__4408\ : InMux
    port map (
            O => \N__19619\,
            I => \N__19616\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19616\,
            I => \Lab_UT.dictrl.g1_2_3\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19610\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__19610\,
            I => \Lab_UT.dictrl.g0_1Z0Z_1\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19604\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19604\,
            I => \Lab_UT.dictrl.g0_i_a3_4\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19601\,
            I => \N__19596\
        );

    \I__4401\ : CascadeMux
    port map (
            O => \N__19600\,
            I => \N__19589\
        );

    \I__4400\ : CascadeMux
    port map (
            O => \N__19599\,
            I => \N__19585\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19596\,
            I => \N__19582\
        );

    \I__4398\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19577\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19594\,
            I => \N__19577\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19593\,
            I => \N__19572\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19592\,
            I => \N__19572\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19589\,
            I => \N__19565\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19565\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19585\,
            I => \N__19565\
        );

    \I__4391\ : Odrv4
    port map (
            O => \N__19582\,
            I => bu_rx_data_4_rep1
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__19577\,
            I => bu_rx_data_4_rep1
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19572\,
            I => bu_rx_data_4_rep1
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19565\,
            I => bu_rx_data_4_rep1
        );

    \I__4387\ : InMux
    port map (
            O => \N__19556\,
            I => \N__19553\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19549\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19546\
        );

    \I__4384\ : Span4Mux_h
    port map (
            O => \N__19549\,
            I => \N__19537\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__19546\,
            I => \N__19534\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19527\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19527\
        );

    \I__4380\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19527\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19542\,
            I => \N__19520\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19520\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19540\,
            I => \N__19520\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__19537\,
            I => bu_rx_data_7_rep1
        );

    \I__4375\ : Odrv12
    port map (
            O => \N__19534\,
            I => bu_rx_data_7_rep1
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__19527\,
            I => bu_rx_data_7_rep1
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19520\,
            I => bu_rx_data_7_rep1
        );

    \I__4372\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19508\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19508\,
            I => \Lab_UT.dictrl.g1_4_0\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__19505\,
            I => \N__19500\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19496\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19503\,
            I => \N__19493\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19490\
        );

    \I__4366\ : CascadeMux
    port map (
            O => \N__19499\,
            I => \N__19487\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19481\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19493\,
            I => \N__19481\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19490\,
            I => \N__19478\
        );

    \I__4362\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19475\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19486\,
            I => \N__19472\
        );

    \I__4360\ : Span4Mux_h
    port map (
            O => \N__19481\,
            I => \N__19469\
        );

    \I__4359\ : Odrv4
    port map (
            O => \N__19478\,
            I => bu_rx_data_2_rep1
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19475\,
            I => bu_rx_data_2_rep1
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19472\,
            I => bu_rx_data_2_rep1
        );

    \I__4356\ : Odrv4
    port map (
            O => \N__19469\,
            I => bu_rx_data_2_rep1
        );

    \I__4355\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19457\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__19457\,
            I => \N__19454\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__19454\,
            I => \N__19446\
        );

    \I__4352\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19443\
        );

    \I__4351\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19438\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19438\
        );

    \I__4349\ : InMux
    port map (
            O => \N__19450\,
            I => \N__19433\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19433\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__19446\,
            I => bu_rx_data_fast_2
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19443\,
            I => bu_rx_data_fast_2
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__19438\,
            I => bu_rx_data_fast_2
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__19433\,
            I => bu_rx_data_fast_2
        );

    \I__4343\ : CascadeMux
    port map (
            O => \N__19424\,
            I => \N__19420\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19415\
        );

    \I__4341\ : InMux
    port map (
            O => \N__19420\,
            I => \N__19408\
        );

    \I__4340\ : InMux
    port map (
            O => \N__19419\,
            I => \N__19403\
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__19418\,
            I => \N__19399\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__19415\,
            I => \N__19396\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19393\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__19413\,
            I => \N__19390\
        );

    \I__4335\ : InMux
    port map (
            O => \N__19412\,
            I => \N__19386\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19411\,
            I => \N__19383\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19408\,
            I => \N__19380\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19407\,
            I => \N__19377\
        );

    \I__4331\ : InMux
    port map (
            O => \N__19406\,
            I => \N__19374\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19403\,
            I => \N__19371\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19402\,
            I => \N__19366\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19399\,
            I => \N__19366\
        );

    \I__4327\ : Span4Mux_v
    port map (
            O => \N__19396\,
            I => \N__19359\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19359\
        );

    \I__4325\ : InMux
    port map (
            O => \N__19390\,
            I => \N__19356\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19389\,
            I => \N__19353\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__19386\,
            I => \N__19347\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19383\,
            I => \N__19347\
        );

    \I__4321\ : Span4Mux_v
    port map (
            O => \N__19380\,
            I => \N__19340\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__19377\,
            I => \N__19340\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19374\,
            I => \N__19340\
        );

    \I__4318\ : Span4Mux_h
    port map (
            O => \N__19371\,
            I => \N__19333\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__19366\,
            I => \N__19333\
        );

    \I__4316\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19330\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19327\
        );

    \I__4314\ : Span4Mux_h
    port map (
            O => \N__19359\,
            I => \N__19317\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19356\,
            I => \N__19317\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19353\,
            I => \N__19314\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19352\,
            I => \N__19311\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__19347\,
            I => \N__19306\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__19340\,
            I => \N__19306\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19301\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19301\
        );

    \I__4306\ : Span4Mux_h
    port map (
            O => \N__19333\,
            I => \N__19294\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19294\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__19327\,
            I => \N__19294\
        );

    \I__4303\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19291\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19325\,
            I => \N__19282\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19324\,
            I => \N__19282\
        );

    \I__4300\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19282\
        );

    \I__4299\ : InMux
    port map (
            O => \N__19322\,
            I => \N__19282\
        );

    \I__4298\ : Span4Mux_v
    port map (
            O => \N__19317\,
            I => \N__19279\
        );

    \I__4297\ : Sp12to4
    port map (
            O => \N__19314\,
            I => \N__19270\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19311\,
            I => \N__19270\
        );

    \I__4295\ : Sp12to4
    port map (
            O => \N__19306\,
            I => \N__19270\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__19301\,
            I => \N__19270\
        );

    \I__4293\ : Span4Mux_v
    port map (
            O => \N__19294\,
            I => \N__19265\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19291\,
            I => \N__19265\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__19282\,
            I => bu_rx_data_3
        );

    \I__4290\ : Odrv4
    port map (
            O => \N__19279\,
            I => bu_rx_data_3
        );

    \I__4289\ : Odrv12
    port map (
            O => \N__19270\,
            I => bu_rx_data_3
        );

    \I__4288\ : Odrv4
    port map (
            O => \N__19265\,
            I => bu_rx_data_3
        );

    \I__4287\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19253\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19250\
        );

    \I__4285\ : Span4Mux_h
    port map (
            O => \N__19250\,
            I => \N__19242\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19249\,
            I => \N__19239\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19234\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19247\,
            I => \N__19234\
        );

    \I__4281\ : InMux
    port map (
            O => \N__19246\,
            I => \N__19229\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19229\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__19242\,
            I => bu_rx_data_fast_1
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19239\,
            I => bu_rx_data_fast_1
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__19234\,
            I => bu_rx_data_fast_1
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__19229\,
            I => bu_rx_data_fast_1
        );

    \I__4275\ : CascadeMux
    port map (
            O => \N__19220\,
            I => \Lab_UT.dictrl.g0_i_a3_0_0_cascade_\
        );

    \I__4274\ : CascadeMux
    port map (
            O => \N__19217\,
            I => \Lab_UT.dictrl.g0_i_a3_0_6_cascade_\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19214\,
            I => \N__19211\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19211\,
            I => \Lab_UT.dictrl.g0_i_a3_0_5\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19202\
        );

    \I__4270\ : InMux
    port map (
            O => \N__19207\,
            I => \N__19202\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19197\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19201\,
            I => \N__19194\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19191\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__19197\,
            I => \Lab_UT.dictrl.N_3\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19194\,
            I => \Lab_UT.dictrl.N_3\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__19191\,
            I => \Lab_UT.dictrl.N_3\
        );

    \I__4263\ : InMux
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__19181\,
            I => \Lab_UT.dictrl.g1_4\
        );

    \I__4261\ : CascadeMux
    port map (
            O => \N__19178\,
            I => \N__19172\
        );

    \I__4260\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19167\
        );

    \I__4259\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19167\
        );

    \I__4258\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19164\
        );

    \I__4257\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19161\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__19167\,
            I => \N__19157\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__19164\,
            I => \N__19152\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19161\,
            I => \N__19152\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19160\,
            I => \N__19149\
        );

    \I__4252\ : Odrv4
    port map (
            O => \N__19157\,
            I => \Lab_UT.dictrl.gZ0Z1\
        );

    \I__4251\ : Odrv4
    port map (
            O => \N__19152\,
            I => \Lab_UT.dictrl.gZ0Z1\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__19149\,
            I => \Lab_UT.dictrl.gZ0Z1\
        );

    \I__4249\ : InMux
    port map (
            O => \N__19142\,
            I => \N__19134\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19131\
        );

    \I__4247\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19128\
        );

    \I__4246\ : InMux
    port map (
            O => \N__19139\,
            I => \N__19125\
        );

    \I__4245\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19120\
        );

    \I__4244\ : InMux
    port map (
            O => \N__19137\,
            I => \N__19120\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__19134\,
            I => \N__19115\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__19131\,
            I => \N__19115\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__19128\,
            I => \N__19112\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__19125\,
            I => \N__19109\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19106\
        );

    \I__4238\ : Span4Mux_v
    port map (
            O => \N__19115\,
            I => \N__19103\
        );

    \I__4237\ : Odrv4
    port map (
            O => \N__19112\,
            I => \Lab_UT.dictrl.next_state12_1\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__19109\,
            I => \Lab_UT.dictrl.next_state12_1\
        );

    \I__4235\ : Odrv12
    port map (
            O => \N__19106\,
            I => \Lab_UT.dictrl.next_state12_1\
        );

    \I__4234\ : Odrv4
    port map (
            O => \N__19103\,
            I => \Lab_UT.dictrl.next_state12_1\
        );

    \I__4233\ : InMux
    port map (
            O => \N__19094\,
            I => \N__19089\
        );

    \I__4232\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19086\
        );

    \I__4231\ : InMux
    port map (
            O => \N__19092\,
            I => \N__19083\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__19089\,
            I => \N__19078\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__19086\,
            I => \N__19078\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__19083\,
            I => \N__19075\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__19078\,
            I => \N__19072\
        );

    \I__4226\ : Odrv4
    port map (
            O => \N__19075\,
            I => \Lab_UT.dictrl.next_state32Z0Z_4\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__19072\,
            I => \Lab_UT.dictrl.next_state32Z0Z_4\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__19067\,
            I => \Lab_UT.dictrl.g1Z0Z_0_cascade_\
        );

    \I__4223\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19061\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__19061\,
            I => \Lab_UT.dictrl.N_13_0_0\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__19058\,
            I => \Lab_UT.dictrl.g1_2_2_cascade_\
        );

    \I__4220\ : InMux
    port map (
            O => \N__19055\,
            I => \N__19052\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__19052\,
            I => \Lab_UT.dictrl.g2_1_1\
        );

    \I__4218\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19046\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__19046\,
            I => \Lab_UT.dictrl.g2_0\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4215\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__19037\,
            I => \N__19033\
        );

    \I__4213\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19030\
        );

    \I__4212\ : Odrv4
    port map (
            O => \N__19033\,
            I => \Lab_UT.dictrl.i6_mux\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__19030\,
            I => \Lab_UT.dictrl.i6_mux\
        );

    \I__4210\ : CascadeMux
    port map (
            O => \N__19025\,
            I => \Lab_UT.dictrl.N_15_0_cascade_\
        );

    \I__4209\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19019\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__19014\
        );

    \I__4207\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19006\
        );

    \I__4206\ : InMux
    port map (
            O => \N__19017\,
            I => \N__19006\
        );

    \I__4205\ : Span4Mux_h
    port map (
            O => \N__19014\,
            I => \N__19002\
        );

    \I__4204\ : InMux
    port map (
            O => \N__19013\,
            I => \N__18997\
        );

    \I__4203\ : InMux
    port map (
            O => \N__19012\,
            I => \N__18997\
        );

    \I__4202\ : InMux
    port map (
            O => \N__19011\,
            I => \N__18994\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__19006\,
            I => \N__18991\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19005\,
            I => \N__18988\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__19002\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__18997\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__18994\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__18991\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__18988\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__18977\,
            I => \N__18973\
        );

    \I__4193\ : CascadeMux
    port map (
            O => \N__18976\,
            I => \N__18970\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18973\,
            I => \N__18962\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18962\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18955\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18955\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18967\,
            I => \N__18955\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__18962\,
            I => \N__18952\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18949\
        );

    \I__4185\ : Span4Mux_h
    port map (
            O => \N__18952\,
            I => \N__18946\
        );

    \I__4184\ : Odrv4
    port map (
            O => \N__18949\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_0\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__18946\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_0\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__18941\,
            I => \N__18935\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18940\,
            I => \N__18931\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18939\,
            I => \N__18926\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18938\,
            I => \N__18926\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18921\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18921\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__18931\,
            I => \N__18918\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__18926\,
            I => \N__18915\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__18921\,
            I => \N__18912\
        );

    \I__4173\ : Span4Mux_v
    port map (
            O => \N__18918\,
            I => \N__18905\
        );

    \I__4172\ : Span4Mux_v
    port map (
            O => \N__18915\,
            I => \N__18905\
        );

    \I__4171\ : Span4Mux_h
    port map (
            O => \N__18912\,
            I => \N__18905\
        );

    \I__4170\ : Odrv4
    port map (
            O => \N__18905\,
            I => \Lab_UT.LdMtens\
        );

    \I__4169\ : CascadeMux
    port map (
            O => \N__18902\,
            I => \Lab_UT.dictrl.g0_6_o3_2_0_cascade_\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__18899\,
            I => \Lab_UT.dictrl.N_5_0_cascade_\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18893\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__18893\,
            I => \Lab_UT.dictrl.g1_3_0\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18890\,
            I => \N__18887\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18884\
        );

    \I__4163\ : Span4Mux_h
    port map (
            O => \N__18884\,
            I => \N__18881\
        );

    \I__4162\ : Odrv4
    port map (
            O => \N__18881\,
            I => \Lab_UT.dictrl.g2_2\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18878\,
            I => \N__18872\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18867\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18867\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18864\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18859\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__18867\,
            I => \N__18859\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__18864\,
            I => \N__18856\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__18859\,
            I => \Lab_UT.dictrl.N_16_0_0\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__18856\,
            I => \Lab_UT.dictrl.N_16_0_0\
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__18851\,
            I => \Lab_UT.dictrl.N_19_cascade_\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__18848\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18842\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__18842\,
            I => \Lab_UT.dictrl.N_19\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18835\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18832\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__18835\,
            I => \N__18826\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__18832\,
            I => \N__18826\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18823\
        );

    \I__4143\ : Span4Mux_h
    port map (
            O => \N__18826\,
            I => \N__18820\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18823\,
            I => \Lab_UT.dictrl.N_11_0_0\
        );

    \I__4141\ : Odrv4
    port map (
            O => \N__18820\,
            I => \Lab_UT.dictrl.N_11_0_0\
        );

    \I__4140\ : CascadeMux
    port map (
            O => \N__18815\,
            I => \Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4138\ : LocalMux
    port map (
            O => \N__18809\,
            I => \Lab_UT.dictrl.state_ret_5_RNOZ0Z_1\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18799\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18799\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18796\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__18799\,
            I => \Lab_UT.dicRun_1\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__18796\,
            I => \Lab_UT.dicRun_1\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18788\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18785\
        );

    \I__4130\ : Odrv4
    port map (
            O => \N__18785\,
            I => \Lab_UT.dictrl.N_10\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18779\
        );

    \I__4128\ : LocalMux
    port map (
            O => \N__18779\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_2\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18776\,
            I => \Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18766\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18763\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18760\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18757\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18754\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__18766\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__18763\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4119\ : LocalMux
    port map (
            O => \N__18760\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__18757\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__18754\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18740\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__18740\,
            I => \N__18737\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__18737\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_3\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__18734\,
            I => \Lab_UT.dictrl.N_14_cascade_\
        );

    \I__4112\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18728\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18728\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_3\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__18725\,
            I => \Lab_UT.dictrl.N_7_cascade_\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__18722\,
            I => \Lab_UT.dictrl.N_13_0_cascade_\
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__18719\,
            I => \Lab_UT.dictrl.N_6_cascade_\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__18716\,
            I => \N__18713\
        );

    \I__4106\ : InMux
    port map (
            O => \N__18713\,
            I => \N__18709\
        );

    \I__4105\ : InMux
    port map (
            O => \N__18712\,
            I => \N__18706\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__18709\,
            I => \N__18701\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18698\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__18705\,
            I => \N__18695\
        );

    \I__4101\ : InMux
    port map (
            O => \N__18704\,
            I => \N__18692\
        );

    \I__4100\ : Span4Mux_v
    port map (
            O => \N__18701\,
            I => \N__18687\
        );

    \I__4099\ : Span4Mux_s3_v
    port map (
            O => \N__18698\,
            I => \N__18687\
        );

    \I__4098\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18684\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18681\
        );

    \I__4096\ : Span4Mux_v
    port map (
            O => \N__18687\,
            I => \N__18676\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18684\,
            I => \N__18676\
        );

    \I__4094\ : Odrv12
    port map (
            O => \N__18681\,
            I => \Lab_UT.LdStens\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__18676\,
            I => \Lab_UT.LdStens\
        );

    \I__4092\ : InMux
    port map (
            O => \N__18671\,
            I => \N__18666\
        );

    \I__4091\ : InMux
    port map (
            O => \N__18670\,
            I => \N__18661\
        );

    \I__4090\ : InMux
    port map (
            O => \N__18669\,
            I => \N__18661\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18666\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__18661\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__18656\,
            I => \N__18653\
        );

    \I__4086\ : InMux
    port map (
            O => \N__18653\,
            I => \N__18650\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18650\,
            I => \Lab_UT.LdStens_i_3\
        );

    \I__4084\ : InMux
    port map (
            O => \N__18647\,
            I => \N__18641\
        );

    \I__4083\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18641\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18638\
        );

    \I__4081\ : Span4Mux_v
    port map (
            O => \N__18638\,
            I => \N__18635\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__18635\,
            I => \Lab_UT.didp.ce_10_0_1\
        );

    \I__4079\ : InMux
    port map (
            O => \N__18632\,
            I => \N__18629\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__18629\,
            I => \N__18626\
        );

    \I__4077\ : Span4Mux_v
    port map (
            O => \N__18626\,
            I => \N__18623\
        );

    \I__4076\ : Span4Mux_h
    port map (
            O => \N__18623\,
            I => \N__18620\
        );

    \I__4075\ : Odrv4
    port map (
            O => \N__18620\,
            I => \Lab_UT.dictrl.m27_1\
        );

    \I__4074\ : InMux
    port map (
            O => \N__18617\,
            I => \N__18614\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__18614\,
            I => \N__18611\
        );

    \I__4072\ : Odrv12
    port map (
            O => \N__18611\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_0\
        );

    \I__4071\ : InMux
    port map (
            O => \N__18608\,
            I => \N__18605\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__18605\,
            I => \N__18602\
        );

    \I__4069\ : Odrv4
    port map (
            O => \N__18602\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_3\
        );

    \I__4068\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18596\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__4066\ : Span4Mux_v
    port map (
            O => \N__18593\,
            I => \N__18590\
        );

    \I__4065\ : Odrv4
    port map (
            O => \N__18590\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_2\
        );

    \I__4064\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18584\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__18584\,
            I => \N__18581\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__18581\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_5\
        );

    \I__4061\ : InMux
    port map (
            O => \N__18578\,
            I => \N__18575\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__18575\,
            I => \N__18572\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__18572\,
            I => \N__18569\
        );

    \I__4058\ : Odrv4
    port map (
            O => \N__18569\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_6\
        );

    \I__4057\ : InMux
    port map (
            O => \N__18566\,
            I => \N__18563\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__18563\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_0\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18560\,
            I => \N__18557\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18557\,
            I => \N__18554\
        );

    \I__4053\ : Span4Mux_h
    port map (
            O => \N__18554\,
            I => \N__18551\
        );

    \I__4052\ : Odrv4
    port map (
            O => \N__18551\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_1\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18548\,
            I => \N__18527\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18547\,
            I => \N__18527\
        );

    \I__4049\ : InMux
    port map (
            O => \N__18546\,
            I => \N__18527\
        );

    \I__4048\ : InMux
    port map (
            O => \N__18545\,
            I => \N__18527\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18544\,
            I => \N__18527\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18543\,
            I => \N__18527\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18542\,
            I => \N__18527\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18527\,
            I => \N__18520\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18517\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18512\
        );

    \I__4041\ : InMux
    port map (
            O => \N__18524\,
            I => \N__18512\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18509\
        );

    \I__4039\ : Span4Mux_h
    port map (
            O => \N__18520\,
            I => \N__18506\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18517\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18512\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__18509\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4035\ : Odrv4
    port map (
            O => \N__18506\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4034\ : CascadeMux
    port map (
            O => \N__18497\,
            I => \N__18491\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__18496\,
            I => \N__18488\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__18495\,
            I => \N__18484\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18494\,
            I => \N__18466\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18491\,
            I => \N__18466\
        );

    \I__4029\ : InMux
    port map (
            O => \N__18488\,
            I => \N__18466\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18466\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18484\,
            I => \N__18466\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18483\,
            I => \N__18466\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18466\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18459\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18456\
        );

    \I__4022\ : InMux
    port map (
            O => \N__18465\,
            I => \N__18453\
        );

    \I__4021\ : InMux
    port map (
            O => \N__18464\,
            I => \N__18448\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18463\,
            I => \N__18448\
        );

    \I__4019\ : InMux
    port map (
            O => \N__18462\,
            I => \N__18445\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18459\,
            I => \N__18440\
        );

    \I__4017\ : Span4Mux_v
    port map (
            O => \N__18456\,
            I => \N__18440\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18453\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__18448\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18445\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4013\ : Odrv4
    port map (
            O => \N__18440\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__18431\,
            I => \N__18425\
        );

    \I__4011\ : CascadeMux
    port map (
            O => \N__18430\,
            I => \N__18422\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__18429\,
            I => \N__18419\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__18428\,
            I => \N__18416\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18425\,
            I => \N__18398\
        );

    \I__4007\ : InMux
    port map (
            O => \N__18422\,
            I => \N__18398\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18398\
        );

    \I__4005\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18398\
        );

    \I__4004\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18398\
        );

    \I__4003\ : InMux
    port map (
            O => \N__18414\,
            I => \N__18398\
        );

    \I__4002\ : InMux
    port map (
            O => \N__18413\,
            I => \N__18398\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__18398\,
            I => \N__18392\
        );

    \I__4000\ : InMux
    port map (
            O => \N__18397\,
            I => \N__18389\
        );

    \I__3999\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18386\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18383\
        );

    \I__3997\ : Span4Mux_h
    port map (
            O => \N__18392\,
            I => \N__18380\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18389\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__18386\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__18383\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3993\ : Odrv4
    port map (
            O => \N__18380\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18349\
        );

    \I__3991\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18349\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18369\,
            I => \N__18349\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18368\,
            I => \N__18349\
        );

    \I__3988\ : InMux
    port map (
            O => \N__18367\,
            I => \N__18349\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18366\,
            I => \N__18349\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18365\,
            I => \N__18349\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__18364\,
            I => \N__18341\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__18349\,
            I => \N__18338\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18331\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18331\
        );

    \I__3981\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18331\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18328\
        );

    \I__3979\ : InMux
    port map (
            O => \N__18344\,
            I => \N__18323\
        );

    \I__3978\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18323\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__18338\,
            I => \N__18320\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18331\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18328\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__18323\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3973\ : Odrv4
    port map (
            O => \N__18320\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__18311\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\
        );

    \I__3971\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18305\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__18305\,
            I => \N__18302\
        );

    \I__3969\ : Odrv4
    port map (
            O => \N__18302\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__3968\ : CascadeMux
    port map (
            O => \N__18299\,
            I => \uu2.mem0.bitmap_pmux_16_ns_1_cascade_\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__18293\,
            I => \N__18289\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18285\
        );

    \I__3964\ : Span4Mux_h
    port map (
            O => \N__18289\,
            I => \N__18281\
        );

    \I__3963\ : InMux
    port map (
            O => \N__18288\,
            I => \N__18278\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18275\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18284\,
            I => \N__18272\
        );

    \I__3960\ : Odrv4
    port map (
            O => \N__18281\,
            I => \uu2.N_30_i\
        );

    \I__3959\ : LocalMux
    port map (
            O => \N__18278\,
            I => \uu2.N_30_i\
        );

    \I__3958\ : Odrv12
    port map (
            O => \N__18275\,
            I => \uu2.N_30_i\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__18272\,
            I => \uu2.N_30_i\
        );

    \I__3956\ : CascadeMux
    port map (
            O => \N__18263\,
            I => \uu2.mem0.N_22_cascade_\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18260\,
            I => \N__18257\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18254\
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__18254\,
            I => \uu2.mem0.G_11_0_0_a3_6_0\
        );

    \I__3952\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18245\
        );

    \I__3951\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18245\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__18245\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__18242\,
            I => \N__18238\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18241\,
            I => \N__18232\
        );

    \I__3947\ : InMux
    port map (
            O => \N__18238\,
            I => \N__18227\
        );

    \I__3946\ : InMux
    port map (
            O => \N__18237\,
            I => \N__18227\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__18236\,
            I => \N__18223\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18220\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__18232\,
            I => \N__18215\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18215\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18226\,
            I => \N__18212\
        );

    \I__3940\ : InMux
    port map (
            O => \N__18223\,
            I => \N__18209\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18220\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__18215\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18212\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18209\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__3935\ : CascadeMux
    port map (
            O => \N__18200\,
            I => \N__18197\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18191\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18196\,
            I => \N__18191\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18191\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__3931\ : CascadeMux
    port map (
            O => \N__18188\,
            I => \N__18184\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18176\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18173\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18183\,
            I => \N__18170\
        );

    \I__3927\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18165\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18165\
        );

    \I__3925\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18160\
        );

    \I__3924\ : InMux
    port map (
            O => \N__18179\,
            I => \N__18160\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__18176\,
            I => \N__18157\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__18173\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__18170\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__18165\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__18160\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3918\ : Odrv4
    port map (
            O => \N__18157\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18140\
        );

    \I__3916\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18140\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__18140\,
            I => \N__18137\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__18137\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__3913\ : CascadeMux
    port map (
            O => \N__18134\,
            I => \uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_\
        );

    \I__3912\ : InMux
    port map (
            O => \N__18131\,
            I => \N__18127\
        );

    \I__3911\ : InMux
    port map (
            O => \N__18130\,
            I => \N__18124\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__18127\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__18124\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__18119\,
            I => \N__18108\
        );

    \I__3907\ : CascadeMux
    port map (
            O => \N__18118\,
            I => \N__18105\
        );

    \I__3906\ : CascadeMux
    port map (
            O => \N__18117\,
            I => \N__18099\
        );

    \I__3905\ : CascadeMux
    port map (
            O => \N__18116\,
            I => \N__18096\
        );

    \I__3904\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18091\
        );

    \I__3903\ : InMux
    port map (
            O => \N__18114\,
            I => \N__18091\
        );

    \I__3902\ : InMux
    port map (
            O => \N__18113\,
            I => \N__18088\
        );

    \I__3901\ : InMux
    port map (
            O => \N__18112\,
            I => \N__18081\
        );

    \I__3900\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18081\
        );

    \I__3899\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18081\
        );

    \I__3898\ : InMux
    port map (
            O => \N__18105\,
            I => \N__18076\
        );

    \I__3897\ : InMux
    port map (
            O => \N__18104\,
            I => \N__18076\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__18103\,
            I => \N__18073\
        );

    \I__3895\ : InMux
    port map (
            O => \N__18102\,
            I => \N__18069\
        );

    \I__3894\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18066\
        );

    \I__3893\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18063\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__18091\,
            I => \N__18060\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__18088\,
            I => \N__18053\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__18081\,
            I => \N__18053\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__18076\,
            I => \N__18053\
        );

    \I__3888\ : InMux
    port map (
            O => \N__18073\,
            I => \N__18050\
        );

    \I__3887\ : InMux
    port map (
            O => \N__18072\,
            I => \N__18047\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__18069\,
            I => \N__18042\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__18066\,
            I => \N__18042\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__18063\,
            I => \N__18033\
        );

    \I__3883\ : Span4Mux_v
    port map (
            O => \N__18060\,
            I => \N__18033\
        );

    \I__3882\ : Span4Mux_v
    port map (
            O => \N__18053\,
            I => \N__18033\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__18050\,
            I => \N__18033\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__18047\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3879\ : Odrv4
    port map (
            O => \N__18042\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3878\ : Odrv4
    port map (
            O => \N__18033\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__3877\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18022\
        );

    \I__3876\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18019\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__18022\,
            I => \N__18016\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__18019\,
            I => \uu2.N_30_i_1\
        );

    \I__3873\ : Odrv4
    port map (
            O => \N__18016\,
            I => \uu2.N_30_i_1\
        );

    \I__3872\ : CascadeMux
    port map (
            O => \N__18011\,
            I => \uu2.mem0.N_22_0_cascade_\
        );

    \I__3871\ : InMux
    port map (
            O => \N__18008\,
            I => \N__18005\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18005\,
            I => \N__18002\
        );

    \I__3869\ : Odrv12
    port map (
            O => \N__18002\,
            I => \uu2.N_104\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17996\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__17996\,
            I => \uu2.mem0.bitmap_pmux_27_ns_1_0\
        );

    \I__3866\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17978\
        );

    \I__3865\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17978\
        );

    \I__3864\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17978\
        );

    \I__3863\ : InMux
    port map (
            O => \N__17990\,
            I => \N__17973\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17989\,
            I => \N__17970\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17988\,
            I => \N__17963\
        );

    \I__3860\ : InMux
    port map (
            O => \N__17987\,
            I => \N__17963\
        );

    \I__3859\ : InMux
    port map (
            O => \N__17986\,
            I => \N__17963\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17985\,
            I => \N__17960\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__17978\,
            I => \N__17957\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17952\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17976\,
            I => \N__17952\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17973\,
            I => \N__17947\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17970\,
            I => \N__17947\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__17963\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__17960\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__17957\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17952\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__17947\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17933\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__17933\,
            I => \uu2.mem0.N_109\
        );

    \I__3845\ : InMux
    port map (
            O => \N__17930\,
            I => \N__17924\
        );

    \I__3844\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17924\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__17924\,
            I => \uu2.bitmap_pmux_19_ns_1\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__17921\,
            I => \N__17914\
        );

    \I__3841\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17905\
        );

    \I__3840\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17905\
        );

    \I__3839\ : InMux
    port map (
            O => \N__17918\,
            I => \N__17900\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17917\,
            I => \N__17891\
        );

    \I__3837\ : InMux
    port map (
            O => \N__17914\,
            I => \N__17891\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17913\,
            I => \N__17891\
        );

    \I__3835\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17891\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__17911\,
            I => \N__17885\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \N__17881\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__17905\,
            I => \N__17877\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__17904\,
            I => \N__17874\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17871\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17900\,
            I => \N__17866\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17891\,
            I => \N__17866\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__17890\,
            I => \N__17861\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__17889\,
            I => \N__17858\
        );

    \I__3825\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17855\
        );

    \I__3824\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17848\
        );

    \I__3823\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17848\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17848\
        );

    \I__3821\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17845\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__17877\,
            I => \N__17842\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17839\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__17871\,
            I => \N__17836\
        );

    \I__3817\ : Span4Mux_h
    port map (
            O => \N__17866\,
            I => \N__17833\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17824\
        );

    \I__3815\ : InMux
    port map (
            O => \N__17864\,
            I => \N__17824\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17824\
        );

    \I__3813\ : InMux
    port map (
            O => \N__17858\,
            I => \N__17824\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17855\,
            I => \N__17821\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__17848\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__17845\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__17842\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__17839\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__17836\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__17833\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17824\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__17821\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__17804\,
            I => \N__17801\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17795\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__17795\,
            I => \N__17792\
        );

    \I__3799\ : Span4Mux_s3_h
    port map (
            O => \N__17792\,
            I => \N__17789\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__17789\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__17786\,
            I => \N__17782\
        );

    \I__3796\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17777\
        );

    \I__3795\ : InMux
    port map (
            O => \N__17782\,
            I => \N__17777\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17777\,
            I => \N__17774\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__17774\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17768\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17768\,
            I => \uu2.mem0.N_109_0\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17765\,
            I => \N__17759\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__17764\,
            I => \N__17754\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__17763\,
            I => \N__17751\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17762\,
            I => \N__17745\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17759\,
            I => \N__17742\
        );

    \I__3785\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17738\
        );

    \I__3784\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17735\
        );

    \I__3783\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17728\
        );

    \I__3782\ : InMux
    port map (
            O => \N__17751\,
            I => \N__17728\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17750\,
            I => \N__17728\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17723\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17723\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17745\,
            I => \N__17718\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__17742\,
            I => \N__17718\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17715\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__17738\,
            I => \N__17710\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17735\,
            I => \N__17710\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17728\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__17723\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__17718\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17715\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__3769\ : Odrv4
    port map (
            O => \N__17710\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__17699\,
            I => \N__17696\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17696\,
            I => \N__17693\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__17693\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__3765\ : InMux
    port map (
            O => \N__17690\,
            I => \N__17687\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17687\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__17684\,
            I => \uu2.bitmap_pmux_20_ns_1_cascade_\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17681\,
            I => \N__17678\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17678\,
            I => \N__17675\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__17675\,
            I => \uu2.mem0.N_108\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17672\,
            I => \N__17666\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17671\,
            I => \N__17666\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17666\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17663\,
            I => \N__17657\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17662\,
            I => \N__17657\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__17657\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17651\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17651\,
            I => \uu2.bitmap_pmux_20_ns_1\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__17648\,
            I => \uu2.mem0.N_108_0_cascade_\
        );

    \I__3750\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17642\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17642\,
            I => \N__17639\
        );

    \I__3748\ : Span4Mux_h
    port map (
            O => \N__17639\,
            I => \N__17636\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__17636\,
            I => \uu2.mem0.N_404_0\
        );

    \I__3746\ : CascadeMux
    port map (
            O => \N__17633\,
            I => \N__17624\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17632\,
            I => \N__17619\
        );

    \I__3744\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17619\
        );

    \I__3743\ : CascadeMux
    port map (
            O => \N__17630\,
            I => \N__17616\
        );

    \I__3742\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17612\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17609\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17627\,
            I => \N__17606\
        );

    \I__3739\ : InMux
    port map (
            O => \N__17624\,
            I => \N__17603\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17619\,
            I => \N__17600\
        );

    \I__3737\ : InMux
    port map (
            O => \N__17616\,
            I => \N__17597\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17615\,
            I => \N__17594\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17612\,
            I => \N__17591\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__17609\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17606\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__17603\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__17600\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__17597\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17594\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__17591\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__17576\,
            I => \uu2.N_104_cascade_\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__17573\,
            I => \uu2.mem0.G_11_0_0_a3_5_0_cascade_\
        );

    \I__3725\ : InMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17567\,
            I => \uu2.mem0.N_40\
        );

    \I__3723\ : InMux
    port map (
            O => \N__17564\,
            I => \N__17561\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__17561\,
            I => \uu2.mem0.N_30\
        );

    \I__3721\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17552\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17552\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17552\,
            I => \N__17548\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17542\
        );

    \I__3717\ : Span4Mux_h
    port map (
            O => \N__17548\,
            I => \N__17538\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17531\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17531\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17531\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__17542\,
            I => \N__17528\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17541\,
            I => \N__17525\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__17538\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17531\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3709\ : Odrv4
    port map (
            O => \N__17528\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17525\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17516\,
            I => \N__17508\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17508\
        );

    \I__3705\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17501\
        );

    \I__3704\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17501\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17508\,
            I => \N__17498\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17507\,
            I => \N__17493\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17506\,
            I => \N__17493\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__17501\,
            I => \N__17477\
        );

    \I__3699\ : Span4Mux_v
    port map (
            O => \N__17498\,
            I => \N__17477\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__17493\,
            I => \N__17477\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17473\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17491\,
            I => \N__17468\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17490\,
            I => \N__17468\
        );

    \I__3694\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17459\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17459\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17459\
        );

    \I__3691\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17459\
        );

    \I__3690\ : InMux
    port map (
            O => \N__17485\,
            I => \N__17454\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17454\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__17477\,
            I => \N__17451\
        );

    \I__3687\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17448\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__17473\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17468\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17459\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17454\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__17451\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__17448\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__3680\ : InMux
    port map (
            O => \N__17435\,
            I => \N__17432\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__17432\,
            I => \N__17429\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__17429\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_41\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17426\,
            I => \N__17411\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17425\,
            I => \N__17411\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17424\,
            I => \N__17411\
        );

    \I__3674\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17406\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17422\,
            I => \N__17406\
        );

    \I__3672\ : InMux
    port map (
            O => \N__17421\,
            I => \N__17403\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17420\,
            I => \N__17400\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17397\
        );

    \I__3669\ : CascadeMux
    port map (
            O => \N__17418\,
            I => \N__17392\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__17411\,
            I => \N__17382\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__17406\,
            I => \N__17382\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__17403\,
            I => \N__17379\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__17400\,
            I => \N__17374\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17397\,
            I => \N__17374\
        );

    \I__3663\ : InMux
    port map (
            O => \N__17396\,
            I => \N__17369\
        );

    \I__3662\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17369\
        );

    \I__3661\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17366\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17359\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17359\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17359\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17354\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17354\
        );

    \I__3655\ : Span4Mux_h
    port map (
            O => \N__17382\,
            I => \N__17351\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__17379\,
            I => \N__17344\
        );

    \I__3653\ : Span4Mux_v
    port map (
            O => \N__17374\,
            I => \N__17344\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__17369\,
            I => \N__17344\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__17366\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17359\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17354\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__17351\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__17344\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17333\,
            I => \N__17329\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17332\,
            I => \N__17326\
        );

    \I__3644\ : LocalMux
    port map (
            O => \N__17329\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17326\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__17321\,
            I => \N__17317\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17307\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17307\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17316\,
            I => \N__17307\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__17315\,
            I => \N__17304\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__17314\,
            I => \N__17299\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__17307\,
            I => \N__17293\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17282\
        );

    \I__3634\ : InMux
    port map (
            O => \N__17303\,
            I => \N__17282\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17282\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17282\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17282\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17297\,
            I => \N__17276\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17296\,
            I => \N__17276\
        );

    \I__3628\ : Span4Mux_h
    port map (
            O => \N__17293\,
            I => \N__17271\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17271\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17268\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17276\,
            I => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5\
        );

    \I__3624\ : Odrv4
    port map (
            O => \N__17271\,
            I => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17268\,
            I => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17261\,
            I => \N__17258\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__17258\,
            I => \N__17250\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17243\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17256\,
            I => \N__17243\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17255\,
            I => \N__17240\
        );

    \I__3617\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17237\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17234\
        );

    \I__3615\ : Span4Mux_h
    port map (
            O => \N__17250\,
            I => \N__17231\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17228\
        );

    \I__3613\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17225\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__17243\,
            I => \N__17222\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17240\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__17237\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__17234\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3608\ : Odrv4
    port map (
            O => \N__17231\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17228\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__17225\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__17222\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__17207\,
            I => \N__17199\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__17206\,
            I => \N__17196\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17189\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17204\,
            I => \N__17189\
        );

    \I__3600\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17189\
        );

    \I__3599\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17186\
        );

    \I__3598\ : InMux
    port map (
            O => \N__17199\,
            I => \N__17181\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17196\,
            I => \N__17181\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__17189\,
            I => \N__17175\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17166\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__17181\,
            I => \N__17166\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17180\,
            I => \N__17161\
        );

    \I__3592\ : InMux
    port map (
            O => \N__17179\,
            I => \N__17161\
        );

    \I__3591\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17158\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__17175\,
            I => \N__17155\
        );

    \I__3589\ : InMux
    port map (
            O => \N__17174\,
            I => \N__17152\
        );

    \I__3588\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17147\
        );

    \I__3587\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17147\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17171\,
            I => \N__17144\
        );

    \I__3585\ : Span4Mux_h
    port map (
            O => \N__17166\,
            I => \N__17139\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__17161\,
            I => \N__17139\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17158\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__17155\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__17152\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__17147\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__17144\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__17139\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3577\ : InMux
    port map (
            O => \N__17126\,
            I => \N__17123\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__17123\,
            I => \uu2.mem0.G_11_0_0_a2_3_4\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__17120\,
            I => \N__17114\
        );

    \I__3574\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17111\
        );

    \I__3573\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17104\
        );

    \I__3572\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17104\
        );

    \I__3571\ : InMux
    port map (
            O => \N__17114\,
            I => \N__17104\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__17111\,
            I => \N__17099\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__17104\,
            I => \N__17099\
        );

    \I__3568\ : Span4Mux_s3_v
    port map (
            O => \N__17099\,
            I => \N__17096\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__17096\,
            I => \N_272_mux\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__17093\,
            I => \uu2.mem0.G_11_0_0_a2_3_5_cascade_\
        );

    \I__3565\ : InMux
    port map (
            O => \N__17090\,
            I => \N__17087\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__17087\,
            I => \N__17083\
        );

    \I__3563\ : InMux
    port map (
            O => \N__17086\,
            I => \N__17080\
        );

    \I__3562\ : Span4Mux_s3_h
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__3560\ : Span4Mux_h
    port map (
            O => \N__17077\,
            I => \N__17070\
        );

    \I__3559\ : Span4Mux_h
    port map (
            O => \N__17074\,
            I => \N__17067\
        );

    \I__3558\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17064\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__17070\,
            I => \L3_tx_data_1\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__17067\,
            I => \L3_tx_data_1\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__17064\,
            I => \L3_tx_data_1\
        );

    \I__3554\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17054\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__17054\,
            I => \uu2.mem0.G_11_0_0_0\
        );

    \I__3552\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17048\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__17048\,
            I => \N__17045\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__17045\,
            I => \N__17042\
        );

    \I__3549\ : Odrv4
    port map (
            O => \N__17042\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_1\
        );

    \I__3548\ : InMux
    port map (
            O => \N__17039\,
            I => \N__17036\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17036\,
            I => \N__17033\
        );

    \I__3546\ : Span4Mux_v
    port map (
            O => \N__17033\,
            I => \N__17030\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__17030\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_5\
        );

    \I__3544\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17024\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__17024\,
            I => \N__17021\
        );

    \I__3542\ : Span4Mux_h
    port map (
            O => \N__17021\,
            I => \N__17018\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__17018\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_4\
        );

    \I__3540\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17012\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__17012\,
            I => \N__17009\
        );

    \I__3538\ : Span4Mux_h
    port map (
            O => \N__17009\,
            I => \N__17006\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__17006\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_2\
        );

    \I__3536\ : InMux
    port map (
            O => \N__17003\,
            I => \N__17000\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__17000\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__16997\,
            I => \N__16994\
        );

    \I__3533\ : InMux
    port map (
            O => \N__16994\,
            I => \N__16991\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16991\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__3531\ : InMux
    port map (
            O => \N__16988\,
            I => \N__16985\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__16985\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16982\,
            I => \N__16979\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__16979\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \uu2.bitmap_pmux_17_ns_1_cascade_\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__16973\,
            I => \N__16963\
        );

    \I__3525\ : CascadeMux
    port map (
            O => \N__16972\,
            I => \N__16958\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__16971\,
            I => \N__16954\
        );

    \I__3523\ : InMux
    port map (
            O => \N__16970\,
            I => \N__16951\
        );

    \I__3522\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16946\
        );

    \I__3521\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16943\
        );

    \I__3520\ : InMux
    port map (
            O => \N__16967\,
            I => \N__16940\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__16966\,
            I => \N__16937\
        );

    \I__3518\ : InMux
    port map (
            O => \N__16963\,
            I => \N__16932\
        );

    \I__3517\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16932\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16923\
        );

    \I__3515\ : InMux
    port map (
            O => \N__16958\,
            I => \N__16923\
        );

    \I__3514\ : InMux
    port map (
            O => \N__16957\,
            I => \N__16923\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16954\,
            I => \N__16923\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16951\,
            I => \N__16920\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16950\,
            I => \N__16917\
        );

    \I__3510\ : InMux
    port map (
            O => \N__16949\,
            I => \N__16914\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16946\,
            I => \N__16909\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__16943\,
            I => \N__16909\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__16940\,
            I => \N__16906\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16903\
        );

    \I__3505\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16900\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__16923\,
            I => \N__16891\
        );

    \I__3503\ : Span4Mux_h
    port map (
            O => \N__16920\,
            I => \N__16891\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__16917\,
            I => \N__16891\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__16914\,
            I => \N__16891\
        );

    \I__3500\ : Span4Mux_v
    port map (
            O => \N__16909\,
            I => \N__16886\
        );

    \I__3499\ : Span4Mux_v
    port map (
            O => \N__16906\,
            I => \N__16886\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16903\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3497\ : Odrv12
    port map (
            O => \N__16900\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__16891\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__16886\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__16877\,
            I => \Lab_UT.dictrl.g0_8Z0Z_3_cascade_\
        );

    \I__3493\ : CascadeMux
    port map (
            O => \N__16874\,
            I => \N__16871\
        );

    \I__3492\ : InMux
    port map (
            O => \N__16871\,
            I => \N__16868\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16868\,
            I => \N__16865\
        );

    \I__3490\ : Odrv4
    port map (
            O => \N__16865\,
            I => \Lab_UT.dictrl.g2_1_3\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16854\
        );

    \I__3488\ : InMux
    port map (
            O => \N__16861\,
            I => \N__16854\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16851\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16859\,
            I => \N__16848\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__16854\,
            I => \N__16843\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__16851\,
            I => \N__16843\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16848\,
            I => bu_rx_data_1_rep1
        );

    \I__3482\ : Odrv4
    port map (
            O => \N__16843\,
            I => bu_rx_data_1_rep1
        );

    \I__3481\ : InMux
    port map (
            O => \N__16838\,
            I => \N__16835\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16835\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_28\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16829\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__16829\,
            I => \uu2.mem0.N_44\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__16826\,
            I => \uu2.mem0.N_41_cascade_\
        );

    \I__3476\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16820\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16820\,
            I => \N__16817\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__16817\,
            I => \N__16814\
        );

    \I__3473\ : Odrv4
    port map (
            O => \N__16814\,
            I => \uu2.mem0.w_data_1\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16811\,
            I => \N__16805\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16805\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__16805\,
            I => \N__16802\
        );

    \I__3469\ : Span4Mux_h
    port map (
            O => \N__16802\,
            I => \N__16798\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16801\,
            I => \N__16795\
        );

    \I__3467\ : Odrv4
    port map (
            O => \N__16798\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__16795\,
            I => \uu2.bitmap_pmux_sn_N_36\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__16790\,
            I => \uu2.mem0.N_24_i_cascade_\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16787\,
            I => \N__16782\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16779\
        );

    \I__3462\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16776\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16773\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16779\,
            I => \uu2.N_406\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16776\,
            I => \uu2.N_406\
        );

    \I__3458\ : Odrv12
    port map (
            O => \N__16773\,
            I => \uu2.N_406\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16766\,
            I => \N__16763\
        );

    \I__3456\ : LocalMux
    port map (
            O => \N__16763\,
            I => \uu2.mem0.N_45\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16757\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__16757\,
            I => \N__16754\
        );

    \I__3453\ : Odrv12
    port map (
            O => \N__16754\,
            I => \Lab_UT.dictrl.next_alarmstate4Z0Z_3\
        );

    \I__3452\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16748\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16748\,
            I => \N__16745\
        );

    \I__3450\ : Odrv4
    port map (
            O => \N__16745\,
            I => \Lab_UT.dictrl.next_alarmstate4Z0Z_0\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16742\,
            I => \N__16739\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16739\,
            I => \Lab_UT.dictrl.g2_1_2\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__16736\,
            I => \Lab_UT.dictrl.g1_5_1_cascade_\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16730\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__16730\,
            I => \Lab_UT.dictrl.g2_3\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16727\,
            I => \N__16724\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16724\,
            I => \Lab_UT.dictrl.g0Z0Z_1\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__16721\,
            I => \Lab_UT.dictrl.g0_3_cascade_\
        );

    \I__3441\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16708\
        );

    \I__3440\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16703\
        );

    \I__3439\ : InMux
    port map (
            O => \N__16716\,
            I => \N__16703\
        );

    \I__3438\ : InMux
    port map (
            O => \N__16715\,
            I => \N__16696\
        );

    \I__3437\ : InMux
    port map (
            O => \N__16714\,
            I => \N__16696\
        );

    \I__3436\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16696\
        );

    \I__3435\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16691\
        );

    \I__3434\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16691\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__16708\,
            I => bu_rx_data_5_rep1
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__16703\,
            I => bu_rx_data_5_rep1
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__16696\,
            I => bu_rx_data_5_rep1
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__16691\,
            I => bu_rx_data_5_rep1
        );

    \I__3429\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16676\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16676\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__16676\,
            I => \N__16673\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__16673\,
            I => \Lab_UT.dictrl.next_state12_0\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__16670\,
            I => \N__16665\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16669\,
            I => \N__16660\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__16668\,
            I => \N__16656\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16647\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16647\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16647\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16660\,
            I => \N__16644\
        );

    \I__3418\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16637\
        );

    \I__3417\ : InMux
    port map (
            O => \N__16656\,
            I => \N__16637\
        );

    \I__3416\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16637\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16654\,
            I => \N__16634\
        );

    \I__3414\ : LocalMux
    port map (
            O => \N__16647\,
            I => \N__16631\
        );

    \I__3413\ : Odrv4
    port map (
            O => \N__16644\,
            I => bu_rx_data_6_rep1
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16637\,
            I => bu_rx_data_6_rep1
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__16634\,
            I => bu_rx_data_6_rep1
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__16631\,
            I => bu_rx_data_6_rep1
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__16622\,
            I => \N__16619\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16616\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16616\,
            I => \Lab_UT.dictrl.g0_0_0_o4_0\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16613\,
            I => \Lab_UT.dictrl.N_3_0_cascade_\
        );

    \I__3405\ : InMux
    port map (
            O => \N__16610\,
            I => \N__16607\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__16607\,
            I => \Lab_UT.dictrl.g0_0_0_a3_2_0\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16604\,
            I => \N__16601\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16601\,
            I => \N__16598\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__16598\,
            I => \Lab_UT.dictrl.g0_0_i_o4_0\
        );

    \I__3400\ : InMux
    port map (
            O => \N__16595\,
            I => \N__16584\
        );

    \I__3399\ : InMux
    port map (
            O => \N__16594\,
            I => \N__16584\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16584\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16579\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16591\,
            I => \N__16579\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__16584\,
            I => \N__16573\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__16579\,
            I => \N__16570\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16578\,
            I => \N__16563\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16577\,
            I => \N__16563\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16563\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__16573\,
            I => \Lab_UT.dictrl.g0_1Z0Z_2\
        );

    \I__3389\ : Odrv4
    port map (
            O => \N__16570\,
            I => \Lab_UT.dictrl.g0_1Z0Z_2\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16563\,
            I => \Lab_UT.dictrl.g0_1Z0Z_2\
        );

    \I__3387\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16553\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16553\,
            I => \Lab_UT.dictrl.next_state18_0\
        );

    \I__3385\ : CascadeMux
    port map (
            O => \N__16550\,
            I => \Lab_UT.dictrl.next_state18_0_cascade_\
        );

    \I__3384\ : CascadeMux
    port map (
            O => \N__16547\,
            I => \Lab_UT.dictrl.g2_0_0_cascade_\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16544\,
            I => \N__16541\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16541\,
            I => \Lab_UT.dictrl.N_7_0\
        );

    \I__3381\ : InMux
    port map (
            O => \N__16538\,
            I => \N__16535\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16535\,
            I => \N__16532\
        );

    \I__3379\ : Odrv12
    port map (
            O => \N__16532\,
            I => \Lab_UT.dictrl.N_11\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16529\,
            I => \N__16526\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16526\,
            I => \Lab_UT.dictrl.g2_2_0\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16523\,
            I => \N__16520\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__16520\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_3_0\
        );

    \I__3374\ : InMux
    port map (
            O => \N__16517\,
            I => \N__16514\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16514\,
            I => \N__16511\
        );

    \I__3372\ : Odrv4
    port map (
            O => \N__16511\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_4\
        );

    \I__3371\ : InMux
    port map (
            O => \N__16508\,
            I => \N__16505\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16502\
        );

    \I__3369\ : Sp12to4
    port map (
            O => \N__16502\,
            I => \N__16499\
        );

    \I__3368\ : Odrv12
    port map (
            O => \N__16499\,
            I => \Lab_UT.dictrl.N_9_0\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__16496\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16483\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16492\,
            I => \N__16483\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16479\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16476\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16471\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16468\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16465\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16482\,
            I => \N__16462\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16479\,
            I => \N__16459\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__16476\,
            I => \N__16456\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16451\
        );

    \I__3355\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16451\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__16471\,
            I => \N__16447\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__16468\,
            I => \N__16440\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__16465\,
            I => \N__16440\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16440\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__16459\,
            I => \N__16435\
        );

    \I__3349\ : Span4Mux_v
    port map (
            O => \N__16456\,
            I => \N__16435\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__16451\,
            I => \N__16432\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16450\,
            I => \N__16429\
        );

    \I__3346\ : Span4Mux_h
    port map (
            O => \N__16447\,
            I => \N__16424\
        );

    \I__3345\ : Span4Mux_h
    port map (
            O => \N__16440\,
            I => \N__16424\
        );

    \I__3344\ : Odrv4
    port map (
            O => \N__16435\,
            I => bu_rx_data_0
        );

    \I__3343\ : Odrv12
    port map (
            O => \N__16432\,
            I => bu_rx_data_0
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16429\,
            I => bu_rx_data_0
        );

    \I__3341\ : Odrv4
    port map (
            O => \N__16424\,
            I => bu_rx_data_0
        );

    \I__3340\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16409\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16409\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__3337\ : Span4Mux_h
    port map (
            O => \N__16406\,
            I => \N__16403\
        );

    \I__3336\ : Odrv4
    port map (
            O => \N__16403\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z4\
        );

    \I__3335\ : CascadeMux
    port map (
            O => \N__16400\,
            I => \Lab_UT.dictrl.N_5_cascade_\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16394\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__16394\,
            I => \Lab_UT.dictrl.N_10_0\
        );

    \I__3332\ : CascadeMux
    port map (
            O => \N__16391\,
            I => \N__16386\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__16390\,
            I => \N__16382\
        );

    \I__3330\ : InMux
    port map (
            O => \N__16389\,
            I => \N__16375\
        );

    \I__3329\ : InMux
    port map (
            O => \N__16386\,
            I => \N__16375\
        );

    \I__3328\ : InMux
    port map (
            O => \N__16385\,
            I => \N__16375\
        );

    \I__3327\ : InMux
    port map (
            O => \N__16382\,
            I => \N__16372\
        );

    \I__3326\ : LocalMux
    port map (
            O => \N__16375\,
            I => \N__16369\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__16372\,
            I => \N__16366\
        );

    \I__3324\ : Span12Mux_s7_h
    port map (
            O => \N__16369\,
            I => \N__16363\
        );

    \I__3323\ : Span4Mux_v
    port map (
            O => \N__16366\,
            I => \N__16360\
        );

    \I__3322\ : Odrv12
    port map (
            O => \N__16363\,
            I => \Lab_UT.dicRun_2\
        );

    \I__3321\ : Odrv4
    port map (
            O => \N__16360\,
            I => \Lab_UT.dicRun_2\
        );

    \I__3320\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16352\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16352\,
            I => \Lab_UT.didp.ce_9_0_0\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__16349\,
            I => \Lab_UT.dicRun_2_cascade_\
        );

    \I__3317\ : InMux
    port map (
            O => \N__16346\,
            I => \N__16341\
        );

    \I__3316\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16338\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16331\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16326\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16338\,
            I => \N__16326\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16323\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16318\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16335\,
            I => \N__16318\
        );

    \I__3309\ : InMux
    port map (
            O => \N__16334\,
            I => \N__16313\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16331\,
            I => \N__16310\
        );

    \I__3307\ : Span4Mux_v
    port map (
            O => \N__16326\,
            I => \N__16305\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__16323\,
            I => \N__16305\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16318\,
            I => \N__16302\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16317\,
            I => \N__16294\
        );

    \I__3303\ : InMux
    port map (
            O => \N__16316\,
            I => \N__16294\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__16313\,
            I => \N__16289\
        );

    \I__3301\ : Span4Mux_v
    port map (
            O => \N__16310\,
            I => \N__16286\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__16305\,
            I => \N__16281\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__16302\,
            I => \N__16281\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16301\,
            I => \N__16274\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16300\,
            I => \N__16274\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16299\,
            I => \N__16274\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__16294\,
            I => \N__16271\
        );

    \I__3294\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16266\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16266\
        );

    \I__3292\ : Span4Mux_v
    port map (
            O => \N__16289\,
            I => \N__16259\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__16286\,
            I => \N__16259\
        );

    \I__3290\ : Span4Mux_v
    port map (
            O => \N__16281\,
            I => \N__16259\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__16274\,
            I => \oneSecStrb\
        );

    \I__3288\ : Odrv4
    port map (
            O => \N__16271\,
            I => \oneSecStrb\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16266\,
            I => \oneSecStrb\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__16259\,
            I => \oneSecStrb\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16240\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16240\
        );

    \I__3283\ : InMux
    port map (
            O => \N__16248\,
            I => \N__16240\
        );

    \I__3282\ : InMux
    port map (
            O => \N__16247\,
            I => \N__16237\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16237\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__16234\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__3278\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16226\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16226\,
            I => \Lab_UT.dictrl.N_11_0\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__16223\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_\
        );

    \I__3275\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16217\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__16217\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_1\
        );

    \I__3273\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16211\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16211\,
            I => \Lab_UT.dictrl.g0_0_i_a3_3_1\
        );

    \I__3271\ : InMux
    port map (
            O => \N__16208\,
            I => \N__16205\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__16205\,
            I => \Lab_UT.bcd2segment3.segment_0Z0Z_2\
        );

    \I__3269\ : InMux
    port map (
            O => \N__16202\,
            I => \N__16199\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__16199\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_4\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__16193\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_6\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16187\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__16187\,
            I => \N__16184\
        );

    \I__3263\ : Odrv12
    port map (
            O => \N__16184\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__3262\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16178\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16178\,
            I => \Lab_UT.bcd2segment3.segment_0Z0Z_1\
        );

    \I__3260\ : InMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__16172\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_5\
        );

    \I__3258\ : InMux
    port map (
            O => \N__16169\,
            I => \N__16166\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16166\,
            I => \N__16163\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__16163\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__3255\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16157\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__16157\,
            I => \N__16154\
        );

    \I__3253\ : Span4Mux_h
    port map (
            O => \N__16154\,
            I => \N__16151\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__16151\,
            I => \Lab_UT.LdASones\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__16148\,
            I => \Lab_UT.LdASones_cascade_\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16142\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__16142\,
            I => \N__16139\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__16139\,
            I => \N__16136\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__16136\,
            I => \Lab_UT.LdSones_i_3\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16133\,
            I => \N__16130\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__16130\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__3244\ : InMux
    port map (
            O => \N__16127\,
            I => \N__16122\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__16126\,
            I => \N__16110\
        );

    \I__3242\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16106\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16103\
        );

    \I__3240\ : InMux
    port map (
            O => \N__16121\,
            I => \N__16100\
        );

    \I__3239\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16095\
        );

    \I__3238\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16095\
        );

    \I__3237\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16090\
        );

    \I__3236\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16090\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16116\,
            I => \N__16083\
        );

    \I__3234\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16083\
        );

    \I__3233\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16083\
        );

    \I__3232\ : InMux
    port map (
            O => \N__16113\,
            I => \N__16076\
        );

    \I__3231\ : InMux
    port map (
            O => \N__16110\,
            I => \N__16076\
        );

    \I__3230\ : InMux
    port map (
            O => \N__16109\,
            I => \N__16076\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__16106\,
            I => \N__16073\
        );

    \I__3228\ : Odrv4
    port map (
            O => \N__16103\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__16100\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__16095\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16090\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__16083\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__16076\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3222\ : Odrv4
    port map (
            O => \N__16073\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__16058\,
            I => \uu2.N_98_cascade_\
        );

    \I__3220\ : InMux
    port map (
            O => \N__16055\,
            I => \N__16049\
        );

    \I__3219\ : InMux
    port map (
            O => \N__16054\,
            I => \N__16049\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16049\,
            I => \uu2.bitmap_RNI04AD1Z0Z_314\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__16046\,
            I => \N__16043\
        );

    \I__3216\ : InMux
    port map (
            O => \N__16043\,
            I => \N__16036\
        );

    \I__3215\ : InMux
    port map (
            O => \N__16042\,
            I => \N__16033\
        );

    \I__3214\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16028\
        );

    \I__3213\ : InMux
    port map (
            O => \N__16040\,
            I => \N__16028\
        );

    \I__3212\ : InMux
    port map (
            O => \N__16039\,
            I => \N__16025\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__16036\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__16033\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__16028\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__16025\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__3207\ : InMux
    port map (
            O => \N__16016\,
            I => \N__16013\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__16013\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__3205\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16004\
        );

    \I__3204\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16004\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__16004\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3202\ : InMux
    port map (
            O => \N__16001\,
            I => \N__15998\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15998\,
            I => \uu2.N_383\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__15995\,
            I => \N__15989\
        );

    \I__3199\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15974\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15993\,
            I => \N__15969\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15969\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15962\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15962\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15987\,
            I => \N__15962\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15986\,
            I => \N__15958\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15985\,
            I => \N__15955\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15952\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__15983\,
            I => \N__15949\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__15982\,
            I => \N__15944\
        );

    \I__3188\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15933\
        );

    \I__3187\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15933\
        );

    \I__3186\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15933\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15933\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15933\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15930\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__15969\,
            I => \N__15926\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__15962\,
            I => \N__15923\
        );

    \I__3180\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15920\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15958\,
            I => \N__15917\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__15955\,
            I => \N__15912\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__15952\,
            I => \N__15912\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15949\,
            I => \N__15903\
        );

    \I__3175\ : InMux
    port map (
            O => \N__15948\,
            I => \N__15903\
        );

    \I__3174\ : InMux
    port map (
            O => \N__15947\,
            I => \N__15903\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15903\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__15933\,
            I => \N__15898\
        );

    \I__3171\ : Span4Mux_s2_v
    port map (
            O => \N__15930\,
            I => \N__15898\
        );

    \I__3170\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15895\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__15926\,
            I => \N__15892\
        );

    \I__3168\ : Span4Mux_h
    port map (
            O => \N__15923\,
            I => \N__15889\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__15920\,
            I => \N__15886\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__15917\,
            I => \N__15881\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__15912\,
            I => \N__15881\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15876\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__15898\,
            I => \N__15876\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__15895\,
            I => \N__15873\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__15892\,
            I => \L3_tx_data_rdy\
        );

    \I__3160\ : Odrv4
    port map (
            O => \N__15889\,
            I => \L3_tx_data_rdy\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__15886\,
            I => \L3_tx_data_rdy\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__15881\,
            I => \L3_tx_data_rdy\
        );

    \I__3157\ : Odrv4
    port map (
            O => \N__15876\,
            I => \L3_tx_data_rdy\
        );

    \I__3156\ : Odrv12
    port map (
            O => \N__15873\,
            I => \L3_tx_data_rdy\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15845\
        );

    \I__3154\ : InMux
    port map (
            O => \N__15859\,
            I => \N__15845\
        );

    \I__3153\ : InMux
    port map (
            O => \N__15858\,
            I => \N__15845\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15845\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15841\
        );

    \I__3150\ : InMux
    port map (
            O => \N__15855\,
            I => \N__15832\
        );

    \I__3149\ : InMux
    port map (
            O => \N__15854\,
            I => \N__15829\
        );

    \I__3148\ : LocalMux
    port map (
            O => \N__15845\,
            I => \N__15822\
        );

    \I__3147\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15815\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15815\
        );

    \I__3145\ : InMux
    port map (
            O => \N__15840\,
            I => \N__15815\
        );

    \I__3144\ : InMux
    port map (
            O => \N__15839\,
            I => \N__15804\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15804\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15837\,
            I => \N__15804\
        );

    \I__3141\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15804\
        );

    \I__3140\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15804\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__15832\,
            I => \N__15800\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15829\,
            I => \N__15797\
        );

    \I__3137\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15794\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15789\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15789\
        );

    \I__3134\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15786\
        );

    \I__3133\ : Span4Mux_h
    port map (
            O => \N__15822\,
            I => \N__15783\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__15815\,
            I => \N__15778\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__15804\,
            I => \N__15778\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15803\,
            I => \N__15775\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__15800\,
            I => \N__15770\
        );

    \I__3128\ : Span4Mux_s2_v
    port map (
            O => \N__15797\,
            I => \N__15770\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__15794\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__15789\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15786\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__15783\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__15778\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__15775\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3121\ : Odrv4
    port map (
            O => \N__15770\,
            I => uu2_un1_w_user_cr_0
        );

    \I__3120\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15749\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15749\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__15749\,
            I => \N__15745\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15748\,
            I => \N__15742\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__15745\,
            I => \N__15738\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15735\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15741\,
            I => \N__15732\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__15738\,
            I => \uu2.N_57\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__15735\,
            I => \uu2.N_57\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__15732\,
            I => \uu2.N_57\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__15725\,
            I => \N__15719\
        );

    \I__3109\ : InMux
    port map (
            O => \N__15724\,
            I => \N__15709\
        );

    \I__3108\ : InMux
    port map (
            O => \N__15723\,
            I => \N__15709\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15722\,
            I => \N__15709\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15709\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__15718\,
            I => \N__15706\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15709\,
            I => \N__15703\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__3102\ : Span4Mux_h
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15700\,
            I => \uu2.N_38\
        );

    \I__3100\ : Odrv4
    port map (
            O => \N__15697\,
            I => \uu2.N_38\
        );

    \I__3099\ : CascadeMux
    port map (
            O => \N__15692\,
            I => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_\
        );

    \I__3098\ : CascadeMux
    port map (
            O => \N__15689\,
            I => \N__15686\
        );

    \I__3097\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15682\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \N__15675\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15682\,
            I => \N__15672\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15668\
        );

    \I__3093\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15659\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15659\
        );

    \I__3091\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15659\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15659\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__15672\,
            I => \N__15653\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15671\,
            I => \N__15650\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15668\,
            I => \N__15645\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15659\,
            I => \N__15645\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15658\,
            I => \N__15638\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15657\,
            I => \N__15638\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15656\,
            I => \N__15638\
        );

    \I__3082\ : Sp12to4
    port map (
            O => \N__15653\,
            I => \N__15633\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__15650\,
            I => \N__15633\
        );

    \I__3080\ : Span4Mux_h
    port map (
            O => \N__15645\,
            I => \N__15630\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__15638\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3078\ : Odrv12
    port map (
            O => \N__15633\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__15630\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15620\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__15620\,
            I => \uu2.bitmap_pmux_sn_N_54_mux\
        );

    \I__3074\ : InMux
    port map (
            O => \N__15617\,
            I => \N__15614\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15614\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__3072\ : CEMux
    port map (
            O => \N__15611\,
            I => \N__15608\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__15608\,
            I => \N__15604\
        );

    \I__3070\ : CEMux
    port map (
            O => \N__15607\,
            I => \N__15601\
        );

    \I__3069\ : Sp12to4
    port map (
            O => \N__15604\,
            I => \N__15598\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__15601\,
            I => \uu2.N_31_0\
        );

    \I__3067\ : Odrv12
    port map (
            O => \N__15598\,
            I => \uu2.N_31_0\
        );

    \I__3066\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15590\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15590\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15587\,
            I => \N__15584\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15584\,
            I => \N__15581\
        );

    \I__3062\ : Odrv12
    port map (
            O => \N__15581\,
            I => \uu2.mem0.N_36\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__15578\,
            I => \uu2.mem0.N_9_cascade_\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15575\,
            I => \N__15572\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15572\,
            I => \uu2.bitmap_pmux_26_bm_1\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15569\,
            I => \uu2.bitmap_RNI31F32Z0Z_34_cascade_\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__15563\,
            I => \uu2.w_addr_displaying_RNIBICU6_0Z0Z_2\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__15560\,
            I => \uu2.N_401_cascade_\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__15554\,
            I => \uu2.w_addr_displaying_RNIBICU6Z0Z_2\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__3050\ : Odrv4
    port map (
            O => \N__15545\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__3049\ : CascadeMux
    port map (
            O => \N__15542\,
            I => \uu2.N_99_cascade_\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15536\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__15536\,
            I => \uu2.bitmap_RNI2Q8F1Z0Z_111\
        );

    \I__3046\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15530\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15530\,
            I => \uu2.bitmap_pmux_sn_N_15\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__15527\,
            I => \N__15524\
        );

    \I__3043\ : InMux
    port map (
            O => \N__15524\,
            I => \N__15521\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15521\,
            I => bu_rx_data_fast_5
        );

    \I__3041\ : InMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15515\,
            I => bu_rx_data_fast_3
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__15512\,
            I => \uu2.mem0.N_98_0_cascade_\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15506\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__15506\,
            I => \uu2.mem0.G_11_0_0_a3_0_2\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__15503\,
            I => \uu2.mem0.N_62_cascade_\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__15500\,
            I => \Lab_UT.dictrl.g2_1_0_1_cascade_\
        );

    \I__3034\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__15494\,
            I => \Lab_UT.dictrl.N_7_1_0\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__3031\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15484\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15487\,
            I => \N__15481\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15484\,
            I => \N__15478\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__15481\,
            I => bu_rx_data_fast_4
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__15478\,
            I => bu_rx_data_fast_4
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__15473\,
            I => \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15467\,
            I => \Lab_UT.dictrl.next_state18_1_0\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__15464\,
            I => \Lab_UT.dictrl.g1_0_1_cascade_\
        );

    \I__3022\ : InMux
    port map (
            O => \N__15461\,
            I => \N__15458\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15458\,
            I => \Lab_UT.dictrl.g2_1\
        );

    \I__3020\ : InMux
    port map (
            O => \N__15455\,
            I => \N__15449\
        );

    \I__3019\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15446\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15441\
        );

    \I__3017\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15441\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__15449\,
            I => \N__15437\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__15446\,
            I => \N__15432\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__15441\,
            I => \N__15432\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15429\
        );

    \I__3012\ : Span4Mux_h
    port map (
            O => \N__15437\,
            I => \N__15426\
        );

    \I__3011\ : Span4Mux_v
    port map (
            O => \N__15432\,
            I => \N__15421\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__15429\,
            I => \N__15421\
        );

    \I__3009\ : Odrv4
    port map (
            O => \N__15426\,
            I => \Lab_UT.LdMones\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__15421\,
            I => \Lab_UT.LdMones\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15416\,
            I => \Lab_UT.dictrl.g0_1_2_0_cascade_\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__15413\,
            I => \Lab_UT.dictrl.N_29_0_0_cascade_\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15407\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__15407\,
            I => \Lab_UT.dictrl.N_30_0\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15404\,
            I => \Lab_UT.dictrl.N_30_0_cascade_\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15395\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15395\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__15395\,
            I => \Lab_UT.dictrl.i6_mux_0\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15389\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15389\,
            I => \N__15386\
        );

    \I__2997\ : Odrv4
    port map (
            O => \N__15386\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__15383\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__15380\,
            I => \Lab_UT.dictrl.dicLdAMones_0_sx_cascade_\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__15377\,
            I => \N__15373\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15368\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15368\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__15368\,
            I => \N__15365\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__15365\,
            I => \Lab_UT.dicLdAMones_1\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__15362\,
            I => \N__15359\
        );

    \I__2988\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15356\
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__15356\,
            I => \Lab_UT.dictrl.g0_1_3\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__15353\,
            I => \N__15349\
        );

    \I__2985\ : InMux
    port map (
            O => \N__15352\,
            I => \N__15344\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15349\,
            I => \N__15344\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__15344\,
            I => \N__15341\
        );

    \I__2982\ : Odrv4
    port map (
            O => \N__15341\,
            I => \Lab_UT.dicLdSones_1\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__15338\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__15335\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__15332\,
            I => \Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_\
        );

    \I__2978\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15326\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__15326\,
            I => \Lab_UT.dictrl.g0_0_i_a3_2\
        );

    \I__2976\ : CascadeMux
    port map (
            O => \N__15323\,
            I => \Lab_UT.dictrl.g3_0_cascade_\
        );

    \I__2975\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15317\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__15317\,
            I => \Lab_UT.dictrl.g0_0_0_a3_2\
        );

    \I__2973\ : CascadeMux
    port map (
            O => \N__15314\,
            I => \Lab_UT.didp.countrce1.q_5_2_cascade_\
        );

    \I__2972\ : CascadeMux
    port map (
            O => \N__15311\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15308\,
            I => \N__15296\
        );

    \I__2970\ : InMux
    port map (
            O => \N__15307\,
            I => \N__15296\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15296\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15296\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__15296\,
            I => \N__15293\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__15293\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__15290\,
            I => \Lab_UT.didp.countrce1.q_5_3_cascade_\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__15287\,
            I => \N__15284\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15281\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15281\,
            I => \N__15278\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__15278\,
            I => \Lab_UT.didp.countrce1.q_5_1\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__15275\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__15272\,
            I => \Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__15269\,
            I => \N__15264\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__15268\,
            I => \N__15260\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15257\
        );

    \I__2955\ : InMux
    port map (
            O => \N__15264\,
            I => \N__15252\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15263\,
            I => \N__15252\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15249\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15257\,
            I => \Lab_UT.LdSones\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__15252\,
            I => \Lab_UT.LdSones\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__15249\,
            I => \Lab_UT.LdSones\
        );

    \I__2949\ : CascadeMux
    port map (
            O => \N__15242\,
            I => \Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__15233\,
            I => \Lab_UT.bcd2segment3.segment_0Z0Z_0\
        );

    \I__2945\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15224\
        );

    \I__2944\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15224\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__15224\,
            I => \N__15209\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15206\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15203\
        );

    \I__2940\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15200\
        );

    \I__2939\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15195\
        );

    \I__2938\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15195\
        );

    \I__2937\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15180\
        );

    \I__2936\ : InMux
    port map (
            O => \N__15217\,
            I => \N__15180\
        );

    \I__2935\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15180\
        );

    \I__2934\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15180\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15214\,
            I => \N__15180\
        );

    \I__2932\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15180\
        );

    \I__2931\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15180\
        );

    \I__2930\ : Span4Mux_h
    port map (
            O => \N__15209\,
            I => \N__15175\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__15206\,
            I => \N__15175\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__15203\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__15200\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__15195\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__15180\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__15175\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2923\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15143\
        );

    \I__2922\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15143\
        );

    \I__2921\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15143\
        );

    \I__2920\ : InMux
    port map (
            O => \N__15161\,
            I => \N__15143\
        );

    \I__2919\ : InMux
    port map (
            O => \N__15160\,
            I => \N__15143\
        );

    \I__2918\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15143\
        );

    \I__2917\ : InMux
    port map (
            O => \N__15158\,
            I => \N__15143\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__15143\,
            I => \N__15136\
        );

    \I__2915\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15131\
        );

    \I__2914\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15131\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15126\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15139\,
            I => \N__15126\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__15136\,
            I => \N__15123\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__15131\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__15126\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__2908\ : Odrv4
    port map (
            O => \N__15123\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__15116\,
            I => \N__15106\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__15115\,
            I => \N__15103\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__15114\,
            I => \N__15100\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__15113\,
            I => \N__15097\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__15112\,
            I => \N__15094\
        );

    \I__2902\ : CascadeMux
    port map (
            O => \N__15111\,
            I => \N__15091\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__15110\,
            I => \N__15088\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__15109\,
            I => \N__15083\
        );

    \I__2899\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15076\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15103\,
            I => \N__15076\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15076\
        );

    \I__2896\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15067\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15067\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15091\,
            I => \N__15067\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15088\,
            I => \N__15067\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15087\,
            I => \N__15064\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15059\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15083\,
            I => \N__15059\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15054\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15054\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__15064\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__15059\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__15054\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__15047\,
            I => \N__15043\
        );

    \I__2883\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15037\
        );

    \I__2882\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15037\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__15042\,
            I => \N__15034\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__15037\,
            I => \N__15029\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15019\
        );

    \I__2878\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15016\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15032\,
            I => \N__15013\
        );

    \I__2876\ : Span4Mux_h
    port map (
            O => \N__15029\,
            I => \N__15010\
        );

    \I__2875\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15003\
        );

    \I__2874\ : InMux
    port map (
            O => \N__15027\,
            I => \N__15003\
        );

    \I__2873\ : InMux
    port map (
            O => \N__15026\,
            I => \N__15003\
        );

    \I__2872\ : InMux
    port map (
            O => \N__15025\,
            I => \N__14994\
        );

    \I__2871\ : InMux
    port map (
            O => \N__15024\,
            I => \N__14994\
        );

    \I__2870\ : InMux
    port map (
            O => \N__15023\,
            I => \N__14994\
        );

    \I__2869\ : InMux
    port map (
            O => \N__15022\,
            I => \N__14994\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__15019\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__15016\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__15013\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__15010\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__15003\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__14994\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__14981\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__14978\,
            I => \N__14975\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14972\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__14972\,
            I => \N__14969\
        );

    \I__2858\ : Span4Mux_h
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__14966\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__14963\,
            I => \Lab_UT.didp.countrce1.q_5_0_cascade_\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14957\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__14957\,
            I => \Lab_UT.three_2\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14951\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__14951\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_6\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__14948\,
            I => \N__14942\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__14947\,
            I => \N__14938\
        );

    \I__2849\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14935\
        );

    \I__2848\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14932\
        );

    \I__2847\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14929\
        );

    \I__2846\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14926\
        );

    \I__2845\ : InMux
    port map (
            O => \N__14938\,
            I => \N__14923\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14935\,
            I => \N__14920\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__14932\,
            I => \N__14917\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__14929\,
            I => \N__14913\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14926\,
            I => \N__14908\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__14923\,
            I => \N__14908\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__14920\,
            I => \N__14903\
        );

    \I__2838\ : Span4Mux_v
    port map (
            O => \N__14917\,
            I => \N__14903\
        );

    \I__2837\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14900\
        );

    \I__2836\ : Span4Mux_h
    port map (
            O => \N__14913\,
            I => \N__14897\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__14908\,
            I => \N__14894\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__14903\,
            I => \N__14891\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__14900\,
            I => \o_One_Sec_Pulse\
        );

    \I__2832\ : Odrv4
    port map (
            O => \N__14897\,
            I => \o_One_Sec_Pulse\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__14894\,
            I => \o_One_Sec_Pulse\
        );

    \I__2830\ : Odrv4
    port map (
            O => \N__14891\,
            I => \o_One_Sec_Pulse\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14878\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14875\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14872\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14875\,
            I => \N__14867\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__14872\,
            I => \N__14864\
        );

    \I__2824\ : InMux
    port map (
            O => \N__14871\,
            I => \N__14859\
        );

    \I__2823\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14859\
        );

    \I__2822\ : Span12Mux_s10_h
    port map (
            O => \N__14867\,
            I => \N__14856\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__14864\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14859\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2819\ : Odrv12
    port map (
            O => \N__14856\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2818\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__14846\,
            I => \N__14842\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14839\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__14842\,
            I => \N__14836\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__14839\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__14836\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2812\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14828\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14825\
        );

    \I__2810\ : Span4Mux_h
    port map (
            O => \N__14825\,
            I => \N__14822\
        );

    \I__2809\ : Odrv4
    port map (
            O => \N__14822\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__14819\,
            I => \uu2.N_97_cascade_\
        );

    \I__2807\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14810\
        );

    \I__2806\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14810\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__14810\,
            I => \uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14807\,
            I => \N__14804\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__14804\,
            I => \Lab_UT.dictrl.next_alarmstate_1\
        );

    \I__2802\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__14798\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14779\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14779\
        );

    \I__2798\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14779\
        );

    \I__2797\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14779\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14779\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__14790\,
            I => \N__14776\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__14779\,
            I => \N__14771\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14764\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14764\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14764\
        );

    \I__2790\ : Odrv4
    port map (
            O => \N__14771\,
            I => \Lab_UT.dictrl.un1_next_alarmstate21_0\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__14764\,
            I => \Lab_UT.dictrl.un1_next_alarmstate21_0\
        );

    \I__2788\ : InMux
    port map (
            O => \N__14759\,
            I => \N__14756\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__2786\ : Span4Mux_h
    port map (
            O => \N__14753\,
            I => \N__14748\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14752\,
            I => \N__14745\
        );

    \I__2784\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14742\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__14748\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__14745\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__14742\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__2779\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14729\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14729\,
            I => \N__14726\
        );

    \I__2777\ : Odrv12
    port map (
            O => \N__14726\,
            I => \Lab_UT.sec1Z0Z_1\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14719\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14715\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14719\,
            I => \N__14710\
        );

    \I__2773\ : IoInMux
    port map (
            O => \N__14718\,
            I => \N__14707\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__14715\,
            I => \N__14704\
        );

    \I__2771\ : InMux
    port map (
            O => \N__14714\,
            I => \N__14699\
        );

    \I__2770\ : InMux
    port map (
            O => \N__14713\,
            I => \N__14699\
        );

    \I__2769\ : Span4Mux_s3_v
    port map (
            O => \N__14710\,
            I => \N__14696\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__14707\,
            I => \N__14693\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__14704\,
            I => \N__14690\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14699\,
            I => \N__14687\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__14696\,
            I => \N__14682\
        );

    \I__2764\ : Span4Mux_s3_h
    port map (
            O => \N__14693\,
            I => \N__14682\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__14690\,
            I => rst
        );

    \I__2762\ : Odrv12
    port map (
            O => \N__14687\,
            I => rst
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__14682\,
            I => rst
        );

    \I__2760\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14671\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14668\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14665\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__14668\,
            I => \N__14662\
        );

    \I__2756\ : Odrv4
    port map (
            O => \N__14665\,
            I => \resetGen.un241_ci\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__14662\,
            I => \resetGen.un241_ci\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__14657\,
            I => \N__14654\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14642\
        );

    \I__2752\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14642\
        );

    \I__2751\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14642\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14642\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__14642\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__14639\,
            I => \N__14635\
        );

    \I__2747\ : InMux
    port map (
            O => \N__14638\,
            I => \N__14631\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14626\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14634\,
            I => \N__14626\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__14631\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__14626\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__14621\,
            I => \N__14616\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14613\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14610\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14616\,
            I => \N__14607\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__14613\,
            I => \N__14604\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__14610\,
            I => \N__14601\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14607\,
            I => \N__14594\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__14604\,
            I => \N__14594\
        );

    \I__2734\ : Span4Mux_v
    port map (
            O => \N__14601\,
            I => \N__14594\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__14594\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14582\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14582\
        );

    \I__2730\ : InMux
    port map (
            O => \N__14589\,
            I => \N__14582\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__14582\,
            I => \N__14576\
        );

    \I__2728\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14573\
        );

    \I__2727\ : InMux
    port map (
            O => \N__14580\,
            I => \N__14568\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14568\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__14576\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14573\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14568\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__14561\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__2721\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14549\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14549\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14549\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14549\,
            I => \N__14544\
        );

    \I__2717\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14541\
        );

    \I__2716\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14538\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__14544\,
            I => \N__14535\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__14541\,
            I => \N__14530\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__14538\,
            I => \N__14530\
        );

    \I__2712\ : Span4Mux_v
    port map (
            O => \N__14535\,
            I => \N__14527\
        );

    \I__2711\ : Span4Mux_v
    port map (
            O => \N__14530\,
            I => \N__14524\
        );

    \I__2710\ : Odrv4
    port map (
            O => \N__14527\,
            I => \resetGen.escKeyZ0\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__14524\,
            I => \resetGen.escKeyZ0\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14516\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14513\
        );

    \I__2706\ : Span4Mux_v
    port map (
            O => \N__14513\,
            I => \N__14509\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14512\,
            I => \N__14506\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__14509\,
            I => \N__14503\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14506\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__14503\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__14498\,
            I => \N__14493\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14497\,
            I => \N__14489\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14484\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14484\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14480\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__14489\,
            I => \N__14475\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__14484\,
            I => \N__14475\
        );

    \I__2694\ : InMux
    port map (
            O => \N__14483\,
            I => \N__14472\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14480\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__14475\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14472\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__14465\,
            I => \N__14461\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__14464\,
            I => \N__14456\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14451\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14451\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14446\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14456\,
            I => \N__14446\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__14451\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14446\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14441\,
            I => \N__14438\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__14438\,
            I => \uu2.vbuf_w_addr_user.un448_ci_0\
        );

    \I__2680\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__14432\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__14429\,
            I => \N__14426\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__14423\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_0\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__14420\,
            I => \N__14417\
        );

    \I__2674\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14414\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14411\,
            I => \N__14405\
        );

    \I__2671\ : InMux
    port map (
            O => \N__14410\,
            I => \N__14405\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__14405\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__14402\,
            I => \uu2.bitmap_pmux_sn_N_11_cascade_\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14396\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__14396\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14393\,
            I => \N__14390\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14390\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14381\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14374\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14374\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14374\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14381\,
            I => \N__14371\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14374\,
            I => \N__14363\
        );

    \I__2658\ : Span4Mux_v
    port map (
            O => \N__14371\,
            I => \N__14363\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14360\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14355\
        );

    \I__2655\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14355\
        );

    \I__2654\ : Odrv4
    port map (
            O => \N__14363\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14360\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14355\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__14348\,
            I => \N__14345\
        );

    \I__2650\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14342\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14336\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__14341\,
            I => \N__14333\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14329\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14326\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__14336\,
            I => \N__14323\
        );

    \I__2644\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14320\
        );

    \I__2643\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14317\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14329\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14326\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__14323\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__14320\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__14317\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2637\ : CascadeMux
    port map (
            O => \N__14306\,
            I => \N__14302\
        );

    \I__2636\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14298\
        );

    \I__2635\ : InMux
    port map (
            O => \N__14302\,
            I => \N__14295\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14301\,
            I => \N__14291\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14298\,
            I => \N__14287\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14295\,
            I => \N__14284\
        );

    \I__2631\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14280\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14291\,
            I => \N__14275\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14290\,
            I => \N__14275\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__14287\,
            I => \N__14272\
        );

    \I__2627\ : Span4Mux_h
    port map (
            O => \N__14284\,
            I => \N__14269\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14266\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__14280\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14275\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__2623\ : Odrv4
    port map (
            O => \N__14272\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__2622\ : Odrv4
    port map (
            O => \N__14269\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14266\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__14255\,
            I => \N__14252\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14249\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14245\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14241\
        );

    \I__2616\ : Span4Mux_h
    port map (
            O => \N__14245\,
            I => \N__14238\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__14244\,
            I => \N__14235\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__14241\,
            I => \N__14231\
        );

    \I__2613\ : Sp12to4
    port map (
            O => \N__14238\,
            I => \N__14228\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14223\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14223\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__14231\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2609\ : Odrv12
    port map (
            O => \N__14228\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__14223\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14213\,
            I => \N__14210\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14210\,
            I => \N__14204\
        );

    \I__2604\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14199\
        );

    \I__2603\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14199\
        );

    \I__2602\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14196\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__14204\,
            I => \N__14191\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__14199\,
            I => \N__14191\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14196\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__14191\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__2596\ : InMux
    port map (
            O => \N__14183\,
            I => \N__14178\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__14182\,
            I => \N__14174\
        );

    \I__2594\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14170\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14167\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__14177\,
            I => \N__14164\
        );

    \I__2591\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14159\
        );

    \I__2590\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14159\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14170\,
            I => \N__14154\
        );

    \I__2588\ : Span4Mux_h
    port map (
            O => \N__14167\,
            I => \N__14154\
        );

    \I__2587\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14151\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__14159\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__14154\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__14151\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__14144\,
            I => \uu2.un426_ci_3_cascade_\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2581\ : InMux
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__14135\,
            I => \N__14131\
        );

    \I__2579\ : InMux
    port map (
            O => \N__14134\,
            I => \N__14128\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__14131\,
            I => \uu2.un426_ci_3\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__14128\,
            I => \uu2.un426_ci_3\
        );

    \I__2576\ : InMux
    port map (
            O => \N__14123\,
            I => \N__14112\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14112\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14112\
        );

    \I__2573\ : InMux
    port map (
            O => \N__14120\,
            I => \N__14107\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14119\,
            I => \N__14107\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__14112\,
            I => \N__14104\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__2569\ : Span4Mux_h
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__14101\,
            I => \N__14095\
        );

    \I__2567\ : Odrv4
    port map (
            O => \N__14098\,
            I => \uu2.un404_ci\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__14095\,
            I => \uu2.un404_ci\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__14090\,
            I => \N__14087\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14082\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14079\
        );

    \I__2562\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14076\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__14082\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__14079\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__14076\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__2558\ : CEMux
    port map (
            O => \N__14069\,
            I => \N__14066\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__14066\,
            I => \N__14063\
        );

    \I__2556\ : Span4Mux_v
    port map (
            O => \N__14063\,
            I => \N__14060\
        );

    \I__2555\ : Span4Mux_s0_v
    port map (
            O => \N__14060\,
            I => \N__14057\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__14057\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2553\ : SRMux
    port map (
            O => \N__14054\,
            I => \N__14051\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__14051\,
            I => \N__14048\
        );

    \I__2551\ : Span4Mux_s1_v
    port map (
            O => \N__14048\,
            I => \N__14043\
        );

    \I__2550\ : SRMux
    port map (
            O => \N__14047\,
            I => \N__14040\
        );

    \I__2549\ : SRMux
    port map (
            O => \N__14046\,
            I => \N__14037\
        );

    \I__2548\ : Span4Mux_h
    port map (
            O => \N__14043\,
            I => \N__14032\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__14040\,
            I => \N__14032\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__14037\,
            I => \N__14029\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__14029\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__14026\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__14021\,
            I => \N__14018\
        );

    \I__2541\ : InMux
    port map (
            O => \N__14018\,
            I => \N__14015\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__14015\,
            I => \N__14012\
        );

    \I__2539\ : Span4Mux_s3_v
    port map (
            O => \N__14012\,
            I => \N__14009\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__14009\,
            I => \N__14006\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__14006\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__2536\ : CascadeMux
    port map (
            O => \N__14003\,
            I => \N__14000\
        );

    \I__2535\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13997\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__13997\,
            I => \N__13994\
        );

    \I__2533\ : Span4Mux_h
    port map (
            O => \N__13994\,
            I => \N__13991\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__13991\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__2531\ : InMux
    port map (
            O => \N__13988\,
            I => \N__13985\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__13985\,
            I => \uu2.mem0.bitmap_pmux_sn_N_42\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13979\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13979\,
            I => \N__13976\
        );

    \I__2527\ : Odrv4
    port map (
            O => \N__13976\,
            I => \uu2.un1_w_user_lf_0_0\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__13973\,
            I => \N__13970\
        );

    \I__2525\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13967\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13964\
        );

    \I__2523\ : Span4Mux_s1_v
    port map (
            O => \N__13964\,
            I => \N__13961\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__13961\,
            I => \N__13958\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__13958\,
            I => \uu2.un1_w_user_lfZ0Z_4\
        );

    \I__2520\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13952\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__13952\,
            I => \uu2.un20_w_addr_userZ0Z_1\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13943\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13943\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__13943\,
            I => \uu2.un3_w_addr_user\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__13940\,
            I => \uu2.un20_w_addr_userZ0Z_1_cascade_\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__13937\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2_cascade_\
        );

    \I__2513\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13921\
        );

    \I__2512\ : InMux
    port map (
            O => \N__13933\,
            I => \N__13921\
        );

    \I__2511\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13921\
        );

    \I__2510\ : InMux
    port map (
            O => \N__13931\,
            I => \N__13912\
        );

    \I__2509\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13912\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13912\
        );

    \I__2507\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13912\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__13921\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__13912\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13907\,
            I => \N__13904\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__13904\,
            I => \N__13901\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__13901\,
            I => \uu2.un3_w_addr_user_5\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13895\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__13895\,
            I => \N__13892\
        );

    \I__2499\ : Span4Mux_v
    port map (
            O => \N__13892\,
            I => \N__13889\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__13889\,
            I => bu_rx_data_fast_6
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \N__13883\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__13880\,
            I => bu_rx_data_fast_7
        );

    \I__2494\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13868\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13868\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13868\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__13868\,
            I => \N__13864\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13861\
        );

    \I__2489\ : Span4Mux_s3_v
    port map (
            O => \N__13864\,
            I => \N__13856\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__13861\,
            I => \N__13856\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__13856\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13853\,
            I => \N__13850\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13850\,
            I => \Lab_UT.dictrl.g2_1_0_0\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13847\,
            I => \N__13837\
        );

    \I__2483\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13837\
        );

    \I__2482\ : InMux
    port map (
            O => \N__13845\,
            I => \N__13828\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13844\,
            I => \N__13828\
        );

    \I__2480\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13828\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13828\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__13837\,
            I => \N__13823\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__13828\,
            I => \N__13823\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__13823\,
            I => \Lab_UT.nine\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__13820\,
            I => \N__13814\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13819\,
            I => \N__13809\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13809\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13806\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13803\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__13809\,
            I => \N__13796\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__13806\,
            I => \N__13796\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13803\,
            I => \N__13796\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__13796\,
            I => \Lab_UT.five\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__13793\,
            I => \N__13787\
        );

    \I__2465\ : InMux
    port map (
            O => \N__13792\,
            I => \N__13777\
        );

    \I__2464\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13777\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13777\
        );

    \I__2462\ : InMux
    port map (
            O => \N__13787\,
            I => \N__13777\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__13786\,
            I => \N__13773\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13777\,
            I => \N__13770\
        );

    \I__2459\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13765\
        );

    \I__2458\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13765\
        );

    \I__2457\ : Span4Mux_h
    port map (
            O => \N__13770\,
            I => \N__13759\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__2455\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13756\
        );

    \I__2454\ : Span4Mux_v
    port map (
            O => \N__13759\,
            I => \N__13753\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__13756\,
            I => \N__13750\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__2451\ : Span4Mux_v
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__13747\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__13744\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__2448\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13734\
        );

    \I__2447\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13729\
        );

    \I__2446\ : InMux
    port map (
            O => \N__13737\,
            I => \N__13729\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__13734\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13729\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__13724\,
            I => \N__13719\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13714\
        );

    \I__2441\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13714\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13710\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__13714\,
            I => \N__13707\
        );

    \I__2438\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13704\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13701\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__13707\,
            I => \N__13698\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13704\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__13701\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__13698\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13691\,
            I => \N__13686\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13690\,
            I => \N__13681\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13689\,
            I => \N__13681\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__13686\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__13681\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13673\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__13673\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__2425\ : InMux
    port map (
            O => \N__13670\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13663\
        );

    \I__2423\ : InMux
    port map (
            O => \N__13666\,
            I => \N__13660\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__13663\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__13660\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13655\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13652\,
            I => \N__13647\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13651\,
            I => \N__13642\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13650\,
            I => \N__13642\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13647\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__13642\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13637\,
            I => \N__13634\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__13634\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13631\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13624\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__13627\,
            I => \N__13620\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__13624\,
            I => \N__13616\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13623\,
            I => \N__13613\
        );

    \I__2407\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13608\
        );

    \I__2406\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13608\
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__13616\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__13613\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13608\,
            I => \buart.Z_rx.ser_clk\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13601\,
            I => \N__13595\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13590\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13590\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__13598\,
            I => \N__13582\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__13595\,
            I => \N__13577\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13574\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13571\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13568\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13587\,
            I => \N__13565\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13560\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13560\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13582\,
            I => \N__13553\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13581\,
            I => \N__13553\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13580\,
            I => \N__13553\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__13577\,
            I => \N__13550\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__13574\,
            I => \N__13547\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__13571\,
            I => \buart.Z_rx.startbit\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__13568\,
            I => \buart.Z_rx.startbit\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__13565\,
            I => \buart.Z_rx.startbit\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__13560\,
            I => \buart.Z_rx.startbit\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13553\,
            I => \buart.Z_rx.startbit\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__13550\,
            I => \buart.Z_rx.startbit\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__13547\,
            I => \buart.Z_rx.startbit\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13532\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__13529\,
            I => \N__13525\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__13528\,
            I => \N__13522\
        );

    \I__2376\ : InMux
    port map (
            O => \N__13525\,
            I => \N__13519\
        );

    \I__2375\ : InMux
    port map (
            O => \N__13522\,
            I => \N__13516\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__13519\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13516\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__13511\,
            I => \Lab_UT.dictrl.g2_0_1_0_cascade_\
        );

    \I__2371\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13505\,
            I => \Lab_UT.didp.countrce4.q_5_0\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13499\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13499\,
            I => \N__13494\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13491\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13488\
        );

    \I__2365\ : Span4Mux_v
    port map (
            O => \N__13494\,
            I => \N__13485\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13491\,
            I => \uu0_sec_clkD\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13488\,
            I => \uu0_sec_clkD\
        );

    \I__2362\ : Odrv4
    port map (
            O => \N__13485\,
            I => \uu0_sec_clkD\
        );

    \I__2361\ : CEMux
    port map (
            O => \N__13478\,
            I => \N__13475\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__13475\,
            I => \N__13472\
        );

    \I__2359\ : Sp12to4
    port map (
            O => \N__13472\,
            I => \N__13469\
        );

    \I__2358\ : Odrv12
    port map (
            O => \N__13469\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13460\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13465\,
            I => \N__13460\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13460\,
            I => \Lab_UT.didp.ce_11_0_2\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__13457\,
            I => \Lab_UT.didp.un26_ce_0_cascade_\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13443\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13443\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13438\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13438\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13433\
        );

    \I__2348\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13433\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13430\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13443\,
            I => \N__13427\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13438\,
            I => \N__13422\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13433\,
            I => \N__13422\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__13430\,
            I => \N__13419\
        );

    \I__2342\ : Span12Mux_s5_h
    port map (
            O => \N__13427\,
            I => \N__13416\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__13422\,
            I => \N__13413\
        );

    \I__2340\ : Odrv4
    port map (
            O => \N__13419\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__13416\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__13413\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__13406\,
            I => \Lab_UT.didp.ce_12_0_3_cascade_\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13400\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__13400\,
            I => \Lab_UT.didp.un26_ce_0\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13391\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13396\,
            I => \N__13391\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13391\,
            I => \N__13384\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13375\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13375\
        );

    \I__2329\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13375\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13387\,
            I => \N__13375\
        );

    \I__2327\ : Span4Mux_h
    port map (
            O => \N__13384\,
            I => \N__13372\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13375\,
            I => \N__13369\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__13372\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__13369\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__2322\ : InMux
    port map (
            O => \N__13361\,
            I => \N__13354\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13354\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13351\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__13354\,
            I => \N__13348\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__13351\,
            I => \N__13343\
        );

    \I__2317\ : Span4Mux_h
    port map (
            O => \N__13348\,
            I => \N__13343\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__13343\,
            I => \Lab_UT.nine_0\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__13340\,
            I => \N__13336\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13329\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13329\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__13335\,
            I => \N__13323\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__13334\,
            I => \N__13320\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__13329\,
            I => \N__13317\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13328\,
            I => \N__13312\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13312\
        );

    \I__2307\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13309\
        );

    \I__2306\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13306\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13303\
        );

    \I__2304\ : Span4Mux_h
    port map (
            O => \N__13317\,
            I => \N__13300\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13312\,
            I => \N__13297\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13290\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__13306\,
            I => \N__13290\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__13303\,
            I => \N__13290\
        );

    \I__2299\ : Odrv4
    port map (
            O => \N__13300\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__13297\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__2297\ : Odrv12
    port map (
            O => \N__13290\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__2295\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13265\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13265\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13278\,
            I => \N__13265\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13265\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13262\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13257\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13257\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__13265\,
            I => \N__13254\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13262\,
            I => \N__13249\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__13257\,
            I => \N__13249\
        );

    \I__2285\ : Sp12to4
    port map (
            O => \N__13254\,
            I => \N__13246\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__13249\,
            I => \N__13243\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__13246\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__13243\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__13238\,
            I => \Lab_UT.three_2_2_cascade_\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__13235\,
            I => \Lab_UT.didp.countrce4.q_5_2_cascade_\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \Lab_UT.didp.reset_12_3_3_cascade_\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__13229\,
            I => \Lab_UT.didp.reset_12_1_3_cascade_\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__13226\,
            I => \N__13222\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__13225\,
            I => \N__13217\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13222\,
            I => \N__13210\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13210\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13201\
        );

    \I__2272\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13201\
        );

    \I__2271\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13201\
        );

    \I__2270\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13201\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__13210\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__13201\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__13196\,
            I => \Lab_UT.didp.countrce4.un20_qPone_cascade_\
        );

    \I__2266\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13189\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13186\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__13189\,
            I => \Lab_UT.didp.countrce4.q_5_3\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__13186\,
            I => \Lab_UT.didp.countrce4.q_5_3\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__13181\,
            I => \N__13177\
        );

    \I__2261\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13174\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13177\,
            I => \N__13171\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__13174\,
            I => \N__13168\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__13171\,
            I => \N__13165\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__2256\ : Odrv12
    port map (
            O => \N__13165\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__13162\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13135\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13135\
        );

    \I__2252\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13135\
        );

    \I__2251\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13135\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13153\,
            I => \N__13135\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13152\,
            I => \N__13135\
        );

    \I__2248\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13135\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13150\,
            I => \N__13128\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__13135\,
            I => \N__13125\
        );

    \I__2245\ : InMux
    port map (
            O => \N__13134\,
            I => \N__13120\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13120\
        );

    \I__2243\ : InMux
    port map (
            O => \N__13132\,
            I => \N__13115\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13115\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13128\,
            I => \N__13110\
        );

    \I__2240\ : Span4Mux_h
    port map (
            O => \N__13125\,
            I => \N__13110\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__13120\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__13115\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__13110\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__13103\,
            I => \N__13097\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__13102\,
            I => \N__13094\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__13101\,
            I => \N__13090\
        );

    \I__2233\ : CascadeMux
    port map (
            O => \N__13100\,
            I => \N__13086\
        );

    \I__2232\ : InMux
    port map (
            O => \N__13097\,
            I => \N__13069\
        );

    \I__2231\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13069\
        );

    \I__2230\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13069\
        );

    \I__2229\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13069\
        );

    \I__2228\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13069\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13086\,
            I => \N__13069\
        );

    \I__2226\ : InMux
    port map (
            O => \N__13085\,
            I => \N__13069\
        );

    \I__2225\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13065\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__13069\,
            I => \N__13058\
        );

    \I__2223\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13055\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__13065\,
            I => \N__13052\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13049\
        );

    \I__2220\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13046\
        );

    \I__2219\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13041\
        );

    \I__2218\ : InMux
    port map (
            O => \N__13061\,
            I => \N__13041\
        );

    \I__2217\ : Span4Mux_h
    port map (
            O => \N__13058\,
            I => \N__13038\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13055\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2215\ : Odrv12
    port map (
            O => \N__13052\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__13049\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__13046\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__13041\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__13038\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__13025\,
            I => \N__13019\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__13024\,
            I => \N__13014\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__13023\,
            I => \N__13010\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__13022\,
            I => \N__13006\
        );

    \I__2206\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13001\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13018\,
            I => \N__12986\
        );

    \I__2204\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12986\
        );

    \I__2203\ : InMux
    port map (
            O => \N__13014\,
            I => \N__12986\
        );

    \I__2202\ : InMux
    port map (
            O => \N__13013\,
            I => \N__12986\
        );

    \I__2201\ : InMux
    port map (
            O => \N__13010\,
            I => \N__12986\
        );

    \I__2200\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12986\
        );

    \I__2199\ : InMux
    port map (
            O => \N__13006\,
            I => \N__12986\
        );

    \I__2198\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12981\
        );

    \I__2197\ : InMux
    port map (
            O => \N__13004\,
            I => \N__12981\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__13001\,
            I => \N__12976\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12986\,
            I => \N__12976\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__12981\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__12976\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12960\
        );

    \I__2191\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12954\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12939\
        );

    \I__2189\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12939\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12939\
        );

    \I__2187\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12939\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12939\
        );

    \I__2185\ : InMux
    port map (
            O => \N__12964\,
            I => \N__12939\
        );

    \I__2184\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12939\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12936\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12933\
        );

    \I__2181\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12928\
        );

    \I__2180\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12928\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__12954\,
            I => \N__12923\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__12939\,
            I => \N__12923\
        );

    \I__2177\ : Span4Mux_h
    port map (
            O => \N__12936\,
            I => \N__12920\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12933\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__12928\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__12923\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__12920\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__2172\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12908\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__12908\,
            I => \Lab_UT.didp.countrce3.q_5_3\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__12905\,
            I => \N__12901\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__12904\,
            I => \N__12898\
        );

    \I__2168\ : InMux
    port map (
            O => \N__12901\,
            I => \N__12895\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12898\,
            I => \N__12892\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12895\,
            I => \Lab_UT.didp.q_fast_1\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__12892\,
            I => \Lab_UT.didp.q_fast_1\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12884\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12884\,
            I => \Lab_UT.didp.countrce4.q_5_1\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__12881\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__2161\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__12875\,
            I => \N__12871\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__12874\,
            I => \N__12868\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__12871\,
            I => \N__12864\
        );

    \I__2157\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12859\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12859\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__12864\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_0\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__12859\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_0\
        );

    \I__2153\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12845\
        );

    \I__2152\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12845\
        );

    \I__2151\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12840\
        );

    \I__2150\ : InMux
    port map (
            O => \N__12851\,
            I => \N__12840\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12837\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12845\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__12840\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12837\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__12830\,
            I => \N__12824\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12816\
        );

    \I__2143\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12816\
        );

    \I__2142\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12816\
        );

    \I__2141\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12811\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12811\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__12816\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__12811\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0\
        );

    \I__2137\ : InMux
    port map (
            O => \N__12806\,
            I => \N__12795\
        );

    \I__2136\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12795\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12795\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12803\,
            I => \N__12790\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12802\,
            I => \N__12790\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__12795\,
            I => \Lab_UT.dictrl.next_alarmstate_1_1\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__12790\,
            I => \Lab_UT.dictrl.next_alarmstate_1_1\
        );

    \I__2130\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12782\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__12782\,
            I => \N__12778\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__12781\,
            I => \N__12774\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__12778\,
            I => \N__12770\
        );

    \I__2126\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12767\
        );

    \I__2125\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12762\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12762\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__12770\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__12767\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__12762\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__2120\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12749\
        );

    \I__2119\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12749\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__12746\,
            I => \N__12739\
        );

    \I__2116\ : InMux
    port map (
            O => \N__12745\,
            I => \N__12736\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12729\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12729\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12742\,
            I => \N__12729\
        );

    \I__2112\ : Odrv4
    port map (
            O => \N__12739\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12736\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__12729\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__2109\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12719\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__12719\,
            I => \Lab_UT.alarmchar_2_1_1\
        );

    \I__2107\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12713\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12708\
        );

    \I__2105\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12705\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12702\
        );

    \I__2103\ : Odrv4
    port map (
            O => \N__12708\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12705\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__12702\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__2100\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12689\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12689\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__12689\,
            I => \Lab_UT.didp.countrce2.q_5_1\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__12686\,
            I => \N__12683\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12680\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__12680\,
            I => \Lab_UT.didp.countrce2.q_5_2\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12674\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__2092\ : IoInMux
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__12668\,
            I => \N__12665\
        );

    \I__2090\ : IoSpan4Mux
    port map (
            O => \N__12665\,
            I => \N__12661\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__12664\,
            I => \N__12658\
        );

    \I__2088\ : Span4Mux_s0_v
    port map (
            O => \N__12661\,
            I => \N__12652\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__12658\,
            I => \N__12652\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12649\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__12652\,
            I => \N__12645\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__12649\,
            I => \N__12642\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12648\,
            I => \N__12639\
        );

    \I__2082\ : Span4Mux_v
    port map (
            O => \N__12645\,
            I => \N__12636\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__12642\,
            I => \N__12633\
        );

    \I__2080\ : InMux
    port map (
            O => \N__12639\,
            I => \N__12630\
        );

    \I__2079\ : Odrv4
    port map (
            O => \N__12636\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__12633\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__12630\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2076\ : CEMux
    port map (
            O => \N__12623\,
            I => \N__12620\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12617\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__12617\,
            I => \Lab_UT.dictrl.G_64\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12608\
        );

    \I__2072\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12608\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__12608\,
            I => \Lab_UT.alarmMatch\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__12605\,
            I => \Lab_UT.dictrl.idle_cascade_\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__12602\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\
        );

    \I__2068\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12596\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__12596\,
            I => \Lab_UT.alarmchar9\
        );

    \I__2066\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12590\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__12587\,
            I => \Lab_UT.alarmchar10\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12578\
        );

    \I__2061\ : Span4Mux_h
    port map (
            O => \N__12578\,
            I => \N__12575\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__12575\,
            I => \Lab_UT.alarmchar10_i_2\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__12572\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__12569\,
            I => \uu2.N_57_cascade_\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12563\,
            I => \N__12557\
        );

    \I__2055\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12557\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__12557\,
            I => \N__12553\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12556\,
            I => \N__12550\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__12553\,
            I => \uu2.w_data_i_a3_0_5\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12550\,
            I => \uu2.w_data_i_a3_0_5\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12545\,
            I => \uu2.mem0.w_data_0_a3_0_6_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__2046\ : Span4Mux_s3_h
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__12530\,
            I => \uu2.mem0.w_data_6\
        );

    \I__2044\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12522\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12517\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12517\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12522\,
            I => \uu2.w_data_displaying_2_i_a2_i_a2_0_0\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__12517\,
            I => \uu2.w_data_displaying_2_i_a2_i_a2_0_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2037\ : Odrv12
    port map (
            O => \N__12506\,
            I => \Lab_UT.alarmcharZ0Z_4\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__12503\,
            I => \N__12498\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12495\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12492\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12489\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12495\,
            I => \L3_tx_data_6\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12492\,
            I => \L3_tx_data_6\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12489\,
            I => \L3_tx_data_6\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12477\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12472\
        );

    \I__2027\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12472\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__12477\,
            I => \L3_tx_data_3\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__12472\,
            I => \L3_tx_data_3\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12464\,
            I => \N__12459\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12456\
        );

    \I__2021\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12453\
        );

    \I__2020\ : Odrv4
    port map (
            O => \N__12459\,
            I => \L3_tx_data_0\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__12456\,
            I => \L3_tx_data_0\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12453\,
            I => \L3_tx_data_0\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12443\,
            I => \uu2.un1_w_user_crZ0Z_4\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__12440\,
            I => \uu2_un1_w_user_cr_0_cascade_\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__12437\,
            I => \N__12433\
        );

    \I__2013\ : CascadeMux
    port map (
            O => \N__12436\,
            I => \N__12429\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12426\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12421\
        );

    \I__2010\ : InMux
    port map (
            O => \N__12429\,
            I => \N__12421\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__12426\,
            I => \L3_tx_data_2\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__12421\,
            I => \L3_tx_data_2\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12413\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12410\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__12407\,
            I => \uu2.mem0.w_data_2\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__12401\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_44\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__12398\,
            I => \N__12395\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12392\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12389\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__12389\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__12386\,
            I => \uu2.mem0.bitmap_pmux_sn_N_33_cascade_\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12383\,
            I => \N__12380\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12380\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__12377\,
            I => \N__12373\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__12376\,
            I => \N__12370\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12367\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12364\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12367\,
            I => \uu2.N_34\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__12364\,
            I => \uu2.N_34\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12356\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__12356\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_42\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12347\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12347\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12347\,
            I => \N__12344\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__12344\,
            I => \uu2.N_49\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__12341\,
            I => \N__12337\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__1980\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__12334\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12331\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12326\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12323\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12320\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__1974\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12308\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12308\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12308\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12308\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1970\ : InMux
    port map (
            O => \N__12305\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12302\,
            I => \N__12299\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12299\,
            I => \uu2.un3_w_addr_user_4\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12296\,
            I => \N__12290\
        );

    \I__1966\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12290\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__12290\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12281\
        );

    \I__1963\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12281\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__12281\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__12278\,
            I => \N__12274\
        );

    \I__1960\ : InMux
    port map (
            O => \N__12277\,
            I => \N__12269\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12269\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__12269\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1957\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12260\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12260\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12260\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12254\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__12254\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__12251\,
            I => \N__12248\
        );

    \I__1951\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__12245\,
            I => \N__12242\
        );

    \I__1949\ : Span4Mux_s3_h
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__12239\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__12236\,
            I => \N__12233\
        );

    \I__1946\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12227\
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__12227\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__12224\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__1942\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12218\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__12218\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__12215\,
            I => \buart.Z_rx.ser_clk_cascade_\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12209\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__12209\,
            I => \N__12202\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12199\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12194\
        );

    \I__1935\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12194\
        );

    \I__1934\ : InMux
    port map (
            O => \N__12205\,
            I => \N__12191\
        );

    \I__1933\ : Span4Mux_v
    port map (
            O => \N__12202\,
            I => \N__12188\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__12199\,
            I => \N__12183\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__12194\,
            I => \N__12183\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__12191\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__12188\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1928\ : Odrv12
    port map (
            O => \N__12183\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__1927\ : IoInMux
    port map (
            O => \N__12176\,
            I => \N__12173\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__12173\,
            I => \N__12170\
        );

    \I__1925\ : Span4Mux_s3_v
    port map (
            O => \N__12170\,
            I => \N__12167\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__12167\,
            I => \buart.Z_rx.sample\
        );

    \I__1923\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12160\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__12157\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1919\ : Odrv12
    port map (
            O => \N__12154\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1918\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12143\
        );

    \I__1917\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12143\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__12143\,
            I => \buart.Z_rx.idle\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__12140\,
            I => \buart.Z_rx.startbit_cascade_\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12132\
        );

    \I__1913\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12129\
        );

    \I__1912\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12126\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__12132\,
            I => bu_rx_data_rdy
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__12129\,
            I => bu_rx_data_rdy
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__12126\,
            I => bu_rx_data_rdy
        );

    \I__1908\ : CEMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__12116\,
            I => \N__12111\
        );

    \I__1906\ : CEMux
    port map (
            O => \N__12115\,
            I => \N__12108\
        );

    \I__1905\ : CEMux
    port map (
            O => \N__12114\,
            I => \N__12105\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__12111\,
            I => \N__12100\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__12108\,
            I => \N__12100\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__12105\,
            I => \N__12097\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__12100\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__12097\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__12092\,
            I => \N__12086\
        );

    \I__1898\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12086\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__1896\ : Span4Mux_v
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__12080\,
            I => \Lab_UT.didp.countrce2.q_5_0\
        );

    \I__1894\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12071\
        );

    \I__1893\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12064\
        );

    \I__1892\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12064\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12064\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12071\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12064\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1888\ : CascadeMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12051\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12046\
        );

    \I__1885\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12046\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__12051\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__12046\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1882\ : InMux
    port map (
            O => \N__12041\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__12038\,
            I => \Lab_UT.dicLdAMones_0_cascade_\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12035\,
            I => \N__12032\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__12032\,
            I => \N__12028\
        );

    \I__1878\ : InMux
    port map (
            O => \N__12031\,
            I => \N__12024\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__12028\,
            I => \N__12021\
        );

    \I__1876\ : InMux
    port map (
            O => \N__12027\,
            I => \N__12018\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__12024\,
            I => \N__12015\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__12021\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__12018\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__12015\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12008\,
            I => \N__12005\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__12005\,
            I => \N__12000\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11997\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11994\
        );

    \I__1867\ : Span4Mux_v
    port map (
            O => \N__12000\,
            I => \N__11989\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11989\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__11994\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__11989\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__1863\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11976\
        );

    \I__1861\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11973\
        );

    \I__1860\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11970\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__11976\,
            I => \N__11965\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11965\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__11970\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__11965\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__11960\,
            I => \N__11956\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11948\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11948\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11948\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11948\,
            I => \Lab_UT.dicLdAMones_0\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__11945\,
            I => \N__11940\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11937\
        );

    \I__1848\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11934\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11931\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__11937\,
            I => \N__11926\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11934\,
            I => \N__11926\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__11931\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__11926\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__1842\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__1839\ : Odrv4
    port map (
            O => \N__11912\,
            I => \resetGen.escKeyZ0Z_5\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__11909\,
            I => \resetGen.escKeyZ0Z_4_cascade_\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__11906\,
            I => \Lab_UT.didp.countrce3.q_5_3_cascade_\
        );

    \I__1836\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11897\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11897\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__11897\,
            I => \Lab_UT.didp.countrce3.q_fastZ0Z_3\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__11894\,
            I => \N__11890\
        );

    \I__1832\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11885\
        );

    \I__1831\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11885\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11885\,
            I => \Lab_UT.didp.q_fast_3\
        );

    \I__1829\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11879\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__11879\,
            I => \Lab_UT.didp.countrce3.did_alarmMatch_0\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11872\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11869\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__11872\,
            I => \N__11866\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11869\,
            I => \N__11863\
        );

    \I__1823\ : Odrv12
    port map (
            O => \N__11866\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__11863\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__1821\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11854\
        );

    \I__1820\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11851\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__11854\,
            I => \N__11848\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11851\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__11848\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__1816\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11837\
        );

    \I__1815\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11837\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__1813\ : Odrv12
    port map (
            O => \N__11834\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11831\,
            I => \N__11828\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__11828\,
            I => \N__11824\
        );

    \I__1810\ : InMux
    port map (
            O => \N__11827\,
            I => \N__11821\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__11824\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__11821\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__11816\,
            I => \Lab_UT.three_2_0_cascade_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11813\,
            I => \N__11809\
        );

    \I__1805\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11806\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__11809\,
            I => \N__11803\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__11806\,
            I => \N__11800\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__11803\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__11800\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11792\,
            I => \Lab_UT.didp.did_alarmMatch_3\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11782\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11785\,
            I => \N__11779\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__11782\,
            I => \Lab_UT.didp.countrce2.q_fastZ0Z_1\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__11779\,
            I => \Lab_UT.didp.countrce2.q_fastZ0Z_1\
        );

    \I__1793\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11770\
        );

    \I__1792\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11767\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__11770\,
            I => \Lab_UT.didp.countrce3.q_fastZ0Z_1\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__11767\,
            I => \Lab_UT.didp.countrce3.q_fastZ0Z_1\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__11762\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \N__11756\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11752\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11748\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11752\,
            I => \N__11745\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11742\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__11748\,
            I => \N__11739\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__11745\,
            I => \Lab_UT.didp.q_fast_0\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__11742\,
            I => \Lab_UT.didp.q_fast_0\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__11739\,
            I => \Lab_UT.didp.q_fast_0\
        );

    \I__1779\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__11729\,
            I => \N__11726\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__11726\,
            I => \Lab_UT.didp.countrce2.un20_qPone\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__11723\,
            I => \Lab_UT.didp.countrce2.q_5_3_cascade_\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11717\,
            I => \N__11712\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11709\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11706\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__11712\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11709\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11706\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__1768\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11696\,
            I => \N__11692\
        );

    \I__1766\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11689\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__11692\,
            I => \Lab_UT.didp.countrce2.q_fastZ0Z_3\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__11689\,
            I => \Lab_UT.didp.countrce2.q_fastZ0Z_3\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11680\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11677\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11680\,
            I => \N__11674\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11671\
        );

    \I__1759\ : Span4Mux_v
    port map (
            O => \N__11674\,
            I => \N__11668\
        );

    \I__1758\ : Span4Mux_h
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__11668\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__1756\ : Odrv4
    port map (
            O => \N__11665\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__1755\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11657\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__11657\,
            I => \Lab_UT.didp.countrce2.q_5_3\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__11651\,
            I => \Lab_UT.didp.did_alarmMatch_2\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__11648\,
            I => \Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_\
        );

    \I__1750\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__11642\,
            I => \Lab_UT.didp.did_alarmMatch_12\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__11636\,
            I => \Lab_UT.min1Z0Z_0\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__11630\,
            I => \N__11627\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__11627\,
            I => \Lab_UT.dispString.m25_ns_1\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11618\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11618\,
            I => \Lab_UT.min1Z0Z_2\
        );

    \I__1740\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__11612\,
            I => \N__11609\
        );

    \I__1738\ : Odrv12
    port map (
            O => \N__11609\,
            I => \Lab_UT.dispString.N_65\
        );

    \I__1737\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11603\,
            I => \Lab_UT.alarmcharZ0Z_6\
        );

    \I__1735\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11597\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__11597\,
            I => \N__11579\
        );

    \I__1733\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11574\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11574\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11594\,
            I => \N__11571\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11564\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11592\,
            I => \N__11564\
        );

    \I__1728\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11564\
        );

    \I__1727\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11555\
        );

    \I__1726\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11555\
        );

    \I__1725\ : InMux
    port map (
            O => \N__11588\,
            I => \N__11555\
        );

    \I__1724\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11555\
        );

    \I__1723\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11548\
        );

    \I__1722\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11548\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11548\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11544\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11582\,
            I => \N__11541\
        );

    \I__1718\ : Span4Mux_h
    port map (
            O => \N__11579\,
            I => \N__11536\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__11574\,
            I => \N__11536\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__11571\,
            I => \N__11527\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11564\,
            I => \N__11527\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__11555\,
            I => \N__11527\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11548\,
            I => \N__11527\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11524\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11544\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__11541\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__11536\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__1708\ : Odrv12
    port map (
            O => \N__11527\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__11524\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__11510\,
            I => \Lab_UT.alarmcharZ0Z_2\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__11495\,
            I => \Lab_UT.sec2Z0Z_2\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__11492\,
            I => \N__11486\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__11491\,
            I => \N__11483\
        );

    \I__1697\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11465\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11465\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11460\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11460\
        );

    \I__1693\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11457\
        );

    \I__1692\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11450\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11450\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11479\,
            I => \N__11450\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11478\,
            I => \N__11443\
        );

    \I__1688\ : InMux
    port map (
            O => \N__11477\,
            I => \N__11443\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11443\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11438\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11431\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11431\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11431\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11426\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11470\,
            I => \N__11426\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11465\,
            I => \N__11423\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__11460\,
            I => \N__11418\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11457\,
            I => \N__11418\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11450\,
            I => \N__11415\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11443\,
            I => \N__11412\
        );

    \I__1675\ : InMux
    port map (
            O => \N__11442\,
            I => \N__11407\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11407\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11438\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11431\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11426\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__11423\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1669\ : Odrv4
    port map (
            O => \N__11418\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__11415\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__11412\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__11407\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11387\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__11387\,
            I => \Lab_UT.dispString.N_68\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11381\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_5\
        );

    \I__1661\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__11375\,
            I => \N__11372\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__11372\,
            I => \Lab_UT.didp.did_alarmMatch_11\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__11369\,
            I => \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__11366\,
            I => \Lab_UT.dispString.N_86_cascade_\
        );

    \I__1656\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__11357\,
            I => \Lab_UT.dispString.N_89\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11351\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11351\,
            I => \Lab_UT.min2Z0Z_0\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11345\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11345\,
            I => \Lab_UT.dispString.m49_ns_1\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__11336\,
            I => \Lab_UT.sec1Z0Z_0\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__11333\,
            I => \N__11322\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__11332\,
            I => \N__11318\
        );

    \I__1644\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11315\
        );

    \I__1643\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11308\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11308\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11308\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11327\,
            I => \N__11305\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11300\
        );

    \I__1638\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11300\
        );

    \I__1637\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11297\
        );

    \I__1636\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11292\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11292\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__11315\,
            I => \N__11287\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11287\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11305\,
            I => \N__11282\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__11300\,
            I => \N__11282\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__11297\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11292\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__11287\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__11282\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__11270\,
            I => \N__11265\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11269\,
            I => \N__11262\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11268\,
            I => \N__11259\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__11265\,
            I => \L3_tx_data_5\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__11262\,
            I => \L3_tx_data_5\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11259\,
            I => \L3_tx_data_5\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11246\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11241\
        );

    \I__1616\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11238\
        );

    \I__1615\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11235\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__11241\,
            I => \L3_tx_data_4\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__11238\,
            I => \L3_tx_data_4\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11235\,
            I => \L3_tx_data_4\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__11228\,
            I => \N__11224\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11221\
        );

    \I__1609\ : InMux
    port map (
            O => \N__11224\,
            I => \N__11218\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__11218\,
            I => \N__11212\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__11215\,
            I => \Lab_UT.alarmcharZ0Z_1\
        );

    \I__1605\ : Odrv4
    port map (
            O => \N__11212\,
            I => \Lab_UT.alarmcharZ0Z_1\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__1601\ : Span4Mux_v
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__11195\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__1599\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__11189\,
            I => \Lab_UT.dispString.m40_ns_1\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__11186\,
            I => \N__11183\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__11180\,
            I => \Lab_UT.min1Z0Z_3\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__11177\,
            I => \Lab_UT.dispString.N_77_cascade_\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11171\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11171\,
            I => \Lab_UT.dispString.N_80\
        );

    \I__1591\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__11165\,
            I => \Lab_UT.sec2Z0Z_3\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__11162\,
            I => \uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_\
        );

    \I__1588\ : InMux
    port map (
            O => \N__11159\,
            I => \N__11156\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__11156\,
            I => \uu2.mem0.w_data_0_1_3\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__1585\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11147\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__1583\ : Odrv12
    port map (
            O => \N__11144\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__1582\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__11138\,
            I => \uu2.mem0.bitmap_pmux_sn_N_33_0\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__11135\,
            I => \uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__11132\,
            I => \uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_\
        );

    \I__1578\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__11126\,
            I => \uu2.mem0.N_409\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__11123\,
            I => \uu2.N_34_cascade_\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11113\
        );

    \I__1573\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__11113\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__11110\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \buart.Z_tx.ser_clk_cascade_\
        );

    \I__1569\ : InMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__11099\,
            I => \buart.Z_tx.uart_busy_0_0\
        );

    \I__1567\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11093\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__11093\,
            I => \N__11087\
        );

    \I__1565\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11084\
        );

    \I__1564\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11078\
        );

    \I__1563\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11078\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__11087\,
            I => \N__11073\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__11084\,
            I => \N__11073\
        );

    \I__1560\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11070\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__11078\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__11073\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__11070\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__11063\,
            I => \N__11059\
        );

    \I__1555\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11051\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11051\
        );

    \I__1553\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11051\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__11051\,
            I => \N__11047\
        );

    \I__1551\ : InMux
    port map (
            O => \N__11050\,
            I => \N__11044\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__11047\,
            I => \N__11041\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__11044\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__11041\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1547\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11032\
        );

    \I__1546\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11026\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__11032\,
            I => \N__11023\
        );

    \I__1544\ : InMux
    port map (
            O => \N__11031\,
            I => \N__11020\
        );

    \I__1543\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11015\
        );

    \I__1542\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11015\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__11026\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__11023\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11020\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__11015\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__11006\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__1536\ : InMux
    port map (
            O => \N__11003\,
            I => \N__10994\
        );

    \I__1535\ : InMux
    port map (
            O => \N__11002\,
            I => \N__10994\
        );

    \I__1534\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10994\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__10994\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1532\ : InMux
    port map (
            O => \N__10991\,
            I => \N__10988\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__10988\,
            I => \buart.Z_tx.un1_bitcount_c3\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10979\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__10976\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__1526\ : IoInMux
    port map (
            O => \N__10973\,
            I => \N__10970\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10966\
        );

    \I__1524\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10963\
        );

    \I__1523\ : Span12Mux_s9_v
    port map (
            O => \N__10966\,
            I => \N__10960\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__10960\,
            I => clk
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__10957\,
            I => clk
        );

    \I__1519\ : CEMux
    port map (
            O => \N__10952\,
            I => \N__10949\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10945\
        );

    \I__1517\ : SRMux
    port map (
            O => \N__10948\,
            I => \N__10942\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__10945\,
            I => \N__10939\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__10942\,
            I => \N__10934\
        );

    \I__1514\ : Span4Mux_s1_h
    port map (
            O => \N__10939\,
            I => \N__10934\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__10934\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__1511\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1509\ : Odrv4
    port map (
            O => \N__10922\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10912\
        );

    \I__1507\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10903\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10917\,
            I => \N__10903\
        );

    \I__1505\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10903\
        );

    \I__1504\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10903\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__10912\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__10903\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10895\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10892\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10882\
        );

    \I__1497\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10879\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10874\
        );

    \I__1495\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10874\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10871\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10882\,
            I => \N__10864\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__10879\,
            I => \N__10864\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10864\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10871\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1489\ : Odrv12
    port map (
            O => \N__10864\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__1487\ : InMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__1485\ : Odrv12
    port map (
            O => \N__10850\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10847\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__10844\,
            I => \N__10838\
        );

    \I__1482\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10834\
        );

    \I__1481\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10825\
        );

    \I__1480\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10825\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10825\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10825\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10834\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10825\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__10820\,
            I => \N__10817\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__10814\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10811\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10802\
        );

    \I__1470\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10802\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__10802\,
            I => \N__10799\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__10799\,
            I => \N__10794\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10791\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10788\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__10794\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__10791\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10788\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10781\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10769\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10774\,
            I => \N__10762\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10762\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10762\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10769\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__10762\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1454\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__10754\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10747\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10750\,
            I => \N__10744\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10747\,
            I => \N__10741\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__10744\,
            I => \N__10738\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__10741\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__10738\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__1446\ : CEMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1443\ : Span4Mux_s0_h
    port map (
            O => \N__10724\,
            I => \N__10720\
        );

    \I__1442\ : CEMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__10720\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__10717\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__10712\,
            I => \buart.Z_rx.valid_0_cascade_\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__10709\,
            I => \buart.Z_rx.idle_0_cascade_\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__10706\,
            I => \buart.Z_rx.idle_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__10703\,
            I => \buart.Z_rx.N_27_0_i_cascade_\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__10700\,
            I => \Lab_UT.three_2_1_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10694\,
            I => \Lab_UT.didp.countrce3.q_5_2\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__10691\,
            I => \Lab_UT.didp.countrce3.q_5_2_cascade_\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__10688\,
            I => \N__10684\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10681\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10678\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__10681\,
            I => \Lab_UT.didp.countrce3.q_fastZ0Z_2\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__10678\,
            I => \Lab_UT.didp.countrce3.q_fastZ0Z_2\
        );

    \I__1426\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10668\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10665\
        );

    \I__1424\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10662\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__10668\,
            I => \N__10659\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10665\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__10662\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__10659\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10652\,
            I => \Lab_UT.didp.did_alarmMatch_6_cascade_\
        );

    \I__1418\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1415\ : Odrv4
    port map (
            O => \N__10640\,
            I => \Lab_UT.min2Z0Z_3\
        );

    \I__1414\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10634\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1412\ : Odrv12
    port map (
            O => \N__10631\,
            I => \Lab_UT.min1Z0Z_1\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10624\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10621\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10624\,
            I => \N__10618\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__10621\,
            I => \N__10615\
        );

    \I__1407\ : Span4Mux_h
    port map (
            O => \N__10618\,
            I => \N__10612\
        );

    \I__1406\ : Odrv4
    port map (
            O => \N__10615\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__10612\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__1404\ : CascadeMux
    port map (
            O => \N__10607\,
            I => \N__10602\
        );

    \I__1403\ : InMux
    port map (
            O => \N__10606\,
            I => \N__10589\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10605\,
            I => \N__10589\
        );

    \I__1401\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10586\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10571\
        );

    \I__1399\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10571\
        );

    \I__1398\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10571\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10571\
        );

    \I__1396\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10571\
        );

    \I__1395\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10571\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10571\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10564\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__10589\,
            I => \N__10561\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10558\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__10571\,
            I => \N__10555\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10548\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10548\
        );

    \I__1387\ : InMux
    port map (
            O => \N__10568\,
            I => \N__10548\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10545\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__10564\,
            I => \N__10539\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__10561\,
            I => \N__10539\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__10558\,
            I => \N__10534\
        );

    \I__1382\ : Span4Mux_s3_h
    port map (
            O => \N__10555\,
            I => \N__10534\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10531\
        );

    \I__1380\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10526\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10526\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__10539\,
            I => vbuf_tx_data_rdy
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__10534\,
            I => vbuf_tx_data_rdy
        );

    \I__1376\ : Odrv4
    port map (
            O => \N__10531\,
            I => vbuf_tx_data_rdy
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10526\,
            I => vbuf_tx_data_rdy
        );

    \I__1374\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10510\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__1371\ : Span4Mux_h
    port map (
            O => \N__10510\,
            I => \N__10502\
        );

    \I__1370\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10495\
        );

    \I__1369\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10495\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10495\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__10502\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10495\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10486\
        );

    \I__1364\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10481\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10476\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10471\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10471\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10468\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10463\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10479\,
            I => \N__10463\
        );

    \I__1357\ : Span4Mux_s1_h
    port map (
            O => \N__10476\,
            I => \N__10460\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10471\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__10468\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__10463\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__10460\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10446\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10441\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10449\,
            I => \N__10438\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10446\,
            I => \N__10435\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10445\,
            I => \N__10430\
        );

    \I__1347\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10430\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10441\,
            I => \N__10427\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__10438\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__10435\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__10430\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__10427\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1341\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__10412\,
            I => \uu0.un143_ci_0\
        );

    \I__1338\ : CEMux
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10402\
        );

    \I__1336\ : CEMux
    port map (
            O => \N__10405\,
            I => \N__10399\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__10402\,
            I => \N__10394\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__10399\,
            I => \N__10394\
        );

    \I__1333\ : Span4Mux_v
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__1332\ : Span4Mux_s2_h
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__10388\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__1327\ : Odrv12
    port map (
            O => \N__10376\,
            I => \resetGen.reset_count_2_0_4\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10370\,
            I => \Lab_UT.dispString.N_46\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1323\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10361\,
            I => \Lab_UT.min2Z0Z_1\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10355\,
            I => \Lab_UT.min2Z0Z_2\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__10346\,
            I => \Lab_UT.sec1Z0Z_2\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \Lab_UT.dicLdAStens_0_cascade_\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__10337\,
            I => \Lab_UT.alarmcharZ0Z_5\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \Lab_UT.dispString.m35_ns_1_cascade_\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__10328\,
            I => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__10319\,
            I => \Lab_UT.sec2Z0Z_0\
        );

    \I__1307\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10313\,
            I => \Lab_UT.alarmcharZ0Z_0\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10310\,
            I => \Lab_UT.dispString.m32_ns_1_cascade_\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1303\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__10301\,
            I => \Lab_UT.sec1Z0Z_3\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \N__10295\
        );

    \I__1300\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10292\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__10292\,
            I => \Lab_UT.sec2Z0Z_1\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__10289\,
            I => \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\
        );

    \I__1297\ : CEMux
    port map (
            O => \N__10286\,
            I => \N__10281\
        );

    \I__1296\ : CEMux
    port map (
            O => \N__10285\,
            I => \N__10278\
        );

    \I__1295\ : CEMux
    port map (
            O => \N__10284\,
            I => \N__10275\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10281\,
            I => \N__10270\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10278\,
            I => \N__10270\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__10275\,
            I => \N__10267\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__10270\,
            I => \N__10264\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__1289\ : Odrv4
    port map (
            O => \N__10264\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__10261\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__10250\,
            I => \N__10246\
        );

    \I__1284\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10243\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__10246\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__10243\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__10235\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10229\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__10229\,
            I => \uu2.mem0.w_data_0\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10223\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__10223\,
            I => \uu2.mem0.N_30_i_0\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__10220\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__10214\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10207\
        );

    \I__1271\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__10207\,
            I => \N__10198\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__10203\,
            I => \N__10194\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__10198\,
            I => \N__10190\
        );

    \I__1266\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10183\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10183\
        );

    \I__1264\ : InMux
    port map (
            O => \N__10193\,
            I => \N__10183\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__10190\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__10183\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \uu2.vbuf_raddr.un448_ci_0_cascade_\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__1259\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10168\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__10168\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__10165\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1255\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10157\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10157\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__10154\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__10151\,
            I => \N__10148\
        );

    \I__1251\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10143\
        );

    \I__1250\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10138\
        );

    \I__1249\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10138\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__10143\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__10138\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1246\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10127\
        );

    \I__1245\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10127\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10122\
        );

    \I__1243\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10117\
        );

    \I__1242\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10117\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__10122\,
            I => \uu2.un404_ci_0\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__10117\,
            I => \uu2.un404_ci_0\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__10112\,
            I => \N__10105\
        );

    \I__1238\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10100\
        );

    \I__1237\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10100\
        );

    \I__1236\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10095\
        );

    \I__1235\ : InMux
    port map (
            O => \N__10108\,
            I => \N__10095\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10092\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__10100\,
            I => \N__10087\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10095\,
            I => \N__10087\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__10092\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__10087\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__10082\,
            I => \uu2.un404_ci_0_cascade_\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__10078\,
            I => \N__10070\
        );

    \I__1226\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10067\
        );

    \I__1225\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10064\
        );

    \I__1224\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10061\
        );

    \I__1223\ : InMux
    port map (
            O => \N__10070\,
            I => \N__10058\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10053\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__10064\,
            I => \N__10053\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__10061\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__10058\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__10053\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \N__10043\
        );

    \I__1216\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10037\
        );

    \I__1215\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10032\
        );

    \I__1214\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10032\
        );

    \I__1213\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10029\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10037\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__10032\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__10029\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__10022\,
            I => \N__10019\
        );

    \I__1208\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10016\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10012\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__10012\,
            I => \N__10004\
        );

    \I__1204\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10001\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10008\,
            I => \N__9996\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9996\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__10004\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__10001\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__9996\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__1197\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__9983\,
            I => \N__9976\
        );

    \I__1195\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9971\
        );

    \I__1194\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9971\
        );

    \I__1193\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9966\
        );

    \I__1192\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9966\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__9976\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__9971\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9966\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__9959\,
            I => \N__9956\
        );

    \I__1187\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9953\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__1185\ : Span4Mux_s3_h
    port map (
            O => \N__9950\,
            I => \N__9942\
        );

    \I__1184\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9935\
        );

    \I__1183\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9935\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9935\
        );

    \I__1181\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9930\
        );

    \I__1180\ : InMux
    port map (
            O => \N__9945\,
            I => \N__9930\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__9942\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__9935\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__9930\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__9923\,
            I => \N__9918\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__9922\,
            I => \N__9915\
        );

    \I__1174\ : CascadeMux
    port map (
            O => \N__9921\,
            I => \N__9912\
        );

    \I__1173\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9909\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9904\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9904\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__9909\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9904\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1168\ : CEMux
    port map (
            O => \N__9899\,
            I => \N__9896\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__1166\ : Span4Mux_v
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__9890\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9887\,
            I => \N__9882\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9886\,
            I => \N__9879\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__9885\,
            I => \N__9875\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9882\,
            I => \N__9870\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__9879\,
            I => \N__9870\
        );

    \I__1159\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9865\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9865\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__9870\,
            I => \uu0.un154_ci_9\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__9865\,
            I => \uu0.un154_ci_9\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9851\
        );

    \I__1154\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9851\
        );

    \I__1153\ : InMux
    port map (
            O => \N__9858\,
            I => \N__9851\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__9851\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9845\,
            I => \N__9842\
        );

    \I__1149\ : Odrv12
    port map (
            O => \N__9842\,
            I => \uu0.un165_ci_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__9833\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1145\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__9827\,
            I => \N__9823\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9820\
        );

    \I__1142\ : Span4Mux_h
    port map (
            O => \N__9823\,
            I => \N__9817\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9820\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__9817\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__9812\,
            I => \uu2.trig_rd_is_det_cascade_\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__9809\,
            I => \N__9804\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__9808\,
            I => \N__9801\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9807\,
            I => \N__9798\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9795\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9792\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9798\,
            I => \N__9789\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9795\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__9792\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__9789\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__9782\,
            I => \N__9779\
        );

    \I__1128\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9773\
        );

    \I__1127\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9770\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9765\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9765\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9762\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9770\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__9765\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__9762\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1120\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9752\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__9752\,
            I => \uu0.un4_l_count_11\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__9746\,
            I => \uu0.un4_l_count_16\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__1115\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9730\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9730\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9730\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9737\,
            I => \N__9727\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9730\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__9727\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__9722\,
            I => \N__9717\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9714\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9707\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9707\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9707\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__9707\,
            I => \N__9704\
        );

    \I__1103\ : Odrv4
    port map (
            O => \N__9704\,
            I => \uu0.un198_ci_2\
        );

    \I__1102\ : CascadeMux
    port map (
            O => \N__9701\,
            I => \N__9696\
        );

    \I__1101\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9691\
        );

    \I__1100\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9691\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9688\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__9691\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9688\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__9683\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9676\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9676\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__9673\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9664\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9661\,
            I => \N__9655\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__9658\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__9655\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9641\
        );

    \I__1084\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9641\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9641\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__9641\,
            I => \N__9637\
        );

    \I__1081\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__9637\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9634\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__9629\,
            I => \N__9624\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9607\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9607\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9607\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9607\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9602\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9602\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9599\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9590\
        );

    \I__1069\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9590\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9590\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9590\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__9607\,
            I => \N__9587\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__9602\,
            I => \uu0.un110_ci\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9599\,
            I => \uu0.un110_ci\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9590\,
            I => \uu0.un110_ci\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__9587\,
            I => \uu0.un110_ci\
        );

    \I__1061\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9572\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9562\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9562\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9562\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9553\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9546\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9546\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9546\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9562\,
            I => \N__9543\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9538\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9538\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9531\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9531\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9531\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9528\
        );

    \I__1046\ : Odrv12
    port map (
            O => \N__9553\,
            I => \uu0.un4_l_count_0\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9546\,
            I => \uu0.un4_l_count_0\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9543\,
            I => \uu0.un4_l_count_0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9538\,
            I => \uu0.un4_l_count_0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9531\,
            I => \uu0.un4_l_count_0\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9528\,
            I => \uu0.un4_l_count_0\
        );

    \I__1040\ : CEMux
    port map (
            O => \N__9515\,
            I => \N__9503\
        );

    \I__1039\ : CEMux
    port map (
            O => \N__9514\,
            I => \N__9503\
        );

    \I__1038\ : CEMux
    port map (
            O => \N__9513\,
            I => \N__9503\
        );

    \I__1037\ : CEMux
    port map (
            O => \N__9512\,
            I => \N__9503\
        );

    \I__1036\ : GlobalMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__1035\ : gio2CtrlBuf
    port map (
            O => \N__9500\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__9497\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9486\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9486\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9483\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9480\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9486\,
            I => \uu0.un66_ci\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__9483\,
            I => \uu0.un66_ci\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9480\,
            I => \uu0.un66_ci\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9461\
        );

    \I__1025\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9461\
        );

    \I__1024\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9461\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9461\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__9461\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__9458\,
            I => \N__9453\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9448\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9448\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9445\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9448\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9445\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9434\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9431\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9438\,
            I => \N__9426\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9426\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9434\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9431\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9426\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1008\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9414\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9411\
        );

    \I__1006\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9408\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__9414\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__9411\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__9408\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9394\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9394\
        );

    \I__1000\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9391\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9394\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9391\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__997\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9383\,
            I => \uu0.un4_l_count_14\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__994\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9364\
        );

    \I__993\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9364\
        );

    \I__992\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9364\
        );

    \I__991\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9364\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__9373\,
            I => \N__9360\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9364\,
            I => \N__9357\
        );

    \I__988\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9354\
        );

    \I__987\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9351\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__9357\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9354\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__9351\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__983\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9341\,
            I => \uu0.un4_l_count_13\
        );

    \I__981\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9335\,
            I => \uu0.un4_l_count_12\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__9332\,
            I => \uu0.un4_l_count_18_cascade_\
        );

    \I__978\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__976\ : Odrv4
    port map (
            O => \N__9323\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__975\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9317\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__973\ : IoInMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9311\,
            I => \N__9308\
        );

    \I__971\ : Span4Mux_s0_h
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__970\ : Span4Mux_v
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__969\ : Odrv4
    port map (
            O => \N__9302\,
            I => o_serial_data_c
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__9299\,
            I => \N__9296\
        );

    \I__967\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9292\
        );

    \I__966\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9289\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9292\,
            I => \uu0.un88_ci_3\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9289\,
            I => \uu0.un88_ci_3\
        );

    \I__963\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9279\
        );

    \I__962\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9276\
        );

    \I__961\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9273\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9279\,
            I => \N__9270\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9276\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9273\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__957\ : Odrv4
    port map (
            O => \N__9270\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__9263\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9257\,
            I => vbuf_tx_data_0
        );

    \I__953\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9251\,
            I => vbuf_tx_data_7
        );

    \I__951\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9245\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__9242\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__948\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9236\,
            I => vbuf_tx_data_1
        );

    \I__946\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9230\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__944\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9224\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__942\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9218\,
            I => vbuf_tx_data_3
        );

    \I__940\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__9212\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__938\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9206\,
            I => vbuf_tx_data_4
        );

    \I__936\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__9200\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__934\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__9191\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__931\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__9185\,
            I => vbuf_tx_data_5
        );

    \I__929\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9179\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__9179\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__927\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9173\,
            I => \N__9170\
        );

    \I__925\ : Span12Mux_s2_h
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__924\ : Odrv12
    port map (
            O => \N__9167\,
            I => \uu2.r_data_wire_2\
        );

    \I__923\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__9161\,
            I => vbuf_tx_data_2
        );

    \I__921\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9151\
        );

    \I__920\ : InMux
    port map (
            O => \N__9157\,
            I => \N__9148\
        );

    \I__919\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9141\
        );

    \I__918\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9141\
        );

    \I__917\ : InMux
    port map (
            O => \N__9154\,
            I => \N__9141\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9151\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9148\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__9141\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9129\
        );

    \I__912\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9123\
        );

    \I__911\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9120\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__9129\,
            I => \N__9117\
        );

    \I__909\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9114\
        );

    \I__908\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9109\
        );

    \I__907\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9109\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__9123\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__9120\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__9117\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__9114\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__9109\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__901\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9092\
        );

    \I__900\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9092\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__9092\,
            I => \uu2.un284_ci\
        );

    \I__898\ : InMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__9083\,
            I => \uu2.r_data_wire_0\
        );

    \I__895\ : InMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__893\ : Odrv4
    port map (
            O => \N__9074\,
            I => \uu2.r_data_wire_1\
        );

    \I__892\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__890\ : Odrv4
    port map (
            O => \N__9065\,
            I => \uu2.r_data_wire_3\
        );

    \I__889\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__9059\,
            I => \uu2.r_data_wire_4\
        );

    \I__887\ : InMux
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__9053\,
            I => \uu2.r_data_wire_5\
        );

    \I__885\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__9047\,
            I => \uu2.r_data_wire_6\
        );

    \I__883\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9041\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__9038\,
            I => vbuf_tx_data_6
        );

    \I__880\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__9032\,
            I => \uu2.r_data_wire_7\
        );

    \I__878\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9026\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9023\
        );

    \I__876\ : IoSpan4Mux
    port map (
            O => \N__9023\,
            I => \N__9020\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__9020\,
            I => \uart_RXD\
        );

    \I__874\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9010\
        );

    \I__873\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9007\
        );

    \I__872\ : InMux
    port map (
            O => \N__9015\,
            I => \N__9000\
        );

    \I__871\ : InMux
    port map (
            O => \N__9014\,
            I => \N__9000\
        );

    \I__870\ : InMux
    port map (
            O => \N__9013\,
            I => \N__9000\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__9010\,
            I => \uu2.un306_ci\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9007\,
            I => \uu2.un306_ci\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__9000\,
            I => \uu2.un306_ci\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__8993\,
            I => \N__8987\
        );

    \I__865\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8983\
        );

    \I__864\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8980\
        );

    \I__863\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8977\
        );

    \I__862\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8972\
        );

    \I__861\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8972\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__8983\,
            I => \N__8969\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__8980\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__8977\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__8972\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__8969\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__855\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8955\
        );

    \I__854\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8952\
        );

    \I__853\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8949\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__8955\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__8952\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__8949\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__849\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8937\
        );

    \I__848\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8934\
        );

    \I__847\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8931\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__8937\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8934\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__8931\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8924\,
            I => \N__8919\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__8923\,
            I => \N__8916\
        );

    \I__841\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8909\
        );

    \I__840\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8909\
        );

    \I__839\ : InMux
    port map (
            O => \N__8916\,
            I => \N__8909\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__8909\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__8906\,
            I => \N__8900\
        );

    \I__836\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8890\
        );

    \I__835\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8890\
        );

    \I__834\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8890\
        );

    \I__833\ : InMux
    port map (
            O => \N__8900\,
            I => \N__8890\
        );

    \I__832\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8887\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8890\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8887\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__829\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8867\
        );

    \I__828\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8867\
        );

    \I__827\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8867\
        );

    \I__826\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8867\
        );

    \I__825\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8867\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__8867\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__823\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8854\
        );

    \I__822\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8854\
        );

    \I__821\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8854\
        );

    \I__820\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8851\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__8854\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8851\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__8846\,
            I => \N__8840\
        );

    \I__816\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8831\
        );

    \I__815\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8831\
        );

    \I__814\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8831\
        );

    \I__813\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8831\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8831\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__811\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8812\
        );

    \I__810\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8812\
        );

    \I__809\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8812\
        );

    \I__808\ : InMux
    port map (
            O => \N__8825\,
            I => \N__8812\
        );

    \I__807\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8812\
        );

    \I__806\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8809\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8812\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8809\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__803\ : InMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__8801\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__801\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8792\
        );

    \I__800\ : InMux
    port map (
            O => \N__8797\,
            I => \N__8792\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8792\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__798\ : IoInMux
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__796\ : Span4Mux_s0_h
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__8780\,
            I => \uu0.un11_l_count_i\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__8777\,
            I => \uu0.un88_ci_3_cascade_\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__8774\,
            I => \uu0.un55_ci_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__8771\,
            I => \N__8768\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__8768\,
            I => \uu0.un99_ci_0\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__8765\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__789\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8747\
        );

    \I__788\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8747\
        );

    \I__787\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8747\
        );

    \I__786\ : InMux
    port map (
            O => \N__8759\,
            I => \N__8747\
        );

    \I__785\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8747\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__8747\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8744\,
            I => \N__8739\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__8743\,
            I => \N__8736\
        );

    \I__781\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8729\
        );

    \I__780\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8729\
        );

    \I__779\ : InMux
    port map (
            O => \N__8736\,
            I => \N__8729\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__8726\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__776\ : InMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8720\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__773\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8707\
        );

    \I__772\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8707\
        );

    \I__771\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8704\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__8707\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8704\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8699\,
            I => \N__8694\
        );

    \I__767\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8689\
        );

    \I__766\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8689\
        );

    \I__765\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8686\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__8689\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8686\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__761\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8673\
        );

    \I__760\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8668\
        );

    \I__759\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8668\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8673\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__8668\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__755\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__8654\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__8651\,
            I => \N__8644\
        );

    \I__751\ : InMux
    port map (
            O => \N__8650\,
            I => \N__8641\
        );

    \I__750\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8632\
        );

    \I__749\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8632\
        );

    \I__748\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8632\
        );

    \I__747\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8632\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8641\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8632\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8621\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8621\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__8618\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__8615\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__738\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8606\,
            I => \uu2.un350_ci\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__8603\,
            I => \N__8598\
        );

    \I__735\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8591\
        );

    \I__734\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8591\
        );

    \I__733\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8591\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__8591\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__731\ : IoInMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8582\
        );

    \I__729\ : IoSpan4Mux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__8579\,
            I => clk_in_c
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__22346\
        );

    \INVuu2.bitmap_34C\ : INV
    port map (
            O => \INVuu2.bitmap_34C_net\,
            I => \N__22357\
        );

    \INVuu2.bitmap_218C\ : INV
    port map (
            O => \INVuu2.bitmap_218C_net\,
            I => \N__22328\
        );

    \INVuu2.bitmap_194C\ : INV
    port map (
            O => \INVuu2.bitmap_194C_net\,
            I => \N__22340\
        );

    \INVuu2.w_addr_displaying_2_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2_rep1C_net\,
            I => \N__22345\
        );

    \INVuu2.bitmap_87C\ : INV
    port map (
            O => \INVuu2.bitmap_87C_net\,
            I => \N__22351\
        );

    \INVuu2.bitmap_203C\ : INV
    port map (
            O => \INVuu2.bitmap_203C_net\,
            I => \N__22318\
        );

    \INVuu2.w_addr_displaying_fast_7C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_7C_net\,
            I => \N__22327\
        );

    \INVuu2.bitmap_90C\ : INV
    port map (
            O => \INVuu2.bitmap_90C_net\,
            I => \N__22334\
        );

    \INVuu2.w_addr_displaying_fast_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            I => \N__22339\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__22309\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__22317\
        );

    \INVuu2.bitmap_40C\ : INV
    port map (
            O => \INVuu2.bitmap_40C_net\,
            I => \N__22333\
        );

    \INVuu2.w_addr_displaying_nesr_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_8C_net\,
            I => \N__22338\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__22344\
        );

    \INVuu2.w_addr_user_0C\ : INV
    port map (
            O => \INVuu2.w_addr_user_0C_net\,
            I => \N__22350\
        );

    \INVuu2.w_addr_user_5C\ : INV
    port map (
            O => \INVuu2.w_addr_user_5C_net\,
            I => \N__22356\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__22312\
        );

    \INVuu2.w_addr_displaying_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4C_net\,
            I => \N__22337\
        );

    \INVuu2.r_data_reg_2C\ : INV
    port map (
            O => \INVuu2.r_data_reg_2C_net\,
            I => \N__22335\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__22347\
        );

    \IN_MUX_bfv_6_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_2_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_13_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10973\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12176\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8789\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14718\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8959\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8992\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8758\,
            in1 => \N__8986\,
            in2 => \N__8603\,
            in3 => \N__9126\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9013\,
            in1 => \N__8713\,
            in2 => \N__8743\,
            in3 => \N__8760\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8615\,
            in3 => \N__8697\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22361\,
            ce => 'H',
            sr => \N__22000\
        );

    \uu2.l_count_RNIBCGK1_9_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9127\,
            in1 => \N__8759\,
            in2 => \N__8993\,
            in3 => \N__8601\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8602\,
            in1 => \N__8698\,
            in2 => \N__8612\,
            in3 => \N__8942\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22361\,
            ce => 'H',
            sr => \N__22000\
        );

    \uu2.l_count_6_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__9014\,
            in1 => \_gnd_net_\,
            in2 => \N__8744\,
            in3 => \N__8761\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22361\,
            ce => 'H',
            sr => \N__22000\
        );

    \uu2.l_count_7_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8762\,
            in1 => \N__9015\,
            in2 => \N__8717\,
            in3 => \N__8742\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22361\,
            ce => 'H',
            sr => \N__22000\
        );

    \uu2.l_count_3_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__8650\,
            in1 => \N__8941\,
            in2 => \N__8681\,
            in3 => \N__9098\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22359\,
            ce => 'H',
            sr => \N__21997\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8677\,
            in1 => \N__9154\,
            in2 => \N__8651\,
            in3 => \N__9128\,
            lcout => \uu2.un306_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9097\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22359\,
            ce => 'H',
            sr => \N__21997\
        );

    \uu2.l_count_RNI9S834_0_1_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8647\,
            in1 => \N__8723\,
            in2 => \N__8663\,
            in3 => \N__9155\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIFGGK1_3_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8712\,
            in1 => \N__8958\,
            in2 => \N__8699\,
            in3 => \N__8676\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8648\,
            in1 => \N__9156\,
            in2 => \N__8627\,
            in3 => \N__8624\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9016\,
            in2 => \N__8618\,
            in3 => \N__8990\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22359\,
            ce => 'H',
            sr => \N__21997\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9295\,
            in2 => \_gnd_net_\,
            in3 => \N__9777\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9439\,
            in2 => \_gnd_net_\,
            in3 => \N__9282\,
            lcout => \uu0.un88_ci_3\,
            ltout => \uu0.un88_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9491\,
            in1 => \N__9776\,
            in2 => \N__8777\,
            in3 => \N__9418\,
            lcout => \uu0.un110_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8828\,
            in1 => \N__8905\,
            in2 => \_gnd_net_\,
            in3 => \N__8864\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__9513\,
            sr => \N__21990\
        );

    \uu0.l_count_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8827\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__9513\,
            sr => \N__21990\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8825\,
            in1 => \N__8903\,
            in2 => \_gnd_net_\,
            in3 => \N__8863\,
            lcout => OPEN,
            ltout => \uu0.un55_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_3_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9570\,
            in1 => \_gnd_net_\,
            in2 => \N__8774\,
            in3 => \N__9401\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__9513\,
            sr => \N__21990\
        );

    \uu0.l_count_0_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8826\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9569\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__9513\,
            sr => \N__21990\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8862\,
            in1 => \N__8824\,
            in2 => \N__8906\,
            in3 => \N__9400\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_7_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__8771\,
            in1 => \N__9419\,
            in2 => \N__8765\,
            in3 => \N__9571\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__9513\,
            sr => \N__21990\
        );

    \uu0.delay_line_0_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8879\,
            in1 => \N__9374\,
            in2 => \N__8924\,
            in3 => \N__8843\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \N__21992\
        );

    \uu0.l_precount_3_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8845\,
            in1 => \N__8922\,
            in2 => \N__9380\,
            in3 => \N__8882\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \N__21992\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8878\,
            in1 => \N__9284\,
            in2 => \N__8923\,
            in3 => \N__8899\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_1_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9375\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8880\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \N__21992\
        );

    \uu0.l_precount_2_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8881\,
            in1 => \N__9376\,
            in2 => \_gnd_net_\,
            in3 => \N__8844\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \N__21992\
        );

    \uu0.l_precount_RNI3Q7K1_2_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10490\,
            in1 => \N__8861\,
            in2 => \N__8846\,
            in3 => \N__8823\,
            lcout => \uu0.un4_l_count_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_1_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22313\,
            ce => 'H',
            sr => \N__21992\
        );

    \uu0.delay_line_RNILLLG7_1_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__8804\,
            in1 => \N__8797\,
            in2 => \_gnd_net_\,
            in3 => \N__9556\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_0_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9363\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22305\,
            ce => 'H',
            sr => \N__21995\
        );

    \buart.Z_rx.hh_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9029\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22297\,
            ce => 'H',
            sr => \N__21996\
        );

    \uu2.trig_rd_det_1_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9826\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22360\,
            ce => 'H',
            sr => \N__21973\
        );

    \uu2.l_count_5_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__9017\,
            in1 => \N__8960\,
            in2 => \_gnd_net_\,
            in3 => \N__8991\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22360\,
            ce => 'H',
            sr => \N__21973\
        );

    \uu2.l_count_0_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9132\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22360\,
            ce => 'H',
            sr => \N__21973\
        );

    \uu2.r_addr_5_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10133\,
            in1 => \N__10111\,
            in2 => \N__10078\,
            in3 => \N__10211\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \uu2.r_addr_4_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10110\,
            in1 => \N__10132\,
            in2 => \_gnd_net_\,
            in3 => \N__10210\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \uu2.trig_rd_det_0_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14870\,
            in2 => \_gnd_net_\,
            in3 => \N__10249\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \uu2.vram_rd_clk_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__14871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8940\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \uu0.sec_clk_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14916\,
            in2 => \_gnd_net_\,
            in3 => \N__9578\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \uu2.l_count_1_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9158\,
            in2 => \_gnd_net_\,
            in3 => \N__9133\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22358\,
            ce => 'H',
            sr => \N__21972\
        );

    \buart.Z_tx.shifter_7_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9248\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22352\,
            ce => \N__10284\,
            sr => \N__21999\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9134\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9080\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9071\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9056\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9050\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9035\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__10409\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9233\,
            in1 => \N__10596\,
            in2 => \_gnd_net_\,
            in3 => \N__9260\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_8_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10595\,
            in2 => \_gnd_net_\,
            in3 => \N__9254\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10597\,
            in1 => \N__9227\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9215\,
            in1 => \N__9164\,
            in2 => \_gnd_net_\,
            in3 => \N__10598\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_4_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10599\,
            in1 => \N__9203\,
            in2 => \_gnd_net_\,
            in3 => \N__9221\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_5_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9182\,
            in1 => \N__10600\,
            in2 => \_gnd_net_\,
            in3 => \N__9209\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \buart.Z_tx.shifter_6_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10601\,
            in1 => \N__9197\,
            in2 => \_gnd_net_\,
            in3 => \N__9188\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22342\,
            ce => \N__10285\,
            sr => \N__21994\
        );

    \uu2.r_data_reg_2_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9176\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_2C_net\,
            ce => \N__10405\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_0_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9329\,
            in2 => \_gnd_net_\,
            in3 => \N__10605\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => \N__10286\,
            sr => \N__21989\
        );

    \buart.Z_tx.uart_tx_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9320\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22330\,
            ce => \N__10286\,
            sr => \N__21989\
        );

    \uu0.l_count_11_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__10418\,
            in1 => \N__9617\,
            in2 => \N__9809\,
            in3 => \N__9575\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.l_count_8_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9616\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10484\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.l_count_9_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__10485\,
            in1 => \N__9619\,
            in2 => \_gnd_net_\,
            in3 => \N__10449\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.l_count_6_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9577\,
            in1 => \N__9494\,
            in2 => \N__9299\,
            in3 => \N__9778\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.l_count_5_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \N__9440\,
            in2 => \_gnd_net_\,
            in3 => \N__9283\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.l_count_13_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__9848\,
            in1 => \N__9618\,
            in2 => \N__9668\,
            in3 => \N__9576\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22323\,
            ce => \N__9512\,
            sr => \N__21991\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9878\,
            in1 => \N__9472\,
            in2 => \_gnd_net_\,
            in3 => \N__9649\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__9621\,
            in1 => \N__9457\,
            in2 => \N__9263\,
            in3 => \N__9560\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__9514\,
            sr => \N__21993\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9456\,
            in1 => \N__9471\,
            in2 => \N__9885\,
            in3 => \N__9648\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10444\,
            in1 => \N__10506\,
            in2 => \N__9808\,
            in3 => \N__10479\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9620\,
            in1 => \N__9473\,
            in2 => \N__9497\,
            in3 => \N__9650\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__9514\,
            sr => \N__21993\
        );

    \uu0.l_count_4_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9492\,
            in1 => \N__9438\,
            in2 => \_gnd_net_\,
            in3 => \N__9561\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__9514\,
            sr => \N__21993\
        );

    \uu0.l_count_10_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10480\,
            in1 => \N__9622\,
            in2 => \N__10513\,
            in3 => \N__10445\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__9514\,
            sr => \N__21993\
        );

    \uu0.l_count_RNIGTCU_15_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9470\,
            in1 => \N__10505\,
            in2 => \N__9458\,
            in3 => \N__9437\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10450\,
            in1 => \N__9417\,
            in2 => \N__9701\,
            in3 => \N__9399\,
            lcout => \uu0.un4_l_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIO2782_16_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9386\,
            in1 => \N__9737\,
            in2 => \N__9373\,
            in3 => \N__9640\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_15_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9344\,
            in1 => \N__9338\,
            in2 => \N__9332\,
            in3 => \N__9749\,
            lcout => \uu0.un4_l_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIOIDD2_18_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9807\,
            in1 => \N__9679\,
            in2 => \N__9782\,
            in3 => \N__9755\,
            lcout => \uu0.un4_l_count_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_2_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19863\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22306\,
            ce => \N__10733\,
            sr => \N__21970\
        );

    \resetGen.escKey_5_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23079\,
            in1 => \N__22877\,
            in2 => \N__19878\,
            in3 => \N__22546\,
            lcout => \resetGen.escKeyZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__9627\,
            in1 => \N__9739\,
            in2 => \N__9722\,
            in3 => \N__9558\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22298\,
            ce => \N__9515\,
            sr => \N__21998\
        );

    \uu0.l_count_17_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9700\,
            in1 => \N__9720\,
            in2 => \N__9743\,
            in3 => \N__9628\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22298\,
            ce => \N__9515\,
            sr => \N__21998\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9623\,
            in1 => \N__9738\,
            in2 => \N__9721\,
            in3 => \N__9699\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9559\,
            in1 => \_gnd_net_\,
            in2 => \N__9683\,
            in3 => \N__9680\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22298\,
            ce => \N__9515\,
            sr => \N__21998\
        );

    \uu0.l_count_RNIFAQ9_13_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9667\,
            in2 => \_gnd_net_\,
            in3 => \N__9858\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_12_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9860\,
            in1 => \N__9887\,
            in2 => \N__9629\,
            in3 => \N__9557\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22298\,
            ce => \N__9515\,
            sr => \N__21998\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9886\,
            in2 => \_gnd_net_\,
            in3 => \N__9859\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12163\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22291\,
            ce => 'H',
            sr => \N__22001\
        );

    \buart.Z_tx.bitcount_3_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__11091\,
            in1 => \N__10570\,
            in2 => \N__11120\,
            in3 => \N__10991\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \buart.Z_tx.bitcount_0_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__10569\,
            in1 => \N__11035\,
            in2 => \_gnd_net_\,
            in3 => \N__11090\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \buart.Z_tx.bitcount_2_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10568\,
            in2 => \_gnd_net_\,
            in3 => \N__10757\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \uu2.r_addr_2_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9982\,
            in1 => \N__10197\,
            in2 => \N__10015\,
            in3 => \N__9949\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9839\,
            in2 => \_gnd_net_\,
            in3 => \N__9830\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => \uu2.trig_rd_is_det_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9812\,
            in3 => \N__22038\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_1_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__9948\,
            in1 => \_gnd_net_\,
            in2 => \N__10203\,
            in3 => \N__9981\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \uu2.r_addr_0_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10193\,
            in2 => \_gnd_net_\,
            in3 => \N__9947\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22355\,
            ce => 'H',
            sr => \N__21981\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10146\,
            in2 => \_gnd_net_\,
            in3 => \N__10040\,
            lcout => OPEN,
            ltout => \uu2.vbuf_raddr.un448_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__10171\,
            in1 => \N__10160\,
            in2 => \N__10178\,
            in3 => \N__10125\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__9899\,
            sr => \N__21976\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10076\,
            in2 => \_gnd_net_\,
            in3 => \N__10108\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_7_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__10147\,
            in1 => \N__10041\,
            in2 => \N__10154\,
            in3 => \N__10126\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__9899\,
            sr => \N__21976\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10007\,
            in1 => \N__9979\,
            in2 => \N__9921\,
            in3 => \N__9945\,
            lcout => \uu2.un404_ci_0\,
            ltout => \uu2.un404_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10109\,
            in1 => \N__10042\,
            in2 => \N__10082\,
            in3 => \N__10077\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__9899\,
            sr => \N__21976\
        );

    \uu2.r_addr_esr_3_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10008\,
            in1 => \N__9980\,
            in2 => \N__9922\,
            in3 => \N__9946\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__9899\,
            sr => \N__21976\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14248\,
            in1 => \N__14387\,
            in2 => \N__14348\,
            in3 => \N__14305\,
            lcout => \uu2.un404_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10544\,
            in2 => \_gnd_net_\,
            in3 => \N__11092\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__22040\,
            in1 => \N__14882\,
            in2 => \N__10567\,
            in3 => \N__10256\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22343\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__15859\,
            in1 => \N__12352\,
            in2 => \N__11252\,
            in3 => \N__15947\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__12353\,
            in1 => \N__12467\,
            in2 => \N__15983\,
            in3 => \N__15860\,
            lcout => \uu2.mem0.w_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__15858\,
            in1 => \N__15948\,
            in2 => \N__12566\,
            in3 => \N__11273\,
            lcout => \uu2.mem0.N_30_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__12482\,
            in1 => \N__15857\,
            in2 => \N__15982\,
            in3 => \N__16787\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011010110010"
        )
    port map (
            in0 => \N__12562\,
            in1 => \N__11159\,
            in2 => \N__10220\,
            in3 => \N__11129\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec2_1_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11813\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.sec2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110000"
        )
    port map (
            in0 => \N__12512\,
            in1 => \N__13497\,
            in2 => \N__14947\,
            in3 => \N__11586\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m32_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010111111110"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__11594\,
            in2 => \N__10310\,
            in3 => \N__11326\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100110011"
        )
    port map (
            in0 => \N__10649\,
            in1 => \N__11584\,
            in2 => \N__10307\,
            in3 => \N__11479\,
            lcout => \Lab_UT.dispString.m40_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec1_3_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11720\,
            lcout => \Lab_UT.sec1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__11227\,
            in1 => \N__11585\,
            in2 => \N__10298\,
            in3 => \N__11480\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11325\,
            in2 => \N__10289\,
            in3 => \N__10331\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min2_0_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12035\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.min2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_5_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12584\,
            lcout => \Lab_UT.alarmcharZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__14675\,
            in1 => \N__14580\,
            in2 => \N__10385\,
            in3 => \N__14548\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min2_2_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11984\,
            lcout => \Lab_UT.min2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_5_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100110000"
        )
    port map (
            in0 => \N__10340\,
            in1 => \N__13498\,
            in2 => \N__14948\,
            in3 => \N__11589\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m35_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011101111110"
        )
    port map (
            in0 => \N__11590\,
            in1 => \N__11327\,
            in2 => \N__10334\,
            in3 => \N__11478\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__11476\,
            in1 => \N__10316\,
            in2 => \N__10325\,
            in3 => \N__11587\,
            lcout => \Lab_UT.dispString.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110111"
        )
    port map (
            in0 => \N__11588\,
            in1 => \N__11477\,
            in2 => \N__14735\,
            in3 => \N__10373\,
            lcout => \Lab_UT.dispString.dOut_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14579\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22331\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16336\,
            in1 => \N__11583\,
            in2 => \N__11333\,
            in3 => \N__11475\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec1_2_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10672\,
            lcout => \Lab_UT.sec1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec2_0_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10751\,
            lcout => \Lab_UT.sec2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_0_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12878\,
            lcout => \Lab_UT.alarmcharZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12785\,
            in2 => \_gnd_net_\,
            in3 => \N__12754\,
            lcout => \Lab_UT.alarmcharZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__10637\,
            in1 => \N__11442\,
            in2 => \N__10367\,
            in3 => \N__16335\,
            lcout => \Lab_UT.dispString.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min2_1_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12008\,
            lcout => \Lab_UT.min2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110001110111"
        )
    port map (
            in0 => \N__10358\,
            in1 => \N__11441\,
            in2 => \N__10352\,
            in3 => \N__11547\,
            lcout => \Lab_UT.dispString.m25_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110010"
        )
    port map (
            in0 => \N__11591\,
            in1 => \N__11473\,
            in2 => \N__11332\,
            in3 => \N__16344\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \Lab_UT.didp.regrce2.q_2_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__19877\,
            in1 => \N__20725\,
            in2 => \N__16391\,
            in3 => \N__10671\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \Lab_UT.didp.regrce2.q_3_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__20726\,
            in1 => \N__16389\,
            in2 => \N__19424\,
            in3 => \N__11716\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \Lab_UT.dictrl.state_0_RNIRNP_1_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21453\,
            in2 => \_gnd_net_\,
            in3 => \N__21123\,
            lcout => \Lab_UT.dicLdAStens_0\,
            ltout => \Lab_UT.dicLdAStens_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_1_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__22768\,
            in1 => \N__16385\,
            in2 => \N__10343\,
            in3 => \N__14752\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \Lab_UT.dispString.cnt_2_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11472\,
            in1 => \N__11321\,
            in2 => \_gnd_net_\,
            in3 => \N__11593\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \Lab_UT.dispString.cnt_1_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11592\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11474\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \buart.Z_tx.bitcount_1_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111111100"
        )
    port map (
            in0 => \N__11036\,
            in1 => \N__11050\,
            in2 => \N__10607\,
            in3 => \N__11096\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => 'H',
            sr => \N__21969\
        );

    \buart.Z_rx.bitcount_es_2_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001010010111110"
        )
    port map (
            in0 => \N__10808\,
            in1 => \N__10885\,
            in2 => \N__10859\,
            in3 => \N__13600\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => \N__12119\,
            sr => \N__22035\
        );

    \buart.Z_rx.bitcount_es_0_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__13599\,
            in1 => \N__10807\,
            in2 => \N__12648\,
            in3 => \N__12205\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22307\,
            ce => \N__12119\,
            sr => \N__22035\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10517\,
            in1 => \N__10489\,
            in2 => \_gnd_net_\,
            in3 => \N__10451\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14831\,
            in1 => \N__14849\,
            in2 => \_gnd_net_\,
            in3 => \N__22034\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m27_1_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23202\,
            in2 => \_gnd_net_\,
            in3 => \N__20414\,
            lcout => \Lab_UT.dictrl.m27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14519\,
            in2 => \_gnd_net_\,
            in3 => \N__14619\,
            lcout => \resetGen.reset_count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__13454\,
            in1 => \N__10697\,
            in2 => \N__13340\,
            in3 => \N__15142\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.un1_num_5_2_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15046\,
            in2 => \_gnd_net_\,
            in3 => \N__15229\,
            lcout => OPEN,
            ltout => \Lab_UT.three_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIGRQR1_2_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19874\,
            in1 => \N__15453\,
            in2 => \N__10700\,
            in3 => \N__15141\,
            lcout => \Lab_UT.didp.countrce3.q_5_2\,
            ltout => \Lab_UT.didp.countrce3.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_2_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__10687\,
            in1 => \N__13453\,
            in2 => \N__10691\,
            in3 => \N__13339\,
            lcout => \Lab_UT.didp.countrce3.q_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_RNII6JA1_2_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__11755\,
            in1 => \N__10750\,
            in2 => \N__10688\,
            in3 => \N__11980\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.did_alarmMatch_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIQTCC2_2_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__12971\,
            in1 => \N__10673\,
            in2 => \N__10652\,
            in3 => \N__10628\,
            lcout => \Lab_UT.didp.did_alarmMatch_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNISLCD1_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__15230\,
            in1 => \N__15452\,
            in2 => \N__15047\,
            in3 => \N__22766\,
            lcout => \Lab_UT.didp.countrce3.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min2_3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11944\,
            lcout => \Lab_UT.min2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22299\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min1_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11857\,
            lcout => \Lab_UT.min1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec2_2_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10627\,
            lcout => \Lab_UT.sec2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22292\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16160\,
            in2 => \_gnd_net_\,
            in3 => \N__22037\,
            lcout => \Lab_UT.didp.regrce1.LdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_0_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16491\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22286\,
            ce => \N__10723\,
            sr => \N__21974\
        );

    \Lab_UT.didp.regrce1.q_esr_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22286\,
            ce => \N__10723\,
            sr => \N__21974\
        );

    \Lab_UT.didp.regrce1.q_esr_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19419\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22286\,
            ce => \N__10723\,
            sr => \N__21974\
        );

    \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10773\,
            in2 => \_gnd_net_\,
            in3 => \N__12206\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10887\,
            in1 => \N__10841\,
            in2 => \N__10712\,
            in3 => \N__10917\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10916\,
            in1 => \N__10886\,
            in2 => \N__10844\,
            in3 => \N__10772\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOUCP_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10837\,
            in2 => \_gnd_net_\,
            in3 => \N__10915\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10888\,
            in1 => \N__10774\,
            in2 => \N__10709\,
            in3 => \N__12207\,
            lcout => \buart.Z_rx.idle\,
            ltout => \buart.Z_rx.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIOP0V3_1_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10706\,
            in3 => \N__12136\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => \buart.Z_rx.N_27_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_1_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__10898\,
            in2 => \N__10703\,
            in3 => \N__13586\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22281\,
            ce => \N__12114\,
            sr => \N__22002\
        );

    \buart.Z_rx.bitcount_es_3_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__13585\,
            in1 => \N__10797\,
            in2 => \N__10820\,
            in3 => \N__10842\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22281\,
            ce => \N__12114\,
            sr => \N__22002\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12208\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10919\,
            in2 => \_gnd_net_\,
            in3 => \N__10892\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10889\,
            in2 => \_gnd_net_\,
            in3 => \N__10847\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10843\,
            in2 => \_gnd_net_\,
            in3 => \N__10811\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__10798\,
            in1 => \N__13587\,
            in2 => \N__10778\,
            in3 => \N__10781\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22277\,
            ce => \N__12115\,
            sr => \N__22003\
        );

    \buart.Z_rx.shifter_fast_6_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23072\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22273\,
            ce => \N__22073\,
            sr => \N__22004\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100111001100"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__11002\,
            in2 => \N__11063\,
            in3 => \N__11083\,
            lcout => \buart.Z_tx.bitcount_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__12076\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12055\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11116\,
            in2 => \_gnd_net_\,
            in3 => \N__11029\,
            lcout => \buart.Z_tx.uart_busy_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__12054\,
            in1 => \N__12074\,
            in2 => \N__12341\,
            in3 => \N__12257\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => \buart.Z_tx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__11001\,
            in1 => \N__11058\,
            in2 => \N__11105\,
            in3 => \N__11102\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__11062\,
            in1 => \N__11031\,
            in2 => \N__11006\,
            in3 => \N__11003\,
            lcout => \buart.Z_tx.un1_bitcount_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22349\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__15979\,
            in1 => \N__17421\,
            in2 => \N__14306\,
            in3 => \N__15837\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__15836\,
            in1 => \N__10969\,
            in2 => \_gnd_net_\,
            in3 => \N__15978\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__17492\,
            in2 => \N__14186\,
            in3 => \N__15838\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_29_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12359\,
            in1 => \N__12383\,
            in2 => \_gnd_net_\,
            in3 => \N__12404\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_i7_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_19_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001110001001"
        )
    port map (
            in0 => \N__15977\,
            in1 => \N__12556\,
            in2 => \N__11162\,
            in3 => \N__15835\,
            lcout => \uu2.mem0.w_data_0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__15839\,
            in1 => \N__15981\,
            in2 => \N__14216\,
            in3 => \N__17253\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_36_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17424\,
            in2 => \_gnd_net_\,
            in3 => \N__17486\,
            lcout => \uu2.mem0.bitmap_pmux_sn_N_33_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_37_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110111110"
        )
    port map (
            in0 => \N__17487\,
            in1 => \N__17912\,
            in2 => \N__18119\,
            in3 => \N__17173\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_m24_0_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_26_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100000000110"
        )
    port map (
            in0 => \N__17913\,
            in1 => \N__11141\,
            in2 => \N__11135\,
            in3 => \N__18111\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_i5_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__16969\,
            in1 => \N__17645\,
            in2 => \N__11132\,
            in3 => \N__16127\,
            lcout => \uu2.mem0.N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__17172\,
            in1 => \N__18112\,
            in2 => \N__17921\,
            in3 => \N__17425\,
            lcout => \uu2.N_34\,
            ltout => \uu2.N_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010011010100110"
        )
    port map (
            in0 => \N__17488\,
            in1 => \N__17316\,
            in2 => \N__11123\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__21943\
        );

    \uu2.w_addr_displaying_2_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__17917\,
            in1 => \N__17178\,
            in2 => \N__17321\,
            in3 => \N__17426\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__21943\
        );

    \uu2.w_addr_displaying_5_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__17489\,
            in1 => \N__17320\,
            in2 => \N__12377\,
            in3 => \N__17255\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__21943\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__11168\,
            in2 => \N__11228\,
            in3 => \N__11600\,
            lcout => \Lab_UT.dispString.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_4_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11268\,
            in1 => \N__17073\,
            in2 => \N__12503\,
            in3 => \N__11244\,
            lcout => \uu2.un1_w_user_crZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min1_3_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11831\,
            lcout => \Lab_UT.min1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__15961\,
            in1 => \N__18113\,
            in2 => \N__14255\,
            in3 => \N__15825\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14941\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0_sec_clkD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101010101"
        )
    port map (
            in0 => \N__11192\,
            in1 => \N__11490\,
            in2 => \N__11186\,
            in3 => \N__16346\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11331\,
            in2 => \N__11177\,
            in3 => \N__11174\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec2_3_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11684\,
            lcout => \Lab_UT.sec2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22332\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100001010000"
        )
    port map (
            in0 => \N__11348\,
            in1 => \N__11639\,
            in2 => \N__11491\,
            in3 => \N__16345\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__11328\,
            in1 => \_gnd_net_\,
            in2 => \N__11366\,
            in3 => \N__11363\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100110011"
        )
    port map (
            in0 => \N__11354\,
            in1 => \N__11595\,
            in2 => \N__11342\,
            in3 => \N__11482\,
            lcout => \Lab_UT.dispString.m49_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011010010"
        )
    port map (
            in0 => \N__14674\,
            in1 => \N__14581\,
            in2 => \N__14621\,
            in3 => \N__14547\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__11615\,
            in1 => \N__11329\,
            in2 => \_gnd_net_\,
            in3 => \N__11390\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec1_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12716\,
            lcout => \Lab_UT.sec1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11606\,
            in1 => \N__11596\,
            in2 => \N__11492\,
            in3 => \N__11330\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22325\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12463\,
            in1 => \N__11269\,
            in2 => \N__12437\,
            in3 => \N__11245\,
            lcout => \uu2.un1_w_user_lfZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min1_2_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11843\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.min1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNI8QDI1_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__12711\,
            in1 => \N__11842\,
            in2 => \N__20345\,
            in3 => \N__11751\,
            lcout => \Lab_UT.didp.regrce4.did_alarmMatch_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNIJRBC_1_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13150\,
            in1 => \N__13063\,
            in2 => \_gnd_net_\,
            in3 => \N__12970\,
            lcout => \Lab_UT.didp.countrce2.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_2_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12599\,
            lcout => \Lab_UT.alarmcharZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.min1_0_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11876\,
            lcout => \Lab_UT.min1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010001000100"
        )
    port map (
            in0 => \N__11633\,
            in1 => \N__11471\,
            in2 => \N__11624\,
            in3 => \N__16337\,
            lcout => \Lab_UT.dispString.N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12722\,
            lcout => \Lab_UT.alarmcharZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22316\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__11582\,
            in1 => \N__11513\,
            in2 => \N__11507\,
            in3 => \N__11470\,
            lcout => \Lab_UT.dispString.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__15223\,
            in1 => \N__11875\,
            in2 => \N__20140\,
            in3 => \N__12031\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIRSKRA_0_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11384\,
            in1 => \N__11378\,
            in2 => \N__11369\,
            in3 => \N__11645\,
            lcout => \Lab_UT.alarmMatch\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_fast_0_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__13277\,
            in1 => \N__12092\,
            in2 => \N__11759\,
            in3 => \N__13791\,
            lcout => \Lab_UT.didp.q_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNIUST81_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__11732\,
            in1 => \N__19423\,
            in2 => \N__18716\,
            in3 => \N__13004\,
            lcout => \Lab_UT.didp.countrce2.q_5_3\,
            ltout => \Lab_UT.didp.countrce2.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_fast_3_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__13278\,
            in1 => \N__11699\,
            in2 => \N__11723\,
            in3 => \N__13792\,
            lcout => \Lab_UT.didp.countrce2.q_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_fast_RNIOS8A1_3_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__11715\,
            in1 => \N__11695\,
            in2 => \_gnd_net_\,
            in3 => \N__11683\,
            lcout => \Lab_UT.didp.did_alarmMatch_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__13005\,
            in1 => \N__13790\,
            in2 => \N__13283\,
            in3 => \N__11660\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__12091\,
            in1 => \N__13279\,
            in2 => \N__13793\,
            in3 => \N__13068\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22308\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_RNINLQC1_1_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__11773\,
            in1 => \N__11858\,
            in2 => \N__12904\,
            in3 => \N__12004\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.did_alarmMatch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_RNI077E5_1_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11654\,
            in1 => \N__11795\,
            in2 => \N__11648\,
            in3 => \N__11882\,
            lcout => \Lab_UT.didp.did_alarmMatch_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.un1_num_5_2_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13133\,
            in2 => \_gnd_net_\,
            in3 => \N__13064\,
            lcout => OPEN,
            ltout => \Lab_UT.three_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__18704\,
            in1 => \N__19872\,
            in2 => \N__11816\,
            in3 => \N__12959\,
            lcout => \Lab_UT.didp.countrce2.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_fast_RNIIM8A1_1_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__11785\,
            in1 => \N__14751\,
            in2 => \_gnd_net_\,
            in3 => \N__11812\,
            lcout => \Lab_UT.didp.did_alarmMatch_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_fast_1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__13274\,
            in1 => \N__12695\,
            in2 => \N__11789\,
            in3 => \N__13776\,
            lcout => \Lab_UT.didp.countrce2.q_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__12694\,
            in1 => \N__13275\,
            in2 => \N__13786\,
            in3 => \N__13134\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22300\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__13449\,
            in1 => \N__13327\,
            in2 => \N__13181\,
            in3 => \N__11774\,
            lcout => \Lab_UT.didp.countrce3.q_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_fast_3_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__11893\,
            in1 => \N__13396\,
            in2 => \N__13226\,
            in3 => \N__13192\,
            lcout => \Lab_UT.didp.q_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIMAAB1_2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15139\,
            in1 => \N__15033\,
            in2 => \_gnd_net_\,
            in3 => \N__15219\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNI529A2_3_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__15086\,
            in1 => \N__19414\,
            in2 => \N__11762\,
            in3 => \N__15454\,
            lcout => \Lab_UT.didp.countrce3.q_5_3\,
            ltout => \Lab_UT.didp.countrce3.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_3_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__13450\,
            in1 => \N__13328\,
            in2 => \N__11906\,
            in3 => \N__11903\,
            lcout => \Lab_UT.didp.countrce3.q_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_fast_RNIVTQC1_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__11902\,
            in1 => \N__11827\,
            in2 => \N__11894\,
            in3 => \N__11943\,
            lcout => \Lab_UT.didp.countrce3.did_alarmMatch_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__13397\,
            in1 => \N__13508\,
            in2 => \N__20123\,
            in3 => \N__13221\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22293\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.un1_num_11_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15220\,
            in1 => \N__15140\,
            in2 => \N__15109\,
            in3 => \N__15032\,
            lcout => \Lab_UT.nine_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_0_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16489\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22287\,
            ce => \N__13478\,
            sr => \N__21975\
        );

    \Lab_UT.didp.regrce4.q_esr_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22767\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22287\,
            ce => \N__13478\,
            sr => \N__21975\
        );

    \Lab_UT.didp.regrce4.q_esr_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19876\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22287\,
            ce => \N__13478\,
            sr => \N__21975\
        );

    \Lab_UT.didp.regrce4.q_esr_3_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19407\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22287\,
            ce => \N__13478\,
            sr => \N__21975\
        );

    \Lab_UT.didp.ce_11_2_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__15440\,
            in1 => \N__21429\,
            in2 => \N__15377\,
            in3 => \N__20655\,
            lcout => \Lab_UT.didp.ce_11_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_RNI0RGF_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15376\,
            lcout => \Lab_UT.dicLdAMones_0\,
            ltout => \Lab_UT.dicLdAMones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_0_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__16493\,
            in1 => \N__20657\,
            in2 => \N__12038\,
            in3 => \N__12027\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => 'H',
            sr => \N__21977\
        );

    \Lab_UT.didp.regrce3.q_1_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100001000"
        )
    port map (
            in0 => \N__22706\,
            in1 => \N__11955\,
            in2 => \N__20666\,
            in3 => \N__12003\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => 'H',
            sr => \N__21977\
        );

    \Lab_UT.didp.regrce3.q_2_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111100100000"
        )
    port map (
            in0 => \N__19875\,
            in1 => \N__20658\,
            in2 => \N__11960\,
            in3 => \N__11979\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => 'H',
            sr => \N__21977\
        );

    \Lab_UT.didp.regrce3.q_3_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__20656\,
            in1 => \N__19402\,
            in2 => \N__11945\,
            in3 => \N__11959\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => 'H',
            sr => \N__21977\
        );

    \resetGen.escKey_4_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16492\,
            in1 => \N__22705\,
            in2 => \N__19418\,
            in3 => \N__22460\,
            lcout => OPEN,
            ltout => \resetGen.escKeyZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11921\,
            in2 => \N__11909\,
            in3 => \N__12135\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__13580\,
            in1 => \N__13637\,
            in2 => \N__13627\,
            in3 => \N__13651\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__13723\,
            in1 => \N__13581\,
            in2 => \_gnd_net_\,
            in3 => \N__13738\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000010"
        )
    port map (
            in0 => \N__13690\,
            in1 => \N__13628\,
            in2 => \N__13598\,
            in3 => \N__13676\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22278\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__13666\,
            in1 => \N__13689\,
            in2 => \N__13528\,
            in3 => \N__13737\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13650\,
            in2 => \N__12224\,
            in3 => \N__13722\,
            lcout => \buart.Z_rx.ser_clk\,
            ltout => \buart.Z_rx.ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12221\,
            in2 => \N__12215\,
            in3 => \N__12212\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNIJ3K62_0_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13867\,
            in1 => \N__12164\,
            in2 => \_gnd_net_\,
            in3 => \N__12148\,
            lcout => \buart.Z_rx.startbit\,
            ltout => \buart.Z_rx.startbit_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__12149\,
            in1 => \N__13619\,
            in2 => \N__12140\,
            in3 => \N__12137\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI5RHS_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__18712\,
            in1 => \N__16450\,
            in2 => \_gnd_net_\,
            in3 => \N__13084\,
            lcout => \Lab_UT.didp.countrce2.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIINVH_2_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__14332\,
            in1 => \N__13907\,
            in2 => \N__14177\,
            in3 => \N__12302\,
            lcout => \uu2.un3_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12077\,
            in2 => \N__12059\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_2_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12266\,
            in2 => \_gnd_net_\,
            in3 => \N__12041\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__22341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12315\,
            in1 => \N__12340\,
            in2 => \_gnd_net_\,
            in3 => \N__12326\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__22341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12287\,
            in2 => \_gnd_net_\,
            in3 => \N__12323\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__22341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12316\,
            in1 => \N__12296\,
            in2 => \_gnd_net_\,
            in3 => \N__12320\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__22341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__12277\,
            in1 => \N__12317\,
            in2 => \_gnd_net_\,
            in3 => \N__12305\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22341\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI9006_8_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__14085\,
            in1 => \N__14483\,
            in2 => \_gnd_net_\,
            in3 => \N__14283\,
            lcout => \uu2.un3_w_addr_user_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12295\,
            in1 => \N__12286\,
            in2 => \N__12278\,
            in3 => \N__12265\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__16118\,
            in1 => \N__14086\,
            in2 => \N__15856\,
            in3 => \N__15988\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__14370\,
            in2 => \N__15995\,
            in3 => \N__15844\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_44_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000100000000"
        )
    port map (
            in0 => \N__17558\,
            in1 => \N__17919\,
            in2 => \N__18118\,
            in3 => \N__13988\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__15987\,
            in1 => \N__17174\,
            in2 => \N__14341\,
            in3 => \N__15840\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_31_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__17249\,
            in1 => \N__16970\,
            in2 => \N__15689\,
            in3 => \N__16117\,
            lcout => \uu2.mem0.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_51_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17476\,
            in2 => \_gnd_net_\,
            in3 => \N__17765\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_43_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010101000"
        )
    port map (
            in0 => \N__16801\,
            in1 => \N__18104\,
            in2 => \N__12386\,
            in3 => \N__17557\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_RNIGIDK3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15984\,
            in2 => \_gnd_net_\,
            in3 => \N__15803\,
            lcout => \N_272_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI17I72_5_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__17491\,
            in1 => \_gnd_net_\,
            in2 => \N__12376\,
            in3 => \N__17254\,
            lcout => \uu2.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_42_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110001000"
        )
    port map (
            in0 => \N__17171\,
            in1 => \N__17422\,
            in2 => \_gnd_net_\,
            in3 => \N__17490\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIB2283_5_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15741\,
            in1 => \N__12526\,
            in2 => \_gnd_net_\,
            in3 => \N__18296\,
            lcout => \uu2.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIEHP31_6_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15681\,
            in1 => \N__16968\,
            in2 => \_gnd_net_\,
            in3 => \N__16121\,
            lcout => \uu2.N_57\,
            ltout => \uu2.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIFOBB3_1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__12525\,
            in1 => \N__17918\,
            in2 => \N__12569\,
            in3 => \N__17423\,
            lcout => \uu2.w_data_i_a3_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_21_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__17396\,
            in1 => \_gnd_net_\,
            in2 => \N__15748\,
            in3 => \N__12527\,
            lcout => OPEN,
            ltout => \uu2.mem0.w_data_0_a3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011011000"
        )
    port map (
            in0 => \N__15993\,
            in1 => \N__12502\,
            in2 => \N__12545\,
            in3 => \N__15828\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNITJLE1_5_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17485\,
            in1 => \N__17180\,
            in2 => \N__18116\,
            in3 => \N__17248\,
            lcout => \uu2.w_data_displaying_2_i_a2_i_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_4_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12593\,
            lcout => \Lab_UT.alarmcharZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22320\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12480\,
            in2 => \_gnd_net_\,
            in3 => \N__12501\,
            lcout => \uu2.un1_w_user_lf_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_cr_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12481\,
            in1 => \N__12462\,
            in2 => \N__12436\,
            in3 => \N__12446\,
            lcout => uu2_un1_w_user_cr_0,
            ltout => \uu2_un1_w_user_cr_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15992\,
            in2 => \N__12440\,
            in3 => \N__12432\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIGEPH1_2_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101000001000"
        )
    port map (
            in0 => \N__17179\,
            in1 => \N__17395\,
            in2 => \N__18103\,
            in3 => \N__17484\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_0_2_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011011110111"
        )
    port map (
            in0 => \N__12968\,
            in1 => \N__13017\,
            in2 => \N__13102\,
            in3 => \N__13156\,
            lcout => \Lab_UT.bcd2segment2.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_4_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__13151\,
            in1 => \N__13085\,
            in2 => \N__13022\,
            in3 => \N__12963\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_5_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110011000"
        )
    port map (
            in0 => \N__12964\,
            in1 => \N__13009\,
            in2 => \N__13100\,
            in3 => \N__13152\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_6_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010100101"
        )
    port map (
            in0 => \N__13153\,
            in1 => \N__13089\,
            in2 => \N__13023\,
            in3 => \N__12965\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_0_0_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111101101101"
        )
    port map (
            in0 => \N__12966\,
            in1 => \N__13013\,
            in2 => \N__13101\,
            in3 => \N__13154\,
            lcout => \Lab_UT.bcd2segment2.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_0_1_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100101111111"
        )
    port map (
            in0 => \N__13155\,
            in1 => \N__13093\,
            in2 => \N__13024\,
            in3 => \N__12967\,
            lcout => \Lab_UT.bcd2segment2.segment_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_3_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011011010"
        )
    port map (
            in0 => \N__12969\,
            in1 => \N__13018\,
            in2 => \N__13103\,
            in3 => \N__13157\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment2.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12572\,
            in3 => \N__20058\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__21940\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__G_64_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__12850\,
            in1 => \N__12803\,
            in2 => \N__14790\,
            in3 => \N__14722\,
            lcout => \Lab_UT.dictrl.G_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.next_alarmstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22304\,
            ce => \N__12623\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__m6_xx_mm_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001110"
        )
    port map (
            in0 => \N__12614\,
            in1 => \N__12743\,
            in2 => \N__12781\,
            in3 => \N__16415\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12773\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__12613\,
            in1 => \N__12867\,
            in2 => \N__12605\,
            in3 => \N__16414\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1_0\,
            ltout => \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNINRI3E_0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14774\,
            in2 => \N__12602\,
            in3 => \N__12823\,
            lcout => \Lab_UT.dictrl.next_alarmstate_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNIT8JUD_0_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__14775\,
            in1 => \_gnd_net_\,
            in2 => \N__12830\,
            in3 => \N__12802\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__12744\,
            in1 => \_gnd_net_\,
            in2 => \N__12874\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmchar9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14794\,
            in1 => \N__12852\,
            in2 => \_gnd_net_\,
            in3 => \N__12805\,
            lcout => \Lab_UT.alarmchar10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.dictrl.alarmstate_ret_2_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__12806\,
            in1 => \N__14795\,
            in2 => \_gnd_net_\,
            in3 => \N__12853\,
            lcout => \Lab_UT.alarmchar10_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.dictrl.alarmstate_0_0_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14791\,
            in1 => \N__12827\,
            in2 => \_gnd_net_\,
            in3 => \N__12851\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.dictrl.alarmstate_ret_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__12829\,
            in1 => \N__14793\,
            in2 => \_gnd_net_\,
            in3 => \N__12854\,
            lcout => \Lab_UT.dictrl.alarmstate_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.dictrl.alarmstate_0_1_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14792\,
            in1 => \N__12828\,
            in2 => \_gnd_net_\,
            in3 => \N__12804\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12777\,
            in2 => \_gnd_net_\,
            in3 => \N__12745\,
            lcout => \Lab_UT.alarmchar_2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__15455\,
            in1 => \N__16474\,
            in2 => \_gnd_net_\,
            in3 => \N__15221\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_0_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__16475\,
            in1 => \N__20727\,
            in2 => \N__16390\,
            in3 => \N__12712\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22295\,
            ce => 'H',
            sr => \N__21971\
        );

    \Lab_UT.didp.countrce2.q_RNINQL01_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__13062\,
            in1 => \N__13132\,
            in2 => \N__18705\,
            in3 => \N__22737\,
            lcout => \Lab_UT.didp.countrce2.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.un1_num_5_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18344\,
            in2 => \_gnd_net_\,
            in3 => \N__18462\,
            lcout => \Lab_UT.three_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__12958\,
            in1 => \N__13764\,
            in2 => \N__12686\,
            in3 => \N__13276\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__13451\,
            in1 => \N__12677\,
            in2 => \N__13335\,
            in3 => \N__15222\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.un1_num_11_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18523\,
            in1 => \N__18481\,
            in2 => \N__18364\,
            in3 => \N__18395\,
            lcout => \Lab_UT.nine\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13713\,
            in2 => \_gnd_net_\,
            in3 => \N__13601\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__13326\,
            in1 => \N__13180\,
            in2 => \N__15042\,
            in3 => \N__13452\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22289\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.un1_num_7_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__13131\,
            in1 => \N__13061\,
            in2 => \N__13025\,
            in3 => \N__12957\,
            lcout => \Lab_UT.five\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__13448\,
            in1 => \N__12911\,
            in2 => \N__13334\,
            in3 => \N__15087\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_fast_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__13387\,
            in1 => \N__12887\,
            in2 => \N__12905\,
            in3 => \N__13220\,
            lcout => \Lab_UT.didp.q_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNI33OG1_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__20110\,
            in1 => \N__18938\,
            in2 => \N__20184\,
            in3 => \N__22736\,
            lcout => \Lab_UT.didp.countrce4.q_5_1\,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__13388\,
            in1 => \N__13215\,
            in2 => \N__12881\,
            in3 => \N__20178\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__13193\,
            in1 => \N__13390\,
            in2 => \N__13225\,
            in3 => \N__20242\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.un1_num_5_2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20177\,
            in2 => \_gnd_net_\,
            in3 => \N__20111\,
            lcout => OPEN,
            ltout => \Lab_UT.three_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__19856\,
            in1 => \N__18939\,
            in2 => \N__13238\,
            in3 => \N__20316\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__13389\,
            in1 => \N__20312\,
            in2 => \N__13235\,
            in3 => \N__13216\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22285\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_1_3_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20240\,
            in2 => \_gnd_net_\,
            in3 => \N__20173\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.reset_12_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16292\,
            in1 => \N__20109\,
            in2 => \N__13232\,
            in3 => \N__20311\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.reset_12_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13847\,
            in1 => \N__13359\,
            in2 => \N__13229\,
            in3 => \N__13817\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => 'H',
            sr => \N__21978\
        );

    \Lab_UT.didp.countrce4.q_RNIPP8Q_1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20172\,
            in1 => \N__20107\,
            in2 => \_gnd_net_\,
            in3 => \N__20310\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNIEP822_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__18934\,
            in1 => \N__19406\,
            in2 => \N__13196\,
            in3 => \N__20241\,
            lcout => \Lab_UT.didp.countrce4.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_0_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__16293\,
            in1 => \N__13846\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22280\,
            ce => 'H',
            sr => \N__21978\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100000101"
        )
    port map (
            in0 => \N__20108\,
            in1 => \_gnd_net_\,
            in2 => \N__18941\,
            in3 => \N__16488\,
            lcout => \Lab_UT.didp.countrce4.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13502\,
            in2 => \_gnd_net_\,
            in3 => \N__14945\,
            lcout => \oneSecStrb\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__21127\,
            in1 => \N__15352\,
            in2 => \N__20665\,
            in3 => \N__22039\,
            lcout => \Lab_UT.didp.regrce4.LdAMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.un26_ce_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__13842\,
            in1 => \N__13465\,
            in2 => \N__13820\,
            in3 => \N__18646\,
            lcout => \Lab_UT.didp.un26_ce_0\,
            ltout => \Lab_UT.didp.un26_ce_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_2_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__13466\,
            in1 => \_gnd_net_\,
            in2 => \N__13457\,
            in3 => \N__16316\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \N__21982\
        );

    \Lab_UT.didp.ce_RNO_0_3_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__18940\,
            in1 => \N__20654\,
            in2 => \N__15353\,
            in3 => \N__21128\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_3_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__16299\,
            in1 => \N__13360\,
            in2 => \N__13406\,
            in3 => \N__13403\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \N__21982\
        );

    \Lab_UT.didp.reset_2_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13845\,
            in1 => \N__13819\,
            in2 => \N__13364\,
            in3 => \N__16301\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \N__21982\
        );

    \Lab_UT.didp.ce_1_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__18647\,
            in1 => \N__16317\,
            in2 => \_gnd_net_\,
            in3 => \N__13843\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \N__21982\
        );

    \Lab_UT.didp.reset_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13844\,
            in1 => \N__13818\,
            in2 => \_gnd_net_\,
            in3 => \N__16300\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22276\,
            ce => 'H',
            sr => \N__21982\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13739\,
            in2 => \N__13724\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13691\,
            in2 => \_gnd_net_\,
            in3 => \N__13670\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13589\,
            in1 => \N__13667\,
            in2 => \_gnd_net_\,
            in3 => \N__13655\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__22272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13652\,
            in2 => \_gnd_net_\,
            in3 => \N__13631\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__13623\,
            in1 => \N__13588\,
            in2 => \N__13529\,
            in3 => \N__13532\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22272\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_19_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21126\,
            in1 => \N__15470\,
            in2 => \_gnd_net_\,
            in3 => \N__13853\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_2_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__21452\,
            in1 => \N__20663\,
            in2 => \N__13511\,
            in3 => \N__15497\,
            lcout => \Lab_UT.dictrl.N_11_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_1_3_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__13898\,
            in1 => \N__15518\,
            in2 => \N__13886\,
            in3 => \N__15487\,
            lcout => \Lab_UT.dictrl.g0_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13875\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22270\,
            ce => \N__22071\,
            sr => \N__22005\
        );

    \buart.Z_rx.shifter_fast_7_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22270\,
            ce => \N__22071\,
            sr => \N__22005\
        );

    \buart.Z_rx.shifter_7_rep1_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13876\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22270\,
            ce => \N__22071\,
            sr => \N__22005\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_22_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__23033\,
            in1 => \N__22876\,
            in2 => \N__16874\,
            in3 => \N__22558\,
            lcout => \Lab_UT.dictrl.g2_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22727\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__22069\,
            sr => \N__22006\
        );

    \buart.Z_rx.shifter_1_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19832\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__22069\,
            sr => \N__22006\
        );

    \buart.Z_rx.shifter_fast_4_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22559\,
            lcout => bu_rx_data_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22269\,
            ce => \N__22069\,
            sr => \N__22006\
        );

    \uu2.w_addr_user_5_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13933\,
            in1 => \N__14122\,
            in2 => \N__14182\,
            in3 => \N__14207\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__14054\
        );

    \uu2.w_addr_user_4_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__14121\,
            in1 => \N__13932\,
            in2 => \_gnd_net_\,
            in3 => \N__14173\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__14054\
        );

    \uu2.w_addr_user_6_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__13934\,
            in1 => \N__14123\,
            in2 => \N__14141\,
            in3 => \N__14492\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__14054\
        );

    \uu2.w_addr_user_RNI93NG7_2_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__13948\,
            in1 => \N__15994\,
            in2 => \_gnd_net_\,
            in3 => \N__13955\,
            lcout => \uu2.un28_w_addr_user_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un20_w_addr_user_1_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__13982\,
            in1 => \N__15854\,
            in2 => \N__13973\,
            in3 => \N__17086\,
            lcout => \uu2.un20_w_addr_userZ0Z_1\,
            ltout => \uu2.un20_w_addr_userZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI43E87_2_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13949\,
            in2 => \N__13940\,
            in3 => \N__14723\,
            lcout => \uu2.w_addr_user_RNI43E87Z0Z_2\,
            ltout => \uu2.w_addr_user_RNI43E87Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNID65PE_2_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13937\,
            in3 => \N__13928\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_0_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14384\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__14047\
        );

    \uu2.w_addr_user_1_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__14385\,
            in1 => \N__14290\,
            in2 => \_gnd_net_\,
            in3 => \N__13930\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__14047\
        );

    \uu2.w_addr_user_2_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__13931\,
            in1 => \N__14339\,
            in2 => \N__14301\,
            in3 => \N__14386\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_0C_net\,
            ce => 'H',
            sr => \N__14047\
        );

    \uu2.w_addr_user_nesr_RNI1VU6_3_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14208\,
            in1 => \N__14234\,
            in2 => \N__14464\,
            in3 => \N__14368\,
            lcout => \uu2.un3_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__14369\,
            in1 => \N__14340\,
            in2 => \N__14244\,
            in3 => \N__14294\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__14069\,
            sr => \N__14046\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14181\,
            lcout => \uu2.un426_ci_3\,
            ltout => \uu2.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_7_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__14119\,
            in1 => \N__14459\,
            in2 => \N__14144\,
            in3 => \N__14497\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__14069\,
            sr => \N__14046\
        );

    \uu2.w_addr_user_nesr_8_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__14134\,
            in1 => \N__14120\,
            in2 => \N__14090\,
            in3 => \N__14441\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__14069\,
            sr => \N__14046\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__15679\,
            in1 => \N__15986\,
            in2 => \N__14498\,
            in3 => \N__15826\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011110000"
        )
    port map (
            in0 => \N__15827\,
            in1 => \N__14460\,
            in2 => \N__16972\,
            in3 => \N__15985\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_52_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__17256\,
            in1 => \N__16957\,
            in2 => \N__15685\,
            in3 => \N__16115\,
            lcout => \uu2.mem0.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI90ME1_5_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__16114\,
            in1 => \N__15678\,
            in2 => \N__16971\,
            in3 => \N__17257\,
            lcout => \uu2.bitmap_pmux_sn_N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_8_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__15680\,
            in1 => \N__16961\,
            in2 => \N__15718\,
            in3 => \N__16116\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_8C_net\,
            ce => \N__15611\,
            sr => \N__21947\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14496\,
            in1 => \_gnd_net_\,
            in2 => \N__14465\,
            in3 => \_gnd_net_\,
            lcout => \uu2.vbuf_w_addr_user.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNILN731_40_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001100101011101"
        )
    port map (
            in0 => \N__16113\,
            in1 => \N__16042\,
            in2 => \N__14978\,
            in3 => \N__14435\,
            lcout => \uu2.bitmap_pmux_26_bm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20052\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__21945\
        );

    \uu2.bitmap_52_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20053\,
            in1 => \_gnd_net_\,
            in2 => \N__14429\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_40C_net\,
            ce => 'H',
            sr => \N__21945\
        );

    \uu2.w_addr_displaying_RNIBICU6_2_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111010101"
        )
    port map (
            in0 => \N__14411\,
            in1 => \N__16055\,
            in2 => \N__14420\,
            in3 => \N__14816\,
            lcout => \uu2.w_addr_displaying_RNIBICU6Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNIF31A1_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000101010"
        )
    port map (
            in0 => \N__17615\,
            in1 => \N__17762\,
            in2 => \N__16126\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => \uu2.bitmap_pmux_sn_N_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIBICU6_0_2_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__14410\,
            in1 => \N__14815\,
            in2 => \N__14402\,
            in3 => \N__16054\,
            lcout => \uu2.w_addr_displaying_RNIBICU6_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIL1MV_52_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16109\,
            in1 => \N__14399\,
            in2 => \_gnd_net_\,
            in3 => \N__14393\,
            lcout => OPEN,
            ltout => \uu2.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_RNICS7L2_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__17629\,
            in1 => \N__16949\,
            in2 => \N__14819\,
            in3 => \N__16001\,
            lcout => \uu2.w_addr_displaying_3_rep1_nesr_RNICS7LZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__14807\,
            in1 => \N__14801\,
            in2 => \_gnd_net_\,
            in3 => \N__14714\,
            lcout => \Lab_UT.dictrl.un1_next_alarmstate21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.sec1_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14759\,
            lcout => \Lab_UT.sec1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI34K17_5_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14713\,
            in2 => \_gnd_net_\,
            in3 => \N__17281\,
            lcout => \uu2.N_31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__14589\,
            in1 => \N__14653\,
            in2 => \_gnd_net_\,
            in3 => \N__14556\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__14557\,
            in1 => \N__14591\,
            in2 => \N__14657\,
            in3 => \N__14638\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14634\,
            in2 => \_gnd_net_\,
            in3 => \N__14651\,
            lcout => \resetGen.un241_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__14652\,
            in1 => \_gnd_net_\,
            in2 => \N__14639\,
            in3 => \N__14620\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011100"
        )
    port map (
            in0 => \N__14590\,
            in1 => \N__14512\,
            in2 => \N__14561\,
            in3 => \N__14558\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18560\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \uu2.bitmap_180_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14954\,
            in2 => \_gnd_net_\,
            in3 => \N__20022\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \uu2.bitmap_111_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14946\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \uu2.vram_rd_clk_det_0_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14881\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \uu2.vram_rd_clk_det_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14845\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \uu2.bitmap_221_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18599\,
            in2 => \_gnd_net_\,
            in3 => \N__20023\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__21941\
        );

    \Lab_UT.bcd2segment3.segment_0_2_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__15217\,
            in1 => \N__15163\,
            in2 => \N__15112\,
            in3 => \N__15024\,
            lcout => \Lab_UT.bcd2segment3.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_4_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__15158\,
            in1 => \N__15027\,
            in2 => \N__15115\,
            in3 => \N__15212\,
            lcout => \Lab_UT.bcd2segment3.segmentUQ_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_5_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111000010"
        )
    port map (
            in0 => \N__15213\,
            in1 => \N__15159\,
            in2 => \N__15111\,
            in3 => \N__15023\,
            lcout => \Lab_UT.bcd2segment3.segmentUQ_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_6_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100111100001"
        )
    port map (
            in0 => \N__15160\,
            in1 => \N__15026\,
            in2 => \N__15114\,
            in3 => \N__15214\,
            lcout => \Lab_UT.bcd2segment3.segmentUQ_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segment_0_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101111001"
        )
    port map (
            in0 => \N__15215\,
            in1 => \N__15161\,
            in2 => \N__15110\,
            in3 => \N__15022\,
            lcout => \Lab_UT.bcd2segment3.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segment_0_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__15162\,
            in1 => \N__15028\,
            in2 => \N__15116\,
            in3 => \N__15216\,
            lcout => \Lab_UT.bcd2segment3.segment_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100110"
        )
    port map (
            in0 => \N__15218\,
            in1 => \N__15164\,
            in2 => \N__15113\,
            in3 => \N__15025\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14981\,
            in3 => \N__19981\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__21938\
        );

    \Lab_UT.didp.countrce1.q_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__18464\,
            in1 => \N__16249\,
            in2 => \N__15287\,
            in3 => \N__15307\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__15263\,
            in1 => \N__16490\,
            in2 => \_gnd_net_\,
            in3 => \N__18347\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__18348\,
            in1 => \N__15306\,
            in2 => \N__14963\,
            in3 => \N__16248\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__18525\,
            in1 => \N__14960\,
            in2 => \N__15269\,
            in3 => \N__19873\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__18526\,
            in1 => \N__16250\,
            in2 => \N__15314\,
            in3 => \N__15308\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18524\,
            in1 => \N__18463\,
            in2 => \_gnd_net_\,
            in3 => \N__18346\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__19412\,
            in2 => \N__15311\,
            in3 => \N__18396\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__15305\,
            in1 => \N__18397\,
            in2 => \N__15290\,
            in3 => \N__16247\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22301\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__22760\,
            in1 => \N__18465\,
            in2 => \N__15268\,
            in3 => \N__18345\,
            lcout => \Lab_UT.didp.countrce1.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001100"
        )
    port map (
            in0 => \N__19411\,
            in1 => \N__18617\,
            in2 => \N__19879\,
            in3 => \N__22759\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_0_a3_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__19138\,
            in1 => \N__16517\,
            in2 => \N__15275\,
            in3 => \N__19177\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_0_a3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001010000"
        )
    port map (
            in0 => \N__19018\,
            in1 => \N__16508\,
            in2 => \N__15272\,
            in3 => \N__15320\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22294\,
            ce => 'H',
            sr => \N__21979\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_8_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__21753\,
            in1 => \N__21465\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_i_a3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_5_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19176\,
            in1 => \N__23210\,
            in2 => \N__15242\,
            in3 => \N__19137\,
            lcout => \Lab_UT.dictrl.N_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15392\,
            in2 => \_gnd_net_\,
            in3 => \N__19017\,
            lcout => \Lab_UT.dicLdSones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22294\,
            ce => 'H',
            sr => \N__21979\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_6_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21063\,
            in1 => \N__21468\,
            in2 => \_gnd_net_\,
            in3 => \N__20828\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_i_a3_0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_4_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__22743\,
            in1 => \N__19880\,
            in2 => \N__15338\,
            in3 => \N__19389\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_i_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_0_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__16523\,
            in1 => \N__19140\,
            in2 => \N__15335\,
            in3 => \N__19175\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_i_a3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000111"
        )
    port map (
            in0 => \N__15329\,
            in1 => \N__16397\,
            in2 => \N__15332\,
            in3 => \N__19022\,
            lcout => \Lab_UT.LdSones_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22288\,
            ce => 'H',
            sr => \N__21983\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__21717\,
            in1 => \N__20829\,
            in2 => \N__20664\,
            in3 => \N__21469\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g3_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21202\,
            in2 => \_gnd_net_\,
            in3 => \N__21062\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_7_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__20395\,
            in1 => \N__21467\,
            in2 => \N__15323\,
            in3 => \N__23222\,
            lcout => \Lab_UT.dictrl.i6_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__21470\,
            in1 => \N__20649\,
            in2 => \N__20854\,
            in3 => \N__21718\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_RNIOF67_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21124\,
            in1 => \N__21427\,
            in2 => \N__21752\,
            in3 => \N__21212\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__20853\,
            in1 => \N__15410\,
            in2 => \N__21763\,
            in3 => \N__15401\,
            lcout => \Lab_UT.dictrl.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22283\,
            ce => 'H',
            sr => \N__21986\
        );

    \Lab_UT.dictrl.g0_1_0_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22974\,
            in1 => \N__19504\,
            in2 => \N__20903\,
            in3 => \N__21572\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_8_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111011101"
        )
    port map (
            in0 => \N__20519\,
            in1 => \N__21125\,
            in2 => \N__15416\,
            in3 => \N__19092\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_29_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_6_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__21428\,
            in1 => \N__21211\,
            in2 => \N__15413\,
            in3 => \N__15461\,
            lcout => \Lab_UT.dictrl.N_30_0\,
            ltout => \Lab_UT.dictrl.N_30_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNI6JM59_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__21711\,
            in1 => \N__20850\,
            in2 => \N__15404\,
            in3 => \N__15400\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_2\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_RNO_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__20851\,
            in1 => \N__21712\,
            in2 => \N__15383\,
            in3 => \N__18875\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.dicLdAMones_0_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__21713\,
            in1 => \N__20852\,
            in2 => \N__15380\,
            in3 => \N__18831\,
            lcout => \Lab_UT.dicLdAMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22283\,
            ce => 'H',
            sr => \N__21986\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_13_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__22531\,
            in1 => \N__19460\,
            in2 => \N__15362\,
            in3 => \N__19256\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111001110"
        )
    port map (
            in0 => \N__23209\,
            in1 => \N__21109\,
            in2 => \N__15500\,
            in3 => \N__16727\,
            lcout => \Lab_UT.dictrl.N_7_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_5_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__16664\,
            in1 => \N__19592\,
            in2 => \N__15527\,
            in3 => \N__19541\,
            lcout => \Lab_UT.dictrl.g2_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_1_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19540\,
            in1 => \N__16663\,
            in2 => \N__15491\,
            in3 => \N__16711\,
            lcout => \Lab_UT.dictrl.g0_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_4_2_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__19593\,
            in2 => \N__16670\,
            in3 => \N__19542\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_4Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_10_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__21569\,
            in1 => \N__20494\,
            in2 => \N__15473\,
            in3 => \N__22969\,
            lcout => \Lab_UT.dictrl.next_state18_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011111"
        )
    port map (
            in0 => \N__22970\,
            in1 => \_gnd_net_\,
            in2 => \N__20498\,
            in3 => \N__21570\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111111111111"
        )
    port map (
            in0 => \N__18890\,
            in1 => \N__22532\,
            in2 => \N__15464\,
            in3 => \N__21110\,
            lcout => \Lab_UT.dictrl.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_2_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19545\,
            in1 => \N__16659\,
            in2 => \N__19600\,
            in3 => \N__16715\,
            lcout => \Lab_UT.dictrl.next_state12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_1_2_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__16714\,
            in1 => \N__19588\,
            in2 => \N__16668\,
            in3 => \N__19544\,
            lcout => \Lab_UT.dictrl.g2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state32_4_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19543\,
            in1 => \N__16655\,
            in2 => \N__19599\,
            in3 => \N__16713\,
            lcout => \Lab_UT.dictrl.next_state32Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_5_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__22870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22274\,
            ce => \N__22068\,
            sr => \N__22007\
        );

    \buart.Z_rx.shifter_5_rep1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22869\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22274\,
            ce => \N__22068\,
            sr => \N__22007\
        );

    \buart.Z_rx.shifter_4_rep1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22545\,
            lcout => bu_rx_data_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22274\,
            ce => \N__22068\,
            sr => \N__22007\
        );

    \buart.Z_rx.shifter_6_rep1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23034\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22271\,
            ce => \N__22067\,
            sr => \N__22008\
        );

    \buart.Z_rx.shifter_fast_3_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22458\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22271\,
            ce => \N__22067\,
            sr => \N__22008\
        );

    \uu2.mem0.ram512X8_inst_RNO_45_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17507\,
            in1 => \N__17888\,
            in2 => \_gnd_net_\,
            in3 => \N__17631\,
            lcout => \uu2.mem0.G_11_0_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_53_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17506\,
            in2 => \_gnd_net_\,
            in3 => \N__17758\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_98_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_46_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17990\,
            in1 => \N__17632\,
            in2 => \N__15512\,
            in3 => \N__17551\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_30_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__15509\,
            in1 => \N__17202\,
            in2 => \N__15503\,
            in3 => \N__17420\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_20_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15587\,
            in1 => \N__17119\,
            in2 => \N__15578\,
            in3 => \N__16785\,
            lcout => \uu2.mem0.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_23_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15671\,
            in1 => \N__16962\,
            in2 => \N__18117\,
            in3 => \N__16119\,
            lcout => \uu2.mem0.G_11_0_0_a2_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_28_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__16120\,
            in1 => \_gnd_net_\,
            in2 => \N__16973\,
            in3 => \_gnd_net_\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI31F32_34_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011111010"
        )
    port map (
            in0 => \N__19922\,
            in1 => \N__19673\,
            in2 => \N__17633\,
            in3 => \N__15575\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNI31F32Z0Z_34_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNII6975_34_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15533\,
            in2 => \N__15569\,
            in3 => \N__15539\,
            lcout => OPEN,
            ltout => \uu2.N_401_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI8B24J_34_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15566\,
            in2 => \N__15560\,
            in3 => \N__15557\,
            lcout => \uu2.N_406\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIJS4P_162_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__16041\,
            in1 => \N__16190\,
            in2 => \_gnd_net_\,
            in3 => \N__19664\,
            lcout => OPEN,
            ltout => \uu2.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI2Q8F1_111_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__15551\,
            in1 => \_gnd_net_\,
            in2 => \N__15542\,
            in3 => \N__15623\,
            lcout => \uu2.bitmap_RNI2Q8F1Z0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNIDBHK1_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110110"
        )
    port map (
            in0 => \N__17741\,
            in1 => \N__17541\,
            in2 => \N__17630\,
            in3 => \N__16950\,
            lcout => \uu2.bitmap_pmux_sn_N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__15617\,
            in1 => \N__16040\,
            in2 => \_gnd_net_\,
            in3 => \N__17332\,
            lcout => \uu2.bitmap_pmux_sn_N_54_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_nesr_3_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__17205\,
            in2 => \N__16046\,
            in3 => \N__17884\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__17203\,
            in1 => \N__17628\,
            in2 => \N__17910\,
            in3 => \N__17390\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.w_addr_displaying_nesr_1_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__17988\,
            in1 => \_gnd_net_\,
            in2 => \N__17764\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17750\,
            in2 => \_gnd_net_\,
            in3 => \N__17986\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.w_addr_displaying_nesr_3_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__17204\,
            in1 => \N__18072\,
            in2 => \N__17911\,
            in3 => \N__17391\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.w_addr_displaying_fast_nesr_1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__17987\,
            in1 => \_gnd_net_\,
            in2 => \N__17763\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_3C_net\,
            ce => \N__15607\,
            sr => \N__21948\
        );

    \uu2.bitmap_RNIFH0N_90_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__18308\,
            in1 => \N__18179\,
            in2 => \N__18236\,
            in3 => \N__15593\,
            lcout => \uu2.bitmap_pmux_19_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_90_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18587\,
            in2 => \_gnd_net_\,
            in3 => \N__20021\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__21946\
        );

    \uu2.bitmap_186_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18578\,
            in2 => \_gnd_net_\,
            in3 => \N__20019\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__21946\
        );

    \uu2.bitmap_RNIKGSI_58_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16169\,
            in1 => \N__18180\,
            in2 => \_gnd_net_\,
            in3 => \N__16133\,
            lcout => OPEN,
            ltout => \uu2.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI04AD1_314_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16125\,
            in2 => \N__16058\,
            in3 => \N__16010\,
            lcout => \uu2.bitmap_RNI04AD1Z0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_314_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20020\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18608\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__21946\
        );

    \uu2.bitmap_RNICM7R_180_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__16039\,
            in1 => \N__16016\,
            in2 => \_gnd_net_\,
            in3 => \N__16009\,
            lcout => \uu2.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_7_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__17297\,
            in1 => \N__15657\,
            in2 => \N__18188\,
            in3 => \N__15724\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_7C_net\,
            ce => 'H',
            sr => \N__21944\
        );

    \uu2.w_addr_displaying_7_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001111000"
        )
    port map (
            in0 => \N__17296\,
            in1 => \N__15656\,
            in2 => \N__16966\,
            in3 => \N__15723\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_7C_net\,
            ce => 'H',
            sr => \N__21944\
        );

    \uu2.w_addr_displaying_RNIVAPV6_5_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011101"
        )
    port map (
            in0 => \N__15929\,
            in1 => \N__15754\,
            in2 => \N__15725\,
            in3 => \N__15855\,
            lcout => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5\,
            ltout => \uu2.w_addr_displaying_RNIVAPV6Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_6_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111110110000"
        )
    port map (
            in0 => \N__15755\,
            in1 => \N__15722\,
            in2 => \N__15692\,
            in3 => \N__15658\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_7C_net\,
            ce => 'H',
            sr => \N__21944\
        );

    \uu2.bitmap_203_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16208\,
            in2 => \_gnd_net_\,
            in3 => \N__19976\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \uu2.bitmap_200_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__19975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16202\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \uu2.bitmap_168_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16196\,
            in2 => \_gnd_net_\,
            in3 => \N__19974\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \uu2.bitmap_75_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19979\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16181\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \uu2.bitmap_72_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16175\,
            in2 => \_gnd_net_\,
            in3 => \N__19978\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \uu2.bitmap_58_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18566\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__21939\
        );

    \Lab_UT.dictrl.state_ret_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101110101111"
        )
    port map (
            in0 => \N__20848\,
            in1 => \N__21269\,
            in2 => \N__19043\,
            in3 => \N__21740\,
            lcout => \Lab_UT.state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22310\,
            ce => 'H',
            sr => \N__21980\
        );

    \Lab_UT.dictrl.state_ret_5_RNIIMGL_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__21738\,
            in1 => \N__18805\,
            in2 => \_gnd_net_\,
            in3 => \N__23181\,
            lcout => \Lab_UT.LdASones\,
            ltout => \Lab_UT.LdASones_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNO_0_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16148\,
            in3 => \N__16145\,
            lcout => \Lab_UT.didp.ce_9_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_RNI0TGF_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18670\,
            in2 => \_gnd_net_\,
            in3 => \N__20606\,
            lcout => \Lab_UT.dicRun_2\,
            ltout => \Lab_UT.dicRun_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__18806\,
            in1 => \N__16355\,
            in2 => \N__16349\,
            in3 => \N__16334\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22310\,
            ce => 'H',
            sr => \N__21980\
        );

    \Lab_UT.dictrl.state_ret_1_RNIKRKU_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__20605\,
            in2 => \_gnd_net_\,
            in3 => \N__18669\,
            lcout => \Lab_UT.Run\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010111010111111"
        )
    port map (
            in0 => \N__20849\,
            in1 => \N__21739\,
            in2 => \N__20534\,
            in3 => \N__16538\,
            lcout => \Lab_UT.dictrl.state_i_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22310\,
            ce => 'H',
            sr => \N__21980\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_3_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__19352\,
            in1 => \N__22765\,
            in2 => \N__19871\,
            in3 => \N__16220\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_i_a3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__16214\,
            in1 => \N__16229\,
            in2 => \N__16223\,
            in3 => \N__18772\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__20811\,
            in1 => \N__18878\,
            in2 => \N__21794\,
            in3 => \N__18838\,
            lcout => \Lab_UT.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22302\,
            ce => 'H',
            sr => \N__21984\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_7_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20795\,
            in1 => \N__21064\,
            in2 => \_gnd_net_\,
            in3 => \N__16593\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_4_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21784\,
            in1 => \N__21369\,
            in2 => \_gnd_net_\,
            in3 => \N__23203\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_3_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__23204\,
            in1 => \N__21786\,
            in2 => \_gnd_net_\,
            in3 => \N__16594\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__21785\,
            in2 => \_gnd_net_\,
            in3 => \N__16595\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110110001"
        )
    port map (
            in0 => \N__21060\,
            in1 => \N__19201\,
            in2 => \N__16622\,
            in3 => \N__18773\,
            lcout => \Lab_UT.dictrl.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_7_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20817\,
            in1 => \N__21059\,
            in2 => \_gnd_net_\,
            in3 => \N__16591\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_0_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__19338\,
            in1 => \N__19833\,
            in2 => \N__16496\,
            in3 => \N__22741\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__16751\,
            in2 => \N__22875\,
            in3 => \N__16482\,
            lcout => \Lab_UT.dictrl.next_alarmstateZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m4_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23192\,
            in2 => \_gnd_net_\,
            in3 => \N__20394\,
            lcout => \Lab_UT.dictrl.N_5\,
            ltout => \Lab_UT.dictrl.N_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000110011"
        )
    port map (
            in0 => \N__16604\,
            in1 => \N__19200\,
            in2 => \N__16400\,
            in3 => \N__21061\,
            lcout => \Lab_UT.dictrl.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_5_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16610\,
            in1 => \N__19139\,
            in2 => \N__19178\,
            in3 => \N__23193\,
            lcout => \Lab_UT.dictrl.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_5_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__22742\,
            in1 => \N__19339\,
            in2 => \N__19870\,
            in3 => \N__16592\,
            lcout => \Lab_UT.dictrl.g0_0_0_o4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__19503\,
            in1 => \N__16860\,
            in2 => \N__22975\,
            in3 => \N__16576\,
            lcout => \Lab_UT.dictrl.next_state18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_11_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111110"
        )
    port map (
            in0 => \N__21209\,
            in1 => \N__19184\,
            in2 => \N__21485\,
            in3 => \N__16681\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_10_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100111"
        )
    port map (
            in0 => \N__21111\,
            in1 => \N__16556\,
            in2 => \N__16613\,
            in3 => \N__18770\,
            lcout => \Lab_UT.dictrl.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_8_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21693\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_RNO_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__22747\,
            in1 => \N__19364\,
            in2 => \N__19855\,
            in3 => \N__16578\,
            lcout => \Lab_UT.dictrl.g0_0_i_o4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_4_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__16577\,
            in1 => \N__21555\,
            in2 => \N__20493\,
            in3 => \N__22965\,
            lcout => \Lab_UT.dictrl.next_state18_0\,
            ltout => \Lab_UT.dictrl.next_state18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_3_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__16682\,
            in1 => \_gnd_net_\,
            in2 => \N__16550\,
            in3 => \N__21112\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_9_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__21432\,
            in1 => \N__20645\,
            in2 => \N__16547\,
            in3 => \N__16544\,
            lcout => \Lab_UT.dictrl.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__21530\,
            in1 => \N__20460\,
            in2 => \N__22971\,
            in3 => \N__16529\,
            lcout => \Lab_UT.dictrl.g2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__19707\,
            in1 => \N__19453\,
            in2 => \_gnd_net_\,
            in3 => \N__19249\,
            lcout => \Lab_UT.dictrl.gZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_3_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16862\,
            in1 => \N__22455\,
            in2 => \N__19505\,
            in3 => \N__19556\,
            lcout => \Lab_UT.dictrl.next_alarmstate4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__19708\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16716\,
            lcout => \Lab_UT.dictrl.next_alarmstate4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_0_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__16742\,
            in1 => \N__22952\,
            in2 => \N__21554\,
            in3 => \N__20461\,
            lcout => \Lab_UT.dictrl.g2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_3_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__16669\,
            in1 => \N__16861\,
            in2 => \N__19712\,
            in3 => \N__16717\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_1_0_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000110101011"
        )
    port map (
            in0 => \N__21108\,
            in1 => \N__19511\,
            in2 => \N__16736\,
            in3 => \N__16733\,
            lcout => \Lab_UT.dictrl.g0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_6_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__19452\,
            in1 => \N__19594\,
            in2 => \N__19699\,
            in3 => \N__19248\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_5_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23046\,
            in1 => \N__22865\,
            in2 => \N__16721\,
            in3 => \N__16718\,
            lcout => \Lab_UT.dictrl.next_state12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_8_3_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__19451\,
            in1 => \N__16654\,
            in2 => \N__19698\,
            in3 => \N__19247\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_8_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__23045\,
            in1 => \N__22430\,
            in2 => \N__16877\,
            in3 => \N__22544\,
            lcout => \Lab_UT.dictrl.next_state12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_1_3_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__19694\,
            in1 => \N__16859\,
            in2 => \N__19499\,
            in3 => \N__19595\,
            lcout => \Lab_UT.dictrl.g2_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19780\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22275\,
            ce => \N__22070\,
            sr => \N__22009\
        );

    \buart.Z_rx.shifter_3_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22457\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22275\,
            ce => \N__22070\,
            sr => \N__22009\
        );

    \uu2.mem0.ram512X8_inst_RNO_18_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16838\,
            in1 => \N__16810\,
            in2 => \N__17120\,
            in3 => \N__17570\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16832\,
            in1 => \N__17057\,
            in2 => \N__16826\,
            in3 => \N__16766\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17757\,
            in2 => \_gnd_net_\,
            in3 => \N__17989\,
            lcout => \uu2.N_30_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_32_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110110110100"
        )
    port map (
            in0 => \N__17514\,
            in1 => \N__18102\,
            in2 => \N__17207\,
            in3 => \N__17419\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_24_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_22_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16811\,
            in1 => \N__17118\,
            in2 => \N__16790\,
            in3 => \N__16786\,
            lcout => \uu2.mem0.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_24_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17513\,
            in1 => \N__17261\,
            in2 => \N__17206\,
            in3 => \N__18288\,
            lcout => OPEN,
            ltout => \uu2.mem0.G_11_0_0_a2_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__17126\,
            in1 => \N__17117\,
            in2 => \N__17093\,
            in3 => \N__17090\,
            lcout => \uu2.mem0.G_11_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17051\,
            in2 => \_gnd_net_\,
            in3 => \N__20057\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__21952\
        );

    \uu2.bitmap_84_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17039\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__21952\
        );

    \uu2.bitmap_212_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17027\,
            in2 => \_gnd_net_\,
            in3 => \N__20054\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__21952\
        );

    \uu2.bitmap_215_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20055\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17015\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__21952\
        );

    \uu2.bitmap_RNIOPSS_212_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__17003\,
            in1 => \N__18187\,
            in2 => \N__16997\,
            in3 => \N__18226\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_17_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIEMII1_84_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__16988\,
            in1 => \N__16982\,
            in2 => \N__16976\,
            in3 => \N__16967\,
            lcout => \uu2.N_104\,
            ltout => \uu2.N_104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_38_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__18284\,
            in1 => \N__17627\,
            in2 => \N__17576\,
            in3 => \N__17681\,
            lcout => OPEN,
            ltout => \uu2.mem0.G_11_0_0_a3_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_27_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__17435\,
            in1 => \N__17564\,
            in2 => \N__17573\,
            in3 => \N__18260\,
            lcout => \uu2.mem0.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_40_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000100001"
        )
    port map (
            in0 => \N__17387\,
            in1 => \N__17545\,
            in2 => \N__17889\,
            in3 => \N__17515\,
            lcout => \uu2.mem0.N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__17547\,
            in1 => \N__17303\,
            in2 => \N__17418\,
            in3 => \N__17865\,
            lcout => \uu2.w_addr_displaying_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__21950\
        );

    \uu2.mem0.ram512X8_inst_RNO_41_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010001000010"
        )
    port map (
            in0 => \N__17749\,
            in1 => \N__17546\,
            in2 => \N__17890\,
            in3 => \N__17516\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17864\,
            in2 => \_gnd_net_\,
            in3 => \N__17298\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__21950\
        );

    \uu2.w_addr_displaying_fast_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__17388\,
            in1 => \N__17880\,
            in2 => \N__17315\,
            in3 => \N__17333\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__21950\
        );

    \uu2.w_addr_displaying_fast_0_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17302\,
            in2 => \_gnd_net_\,
            in3 => \N__18235\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__21950\
        );

    \uu2.w_addr_displaying_0_rep1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__17977\,
            in1 => \_gnd_net_\,
            in2 => \N__17314\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__21950\
        );

    \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_0_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17748\,
            in2 => \_gnd_net_\,
            in3 => \N__17976\,
            lcout => \uu2.N_30_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_194_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19646\,
            in2 => \_gnd_net_\,
            in3 => \N__20030\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__21949\
        );

    \uu2.bitmap_66_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__20032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19637\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__21949\
        );

    \uu2.bitmap_RNILQ2M_66_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__18241\,
            in1 => \N__18183\,
            in2 => \N__17699\,
            in3 => \N__17690\,
            lcout => \uu2.bitmap_pmux_20_ns_1\,
            ltout => \uu2.bitmap_pmux_20_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_48_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__17662\,
            in1 => \N__17671\,
            in2 => \N__17684\,
            in3 => \N__17985\,
            lcout => \uu2.mem0.N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_197_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__19655\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20031\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__21949\
        );

    \uu2.bitmap_69_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20033\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20354\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_194C_net\,
            ce => 'H',
            sr => \N__21949\
        );

    \uu2.mem0.ram512X8_inst_RNO_33_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__17672\,
            in1 => \N__17663\,
            in2 => \N__17904\,
            in3 => \N__17654\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_108_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_25_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__18025\,
            in1 => \N__17771\,
            in2 => \N__17648\,
            in3 => \N__17999\,
            lcout => \uu2.mem0.N_404_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_55_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__18182\,
            in1 => \N__18251\,
            in2 => \N__18242\,
            in3 => \N__18196\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_16_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_49_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__18145\,
            in1 => \N__18130\,
            in2 => \N__18299\,
            in3 => \N__17991\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_39_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__18292\,
            in1 => \N__18114\,
            in2 => \N__18263\,
            in3 => \N__17936\,
            lcout => \uu2.mem0.G_11_0_0_a3_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_54_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__18250\,
            in1 => \N__18237\,
            in2 => \N__18200\,
            in3 => \N__18181\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_16_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_47_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__17992\,
            in1 => \N__18146\,
            in2 => \N__18134\,
            in3 => \N__18131\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_22_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_35_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__18115\,
            in1 => \N__18026\,
            in2 => \N__18011\,
            in3 => \N__18008\,
            lcout => \uu2.mem0.bitmap_pmux_27_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_50_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__17800\,
            in2 => \N__17786\,
            in3 => \N__17929\,
            lcout => \uu2.mem0.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_34_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110010001"
        )
    port map (
            in0 => \N__17930\,
            in1 => \N__17903\,
            in2 => \N__17804\,
            in3 => \N__17785\,
            lcout => \uu2.mem0.N_109_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111100010"
        )
    port map (
            in0 => \N__18546\,
            in1 => \N__18482\,
            in2 => \N__18429\,
            in3 => \N__18369\,
            lcout => \Lab_UT.bcd2segment1.segmentUQ_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_0_2_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__18366\,
            in1 => \N__18414\,
            in2 => \N__18497\,
            in3 => \N__18543\,
            lcout => \Lab_UT.bcd2segment1.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_5_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111100100"
        )
    port map (
            in0 => \N__18545\,
            in1 => \N__18483\,
            in2 => \N__18428\,
            in3 => \N__18368\,
            lcout => \Lab_UT.bcd2segment1.segmentUQ_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_6_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011000011"
        )
    port map (
            in0 => \N__18365\,
            in1 => \N__18413\,
            in2 => \N__18495\,
            in3 => \N__18542\,
            lcout => \Lab_UT.bcd2segment1.segmentUQ_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_0_0_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__18547\,
            in1 => \N__18487\,
            in2 => \N__18430\,
            in3 => \N__18370\,
            lcout => \Lab_UT.bcd2segment1.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_0_1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__18367\,
            in1 => \N__18415\,
            in2 => \N__18496\,
            in3 => \N__18544\,
            lcout => \Lab_UT.bcd2segment1.segment_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_4_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__18548\,
            in1 => \N__18494\,
            in2 => \N__18431\,
            in3 => \N__18371\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_218_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18311\,
            in3 => \N__19980\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_218C_net\,
            ce => 'H',
            sr => \N__21942\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_6_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18968\,
            in1 => \N__21374\,
            in2 => \_gnd_net_\,
            in3 => \N__20951\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__21376\,
            in1 => \N__19208\,
            in2 => \N__18734\,
            in3 => \N__21073\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100010011"
        )
    port map (
            in0 => \N__20741\,
            in1 => \N__18731\,
            in2 => \N__18725\,
            in3 => \N__19013\,
            lcout => \Lab_UT.LdStens_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__21985\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m33_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000001100"
        )
    port map (
            in0 => \N__20952\,
            in1 => \N__20608\,
            in2 => \N__21423\,
            in3 => \N__18969\,
            lcout => \Lab_UT.dictrl.N_39_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_6_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18967\,
            in1 => \N__21373\,
            in2 => \_gnd_net_\,
            in3 => \N__20950\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_2_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__21375\,
            in1 => \N__19207\,
            in2 => \N__18722\,
            in3 => \N__21072\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__20876\,
            in1 => \N__18743\,
            in2 => \N__18719\,
            in3 => \N__19012\,
            lcout => \Lab_UT.LdStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22319\,
            ce => 'H',
            sr => \N__21985\
        );

    \Lab_UT.didp.ce_10_1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001110000"
        )
    port map (
            in0 => \N__20728\,
            in1 => \N__18671\,
            in2 => \N__18656\,
            in3 => \N__20607\,
            lcout => \Lab_UT.didp.ce_10_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m27_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100000010000"
        )
    port map (
            in0 => \N__21067\,
            in1 => \N__21448\,
            in2 => \N__21236\,
            in3 => \N__18632\,
            lcout => \Lab_UT.dictrl.i6_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_9_RNO_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__21446\,
            in1 => \N__20796\,
            in2 => \_gnd_net_\,
            in3 => \N__21065\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m18_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110110101111"
        )
    port map (
            in0 => \N__21066\,
            in1 => \N__18769\,
            in2 => \N__21235\,
            in3 => \N__21601\,
            lcout => \Lab_UT.dictrl.N_19\,
            ltout => \Lab_UT.dictrl.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNICIPPD_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100100010"
        )
    port map (
            in0 => \N__21447\,
            in1 => \N__20797\,
            in2 => \N__18851\,
            in3 => \N__21619\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_1\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_RNO_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__20798\,
            in1 => \N__21793\,
            in2 => \N__18848\,
            in3 => \N__18876\,
            lcout => \Lab_UT.dictrl.state_ret_5_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100110000"
        )
    port map (
            in0 => \N__18845\,
            in1 => \N__20800\,
            in2 => \N__21466\,
            in3 => \N__21620\,
            lcout => \Lab_UT.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22311\,
            ce => 'H',
            sr => \N__21987\
        );

    \Lab_UT.dictrl.state_ret_5_RNO_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__20799\,
            in1 => \N__18877\,
            in2 => \N__21792\,
            in3 => \N__19005\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_ret_5_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18839\,
            in2 => \N__18815\,
            in3 => \N__18812\,
            lcout => \Lab_UT.dicRun_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22311\,
            ce => 'H',
            sr => \N__21987\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_4_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__21777\,
            in1 => \N__21364\,
            in2 => \_gnd_net_\,
            in3 => \N__23195\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_0_a3_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011001000"
        )
    port map (
            in0 => \N__18791\,
            in1 => \N__18782\,
            in2 => \N__18776\,
            in3 => \N__18771\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_2_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011000100"
        )
    port map (
            in0 => \N__21377\,
            in1 => \N__19036\,
            in2 => \N__18977\,
            in3 => \N__20943\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_15_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__19892\,
            in1 => \N__18896\,
            in2 => \N__19025\,
            in3 => \N__19011\,
            lcout => \Lab_UT.dictrl.un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22303\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_RNITITL_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__21363\,
            in2 => \N__18976\,
            in3 => \N__23194\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_4_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__19142\,
            in1 => \N__20491\,
            in2 => \N__19413\,
            in3 => \N__21564\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_6_o3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_3_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100010"
        )
    port map (
            in0 => \N__21071\,
            in1 => \N__23196\,
            in2 => \N__18902\,
            in3 => \N__20410\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_1_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__21365\,
            in1 => \_gnd_net_\,
            in2 => \N__18899\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.g1_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g2_2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__23077\,
            in1 => \N__22862\,
            in2 => \_gnd_net_\,
            in3 => \N__22449\,
            lcout => \Lab_UT.dictrl.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_17_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__20650\,
            in1 => \N__19064\,
            in2 => \N__21433\,
            in3 => \N__19049\,
            lcout => \Lab_UT.dictrl.N_16_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_5_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__22556\,
            in1 => \N__22863\,
            in2 => \N__21571\,
            in3 => \N__22451\,
            lcout => \Lab_UT.dictrl.g0_i_a3_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_0_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21208\,
            in2 => \_gnd_net_\,
            in3 => \N__22610\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_0_6_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__20482\,
            in1 => \N__19365\,
            in2 => \N__19220\,
            in3 => \N__23078\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_a3_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_14_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__19607\,
            in1 => \N__23096\,
            in2 => \N__19217\,
            in3 => \N__19214\,
            lcout => \Lab_UT.dictrl.N_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state32_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22973\,
            in1 => \N__19093\,
            in2 => \N__22615\,
            in3 => \N__21247\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_4_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__22450\,
            in1 => \N__20481\,
            in2 => \N__22557\,
            in3 => \N__22609\,
            lcout => \Lab_UT.dictrl.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__21210\,
            in1 => \N__19160\,
            in2 => \_gnd_net_\,
            in3 => \N__19141\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_23_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010011111100"
        )
    port map (
            in0 => \N__19094\,
            in1 => \N__21133\,
            in2 => \N__19067\,
            in3 => \N__19613\,
            lcout => \Lab_UT.dictrl.N_13_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_2_2_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__22864\,
            in1 => \N__23073\,
            in2 => \_gnd_net_\,
            in3 => \N__22459\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_20_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__19619\,
            in1 => \N__21134\,
            in2 => \N__19058\,
            in3 => \N__19055\,
            lcout => \Lab_UT.dictrl.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state32_1_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19449\,
            in2 => \_gnd_net_\,
            in3 => \N__19245\,
            lcout => \Lab_UT.dictrl.next_state32Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_2_3_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__20462\,
            in1 => \N__21534\,
            in2 => \N__22972\,
            in3 => \N__22527\,
            lcout => \Lab_UT.dictrl.g1_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_1_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22976\,
            in1 => \N__19450\,
            in2 => \N__22616\,
            in3 => \N__19246\,
            lcout => \Lab_UT.dictrl.g0_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_4_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__20463\,
            in1 => \N__19326\,
            in2 => \N__23086\,
            in3 => \N__21535\,
            lcout => \Lab_UT.dictrl.g0_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_2_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__19486\,
            in1 => \N__19601\,
            in2 => \N__22611\,
            in3 => \N__19552\,
            lcout => \Lab_UT.dictrl.g1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_rep1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19324\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_fast_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_2_rep2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19325\,
            lcout => bu_rx_data_2_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_2_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19322\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_fast_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19778\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_1_rep2_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19779\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22284\,
            ce => \N__22074\,
            sr => \N__22010\
        );

    \buart.Z_rx.shifter_3_rep1_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22456\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22279\,
            ce => \N__22072\,
            sr => \N__22012\
        );

    \buart.Z_rx.shifter_fast_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22748\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22279\,
            ce => \N__22072\,
            sr => \N__22012\
        );

    \uu2.bitmap_34_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20363\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__21953\
        );

    \uu2.bitmap_162_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19628\,
            in2 => \_gnd_net_\,
            in3 => \N__20065\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__21953\
        );

    \Lab_UT.bcd2segment4.segment_0_2_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101100111"
        )
    port map (
            in0 => \N__20338\,
            in1 => \N__20272\,
            in2 => \N__20216\,
            in3 => \N__20144\,
            lcout => \Lab_UT.bcd2segment4.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_4_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111101100"
        )
    port map (
            in0 => \N__20213\,
            in1 => \N__20141\,
            in2 => \N__20274\,
            in3 => \N__20341\,
            lcout => \Lab_UT.bcd2segment4.segmentUQ_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_5_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111011000"
        )
    port map (
            in0 => \N__20339\,
            in1 => \N__20264\,
            in2 => \N__20217\,
            in3 => \N__20145\,
            lcout => \Lab_UT.bcd2segment4.segmentUQ_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_6_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010100101"
        )
    port map (
            in0 => \N__20214\,
            in1 => \N__20142\,
            in2 => \N__20275\,
            in3 => \N__20342\,
            lcout => \Lab_UT.bcd2segment4.segmentUQ_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_0_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011011011111101"
        )
    port map (
            in0 => \N__20340\,
            in1 => \N__20268\,
            in2 => \N__20218\,
            in3 => \N__20146\,
            lcout => \Lab_UT.bcd2segment4.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_0_1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100101111111"
        )
    port map (
            in0 => \N__20215\,
            in1 => \N__20143\,
            in2 => \N__20276\,
            in3 => \N__20343\,
            lcout => \Lab_UT.bcd2segment4.segment_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segmentUQ_3_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111001010"
        )
    port map (
            in0 => \N__20344\,
            in1 => \N__20273\,
            in2 => \N__20219\,
            in3 => \N__20147\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment4.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_290_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20069\,
            in3 => \N__20059\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__21951\
        );

    \Lab_UT.dictrl.state_0_3_rep1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19908\,
            in1 => \N__20681\,
            in2 => \N__20866\,
            in3 => \N__21774\,
            lcout => \Lab_UT.dictrl.state_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__21988\
        );

    \Lab_UT.dictrl.state_0_fast_3_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__21773\,
            in1 => \N__20865\,
            in2 => \N__20690\,
            in3 => \N__19910\,
            lcout => \Lab_UT.dictrl.state_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__21988\
        );

    \Lab_UT.dictrl.state_0_3_rep2_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__19909\,
            in1 => \N__20682\,
            in2 => \N__20867\,
            in3 => \N__21775\,
            lcout => \Lab_UT.dictrl.state_3_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__21988\
        );

    \Lab_UT.dictrl.state_0_3_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__21772\,
            in1 => \N__20858\,
            in2 => \N__20689\,
            in3 => \N__19907\,
            lcout => \Lab_UT.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22329\,
            ce => 'H',
            sr => \N__21988\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20855\,
            in1 => \N__20601\,
            in2 => \N__21790\,
            in3 => \N__22036\,
            lcout => \Lab_UT.dictrl.g0_0_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_RNO_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__20856\,
            in1 => \_gnd_net_\,
            in2 => \N__21791\,
            in3 => \N__20603\,
            lcout => \Lab_UT.dictrl.g0_0_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_RNO_1_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__20602\,
            in1 => \N__20857\,
            in2 => \_gnd_net_\,
            in3 => \N__21768\,
            lcout => \Lab_UT.dictrl.g0_0_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m35_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__20732\,
            in1 => \N__20604\,
            in2 => \_gnd_net_\,
            in3 => \N__21605\,
            lcout => \Lab_UT.dictrl.N_40_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m12_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100100010"
        )
    port map (
            in0 => \N__21130\,
            in1 => \N__20954\,
            in2 => \N__20662\,
            in3 => \N__21603\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m15_ns_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21455\,
            in1 => \_gnd_net_\,
            in2 => \N__20537\,
            in3 => \N__20420\,
            lcout => \Lab_UT.dictrl.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_6_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__20512\,
            in1 => \N__20492\,
            in2 => \N__23087\,
            in3 => \N__21113\,
            lcout => \Lab_UT.dictrl.g1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__21604\,
            in1 => \N__23170\,
            in2 => \N__21132\,
            in3 => \N__20409\,
            lcout => \Lab_UT.dictrl.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m20_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101010111"
        )
    port map (
            in0 => \N__21129\,
            in1 => \N__20408\,
            in2 => \N__23197\,
            in3 => \N__20953\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIFHHU6_2_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001110011011"
        )
    port map (
            in0 => \N__21454\,
            in1 => \N__21764\,
            in2 => \N__21623\,
            in3 => \N__21280\,
            lcout => \Lab_UT.dictrl.next_state_latmux_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__21182\,
            in1 => \N__21114\,
            in2 => \_gnd_net_\,
            in3 => \N__21602\,
            lcout => \Lab_UT.dictrl.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__22961\,
            in1 => \N__21568\,
            in2 => \N__22871\,
            in3 => \N__23083\,
            lcout => \Lab_UT.dictrl.g1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20909\,
            in1 => \N__21434\,
            in2 => \_gnd_net_\,
            in3 => \N__21281\,
            lcout => \Lab_UT.dictrl.N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_1_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23084\,
            in2 => \_gnd_net_\,
            in3 => \N__22434\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m17_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22825\,
            in1 => \N__21140\,
            in2 => \N__21257\,
            in3 => \N__21254\,
            lcout => \Lab_UT.dictrl.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__m17_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__22959\,
            in1 => \N__22599\,
            in2 => \N__21198\,
            in3 => \N__22502\,
            lcout => \Lab_UT.dictrl.m17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_5_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__23174\,
            in1 => \N__21131\,
            in2 => \_gnd_net_\,
            in3 => \N__20949\,
            lcout => \Lab_UT.dictrl.N_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22960\,
            in1 => \N__22824\,
            in2 => \N__20899\,
            in3 => \N__22503\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g1_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__22435\,
            in1 => \N__22764\,
            in2 => \N__23231\,
            in3 => \N__23228\,
            lcout => \Lab_UT.dictrl.g1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_3_0__g0_i_a3_3_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22826\,
            in1 => \N__22436\,
            in2 => \N__23198\,
            in3 => \N__22504\,
            lcout => \Lab_UT.dictrl.g0_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23085\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__22076\,
            sr => \N__22011\
        );

    \buart.Z_rx.shifter_3_rep2_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22419\,
            lcout => bu_rx_data_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__22076\,
            sr => \N__22011\
        );

    \buart.Z_rx.shifter_5_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22827\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22296\,
            ce => \N__22076\,
            sr => \N__22011\
        );

    \buart.Z_rx.shifter_0_rep1_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22769\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22290\,
            ce => \N__22075\,
            sr => \N__22013\
        );

    \buart.Z_rx.shifter_4_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22520\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22290\,
            ce => \N__22075\,
            sr => \N__22013\
        );
end \INTERFACE\;
