// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 20 2019 23:10:53

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26833;
    wire N__26832;
    wire N__26831;
    wire N__26824;
    wire N__26823;
    wire N__26822;
    wire N__26815;
    wire N__26814;
    wire N__26813;
    wire N__26806;
    wire N__26805;
    wire N__26804;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26788;
    wire N__26787;
    wire N__26786;
    wire N__26779;
    wire N__26778;
    wire N__26777;
    wire N__26770;
    wire N__26769;
    wire N__26768;
    wire N__26761;
    wire N__26760;
    wire N__26759;
    wire N__26742;
    wire N__26739;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26731;
    wire N__26730;
    wire N__26725;
    wire N__26724;
    wire N__26723;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26693;
    wire N__26690;
    wire N__26689;
    wire N__26688;
    wire N__26687;
    wire N__26686;
    wire N__26681;
    wire N__26672;
    wire N__26669;
    wire N__26668;
    wire N__26667;
    wire N__26664;
    wire N__26655;
    wire N__26652;
    wire N__26651;
    wire N__26650;
    wire N__26649;
    wire N__26644;
    wire N__26639;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26623;
    wire N__26618;
    wire N__26617;
    wire N__26616;
    wire N__26615;
    wire N__26612;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26594;
    wire N__26591;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26571;
    wire N__26570;
    wire N__26567;
    wire N__26566;
    wire N__26563;
    wire N__26562;
    wire N__26555;
    wire N__26552;
    wire N__26545;
    wire N__26538;
    wire N__26537;
    wire N__26532;
    wire N__26531;
    wire N__26530;
    wire N__26529;
    wire N__26528;
    wire N__26527;
    wire N__26524;
    wire N__26521;
    wire N__26518;
    wire N__26511;
    wire N__26508;
    wire N__26499;
    wire N__26498;
    wire N__26497;
    wire N__26494;
    wire N__26493;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26482;
    wire N__26473;
    wire N__26470;
    wire N__26467;
    wire N__26460;
    wire N__26459;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26455;
    wire N__26452;
    wire N__26449;
    wire N__26440;
    wire N__26435;
    wire N__26432;
    wire N__26427;
    wire N__26424;
    wire N__26423;
    wire N__26422;
    wire N__26421;
    wire N__26420;
    wire N__26417;
    wire N__26414;
    wire N__26413;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26391;
    wire N__26390;
    wire N__26389;
    wire N__26388;
    wire N__26381;
    wire N__26378;
    wire N__26373;
    wire N__26372;
    wire N__26371;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26360;
    wire N__26359;
    wire N__26358;
    wire N__26355;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26339;
    wire N__26332;
    wire N__26331;
    wire N__26330;
    wire N__26327;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26309;
    wire N__26302;
    wire N__26299;
    wire N__26294;
    wire N__26289;
    wire N__26282;
    wire N__26277;
    wire N__26268;
    wire N__26267;
    wire N__26262;
    wire N__26259;
    wire N__26258;
    wire N__26257;
    wire N__26256;
    wire N__26253;
    wire N__26248;
    wire N__26243;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26231;
    wire N__26230;
    wire N__26229;
    wire N__26228;
    wire N__26223;
    wire N__26216;
    wire N__26213;
    wire N__26208;
    wire N__26205;
    wire N__26204;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26200;
    wire N__26199;
    wire N__26198;
    wire N__26197;
    wire N__26196;
    wire N__26195;
    wire N__26194;
    wire N__26193;
    wire N__26192;
    wire N__26191;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26186;
    wire N__26185;
    wire N__26184;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26176;
    wire N__26175;
    wire N__26174;
    wire N__26173;
    wire N__26172;
    wire N__26171;
    wire N__26170;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26166;
    wire N__26165;
    wire N__26164;
    wire N__26163;
    wire N__26162;
    wire N__26161;
    wire N__26160;
    wire N__26159;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26152;
    wire N__26151;
    wire N__26150;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26145;
    wire N__26144;
    wire N__26143;
    wire N__26142;
    wire N__26141;
    wire N__26140;
    wire N__26139;
    wire N__26138;
    wire N__26137;
    wire N__26136;
    wire N__26135;
    wire N__26134;
    wire N__26133;
    wire N__26132;
    wire N__26131;
    wire N__26130;
    wire N__26129;
    wire N__26128;
    wire N__26127;
    wire N__26126;
    wire N__26125;
    wire N__26124;
    wire N__26123;
    wire N__26122;
    wire N__26121;
    wire N__26120;
    wire N__26119;
    wire N__26118;
    wire N__26117;
    wire N__26116;
    wire N__26115;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25925;
    wire N__25924;
    wire N__25919;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25899;
    wire N__25896;
    wire N__25891;
    wire N__25888;
    wire N__25881;
    wire N__25880;
    wire N__25879;
    wire N__25878;
    wire N__25877;
    wire N__25876;
    wire N__25875;
    wire N__25874;
    wire N__25873;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25842;
    wire N__25841;
    wire N__25840;
    wire N__25839;
    wire N__25838;
    wire N__25837;
    wire N__25836;
    wire N__25835;
    wire N__25834;
    wire N__25833;
    wire N__25832;
    wire N__25831;
    wire N__25830;
    wire N__25829;
    wire N__25828;
    wire N__25827;
    wire N__25826;
    wire N__25825;
    wire N__25824;
    wire N__25823;
    wire N__25822;
    wire N__25821;
    wire N__25820;
    wire N__25819;
    wire N__25818;
    wire N__25817;
    wire N__25816;
    wire N__25815;
    wire N__25814;
    wire N__25813;
    wire N__25812;
    wire N__25811;
    wire N__25810;
    wire N__25809;
    wire N__25808;
    wire N__25807;
    wire N__25806;
    wire N__25805;
    wire N__25804;
    wire N__25803;
    wire N__25802;
    wire N__25801;
    wire N__25800;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25784;
    wire N__25781;
    wire N__25780;
    wire N__25779;
    wire N__25778;
    wire N__25777;
    wire N__25776;
    wire N__25775;
    wire N__25774;
    wire N__25773;
    wire N__25772;
    wire N__25771;
    wire N__25770;
    wire N__25769;
    wire N__25768;
    wire N__25767;
    wire N__25766;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25598;
    wire N__25595;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25587;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25577;
    wire N__25572;
    wire N__25569;
    wire N__25560;
    wire N__25559;
    wire N__25558;
    wire N__25557;
    wire N__25556;
    wire N__25555;
    wire N__25554;
    wire N__25553;
    wire N__25550;
    wire N__25543;
    wire N__25534;
    wire N__25531;
    wire N__25524;
    wire N__25523;
    wire N__25522;
    wire N__25521;
    wire N__25520;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25504;
    wire N__25503;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25497;
    wire N__25496;
    wire N__25495;
    wire N__25494;
    wire N__25493;
    wire N__25490;
    wire N__25485;
    wire N__25482;
    wire N__25481;
    wire N__25478;
    wire N__25475;
    wire N__25470;
    wire N__25467;
    wire N__25458;
    wire N__25457;
    wire N__25456;
    wire N__25453;
    wire N__25450;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25440;
    wire N__25439;
    wire N__25434;
    wire N__25431;
    wire N__25426;
    wire N__25421;
    wire N__25418;
    wire N__25409;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25394;
    wire N__25389;
    wire N__25386;
    wire N__25379;
    wire N__25374;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25362;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25331;
    wire N__25330;
    wire N__25329;
    wire N__25324;
    wire N__25321;
    wire N__25318;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25299;
    wire N__25298;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25284;
    wire N__25277;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25265;
    wire N__25264;
    wire N__25261;
    wire N__25260;
    wire N__25257;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25227;
    wire N__25226;
    wire N__25223;
    wire N__25222;
    wire N__25221;
    wire N__25220;
    wire N__25217;
    wire N__25212;
    wire N__25209;
    wire N__25206;
    wire N__25203;
    wire N__25200;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25184;
    wire N__25183;
    wire N__25176;
    wire N__25173;
    wire N__25172;
    wire N__25171;
    wire N__25170;
    wire N__25169;
    wire N__25168;
    wire N__25167;
    wire N__25164;
    wire N__25163;
    wire N__25162;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25136;
    wire N__25131;
    wire N__25126;
    wire N__25123;
    wire N__25116;
    wire N__25113;
    wire N__25104;
    wire N__25103;
    wire N__25102;
    wire N__25101;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25090;
    wire N__25089;
    wire N__25088;
    wire N__25087;
    wire N__25080;
    wire N__25079;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25071;
    wire N__25068;
    wire N__25061;
    wire N__25058;
    wire N__25053;
    wire N__25048;
    wire N__25043;
    wire N__25032;
    wire N__25031;
    wire N__25030;
    wire N__25029;
    wire N__25028;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24977;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24954;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24937;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24909;
    wire N__24906;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24893;
    wire N__24892;
    wire N__24891;
    wire N__24890;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24878;
    wire N__24875;
    wire N__24872;
    wire N__24869;
    wire N__24864;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24824;
    wire N__24821;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24795;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24779;
    wire N__24776;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24760;
    wire N__24757;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24741;
    wire N__24740;
    wire N__24739;
    wire N__24736;
    wire N__24731;
    wire N__24730;
    wire N__24727;
    wire N__24724;
    wire N__24723;
    wire N__24720;
    wire N__24719;
    wire N__24718;
    wire N__24713;
    wire N__24710;
    wire N__24703;
    wire N__24696;
    wire N__24695;
    wire N__24694;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24688;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24673;
    wire N__24670;
    wire N__24663;
    wire N__24660;
    wire N__24657;
    wire N__24652;
    wire N__24649;
    wire N__24646;
    wire N__24641;
    wire N__24636;
    wire N__24633;
    wire N__24632;
    wire N__24631;
    wire N__24628;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24603;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24579;
    wire N__24578;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24562;
    wire N__24555;
    wire N__24554;
    wire N__24553;
    wire N__24552;
    wire N__24551;
    wire N__24548;
    wire N__24547;
    wire N__24546;
    wire N__24545;
    wire N__24544;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24536;
    wire N__24535;
    wire N__24534;
    wire N__24533;
    wire N__24528;
    wire N__24525;
    wire N__24524;
    wire N__24523;
    wire N__24522;
    wire N__24521;
    wire N__24518;
    wire N__24515;
    wire N__24512;
    wire N__24509;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24491;
    wire N__24490;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24484;
    wire N__24481;
    wire N__24478;
    wire N__24469;
    wire N__24466;
    wire N__24463;
    wire N__24460;
    wire N__24459;
    wire N__24458;
    wire N__24451;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24406;
    wire N__24401;
    wire N__24394;
    wire N__24383;
    wire N__24372;
    wire N__24369;
    wire N__24368;
    wire N__24365;
    wire N__24362;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24342;
    wire N__24341;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24324;
    wire N__24323;
    wire N__24322;
    wire N__24321;
    wire N__24320;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24313;
    wire N__24310;
    wire N__24309;
    wire N__24308;
    wire N__24307;
    wire N__24306;
    wire N__24305;
    wire N__24304;
    wire N__24303;
    wire N__24300;
    wire N__24295;
    wire N__24294;
    wire N__24293;
    wire N__24292;
    wire N__24283;
    wire N__24280;
    wire N__24279;
    wire N__24278;
    wire N__24277;
    wire N__24272;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24254;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24240;
    wire N__24237;
    wire N__24234;
    wire N__24229;
    wire N__24226;
    wire N__24223;
    wire N__24220;
    wire N__24217;
    wire N__24210;
    wire N__24201;
    wire N__24196;
    wire N__24191;
    wire N__24186;
    wire N__24183;
    wire N__24178;
    wire N__24173;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24145;
    wire N__24144;
    wire N__24141;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24113;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24062;
    wire N__24059;
    wire N__24058;
    wire N__24057;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24053;
    wire N__24052;
    wire N__24051;
    wire N__24050;
    wire N__24049;
    wire N__24048;
    wire N__24045;
    wire N__24042;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24038;
    wire N__24037;
    wire N__24036;
    wire N__24035;
    wire N__24034;
    wire N__24033;
    wire N__24032;
    wire N__24031;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24017;
    wire N__24016;
    wire N__24015;
    wire N__24014;
    wire N__24013;
    wire N__24012;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__24002;
    wire N__24001;
    wire N__24000;
    wire N__23999;
    wire N__23998;
    wire N__23997;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23984;
    wire N__23983;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23966;
    wire N__23965;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23959;
    wire N__23958;
    wire N__23955;
    wire N__23940;
    wire N__23935;
    wire N__23930;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23912;
    wire N__23911;
    wire N__23910;
    wire N__23909;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23893;
    wire N__23890;
    wire N__23883;
    wire N__23876;
    wire N__23869;
    wire N__23866;
    wire N__23859;
    wire N__23854;
    wire N__23849;
    wire N__23840;
    wire N__23833;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23827;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23805;
    wire N__23802;
    wire N__23793;
    wire N__23790;
    wire N__23783;
    wire N__23776;
    wire N__23769;
    wire N__23762;
    wire N__23759;
    wire N__23754;
    wire N__23749;
    wire N__23744;
    wire N__23735;
    wire N__23728;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23694;
    wire N__23693;
    wire N__23692;
    wire N__23691;
    wire N__23684;
    wire N__23681;
    wire N__23680;
    wire N__23677;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23663;
    wire N__23662;
    wire N__23655;
    wire N__23646;
    wire N__23643;
    wire N__23642;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23630;
    wire N__23625;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23609;
    wire N__23608;
    wire N__23607;
    wire N__23606;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23600;
    wire N__23593;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23581;
    wire N__23580;
    wire N__23579;
    wire N__23578;
    wire N__23575;
    wire N__23572;
    wire N__23565;
    wire N__23562;
    wire N__23555;
    wire N__23544;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23489;
    wire N__23488;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23482;
    wire N__23475;
    wire N__23474;
    wire N__23473;
    wire N__23472;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23462;
    wire N__23457;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23418;
    wire N__23417;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23404;
    wire N__23403;
    wire N__23402;
    wire N__23397;
    wire N__23390;
    wire N__23385;
    wire N__23382;
    wire N__23381;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23369;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23354;
    wire N__23349;
    wire N__23344;
    wire N__23343;
    wire N__23342;
    wire N__23335;
    wire N__23334;
    wire N__23331;
    wire N__23330;
    wire N__23329;
    wire N__23328;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23310;
    wire N__23305;
    wire N__23300;
    wire N__23295;
    wire N__23292;
    wire N__23291;
    wire N__23290;
    wire N__23289;
    wire N__23286;
    wire N__23279;
    wire N__23278;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23266;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23252;
    wire N__23251;
    wire N__23250;
    wire N__23249;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23199;
    wire N__23192;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23165;
    wire N__23164;
    wire N__23163;
    wire N__23162;
    wire N__23161;
    wire N__23160;
    wire N__23159;
    wire N__23156;
    wire N__23155;
    wire N__23154;
    wire N__23153;
    wire N__23152;
    wire N__23149;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23133;
    wire N__23132;
    wire N__23129;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23119;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23090;
    wire N__23085;
    wire N__23084;
    wire N__23083;
    wire N__23082;
    wire N__23079;
    wire N__23074;
    wire N__23071;
    wire N__23066;
    wire N__23063;
    wire N__23060;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23041;
    wire N__23036;
    wire N__23029;
    wire N__23026;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22977;
    wire N__22974;
    wire N__22973;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22967;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22952;
    wire N__22949;
    wire N__22948;
    wire N__22947;
    wire N__22946;
    wire N__22945;
    wire N__22944;
    wire N__22943;
    wire N__22940;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22921;
    wire N__22914;
    wire N__22907;
    wire N__22904;
    wire N__22899;
    wire N__22894;
    wire N__22889;
    wire N__22878;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22819;
    wire N__22818;
    wire N__22817;
    wire N__22816;
    wire N__22815;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22809;
    wire N__22802;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22781;
    wire N__22778;
    wire N__22777;
    wire N__22776;
    wire N__22775;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22751;
    wire N__22750;
    wire N__22745;
    wire N__22742;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22721;
    wire N__22718;
    wire N__22713;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22643;
    wire N__22642;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22605;
    wire N__22604;
    wire N__22603;
    wire N__22600;
    wire N__22595;
    wire N__22590;
    wire N__22589;
    wire N__22588;
    wire N__22587;
    wire N__22584;
    wire N__22579;
    wire N__22576;
    wire N__22569;
    wire N__22568;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22560;
    wire N__22553;
    wire N__22552;
    wire N__22551;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22533;
    wire N__22524;
    wire N__22523;
    wire N__22522;
    wire N__22521;
    wire N__22518;
    wire N__22513;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22491;
    wire N__22490;
    wire N__22489;
    wire N__22488;
    wire N__22487;
    wire N__22486;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22463;
    wire N__22462;
    wire N__22459;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22425;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22419;
    wire N__22418;
    wire N__22415;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22388;
    wire N__22383;
    wire N__22380;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22372;
    wire N__22371;
    wire N__22370;
    wire N__22367;
    wire N__22360;
    wire N__22357;
    wire N__22354;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22340;
    wire N__22335;
    wire N__22334;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22308;
    wire N__22305;
    wire N__22304;
    wire N__22303;
    wire N__22302;
    wire N__22299;
    wire N__22298;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22280;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22260;
    wire N__22257;
    wire N__22254;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22237;
    wire N__22234;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22214;
    wire N__22213;
    wire N__22210;
    wire N__22209;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22192;
    wire N__22185;
    wire N__22184;
    wire N__22179;
    wire N__22178;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22149;
    wire N__22148;
    wire N__22147;
    wire N__22146;
    wire N__22145;
    wire N__22144;
    wire N__22143;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22118;
    wire N__22113;
    wire N__22112;
    wire N__22111;
    wire N__22110;
    wire N__22109;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22084;
    wire N__22071;
    wire N__22070;
    wire N__22069;
    wire N__22066;
    wire N__22065;
    wire N__22062;
    wire N__22059;
    wire N__22056;
    wire N__22053;
    wire N__22052;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22017;
    wire N__22012;
    wire N__21999;
    wire N__21998;
    wire N__21997;
    wire N__21994;
    wire N__21987;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21975;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21960;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21952;
    wire N__21949;
    wire N__21948;
    wire N__21943;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21918;
    wire N__21915;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21907;
    wire N__21906;
    wire N__21905;
    wire N__21904;
    wire N__21899;
    wire N__21896;
    wire N__21889;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21848;
    wire N__21847;
    wire N__21844;
    wire N__21839;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21815;
    wire N__21810;
    wire N__21807;
    wire N__21806;
    wire N__21805;
    wire N__21804;
    wire N__21803;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21779;
    wire N__21776;
    wire N__21775;
    wire N__21774;
    wire N__21771;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21730;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21709;
    wire N__21704;
    wire N__21701;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21685;
    wire N__21680;
    wire N__21677;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21624;
    wire N__21621;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21578;
    wire N__21575;
    wire N__21572;
    wire N__21571;
    wire N__21570;
    wire N__21569;
    wire N__21562;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21550;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21538;
    wire N__21531;
    wire N__21530;
    wire N__21529;
    wire N__21526;
    wire N__21525;
    wire N__21518;
    wire N__21517;
    wire N__21514;
    wire N__21513;
    wire N__21510;
    wire N__21505;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21490;
    wire N__21485;
    wire N__21482;
    wire N__21477;
    wire N__21476;
    wire N__21475;
    wire N__21474;
    wire N__21471;
    wire N__21470;
    wire N__21463;
    wire N__21458;
    wire N__21457;
    wire N__21454;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21436;
    wire N__21429;
    wire N__21428;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21420;
    wire N__21417;
    wire N__21410;
    wire N__21409;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21361;
    wire N__21356;
    wire N__21353;
    wire N__21348;
    wire N__21347;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21333;
    wire N__21328;
    wire N__21327;
    wire N__21326;
    wire N__21321;
    wire N__21318;
    wire N__21309;
    wire N__21304;
    wire N__21303;
    wire N__21302;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21277;
    wire N__21264;
    wire N__21263;
    wire N__21260;
    wire N__21259;
    wire N__21258;
    wire N__21257;
    wire N__21256;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21240;
    wire N__21237;
    wire N__21232;
    wire N__21225;
    wire N__21222;
    wire N__21221;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21195;
    wire N__21194;
    wire N__21191;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21178;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21134;
    wire N__21133;
    wire N__21132;
    wire N__21131;
    wire N__21128;
    wire N__21127;
    wire N__21126;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21112;
    wire N__21109;
    wire N__21106;
    wire N__21103;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21080;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21050;
    wire N__21049;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21037;
    wire N__21034;
    wire N__21031;
    wire N__21028;
    wire N__21025;
    wire N__21022;
    wire N__21015;
    wire N__21014;
    wire N__21013;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20999;
    wire N__20996;
    wire N__20991;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20973;
    wire N__20972;
    wire N__20971;
    wire N__20964;
    wire N__20961;
    wire N__20960;
    wire N__20959;
    wire N__20958;
    wire N__20955;
    wire N__20948;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20938;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20922;
    wire N__20921;
    wire N__20920;
    wire N__20917;
    wire N__20912;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20883;
    wire N__20882;
    wire N__20881;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20854;
    wire N__20851;
    wire N__20844;
    wire N__20843;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20789;
    wire N__20788;
    wire N__20785;
    wire N__20784;
    wire N__20783;
    wire N__20778;
    wire N__20775;
    wire N__20770;
    wire N__20763;
    wire N__20762;
    wire N__20761;
    wire N__20760;
    wire N__20759;
    wire N__20758;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20745;
    wire N__20744;
    wire N__20743;
    wire N__20742;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20706;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20643;
    wire N__20634;
    wire N__20633;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20617;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20593;
    wire N__20592;
    wire N__20591;
    wire N__20586;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20578;
    wire N__20577;
    wire N__20576;
    wire N__20567;
    wire N__20562;
    wire N__20555;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20541;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20504;
    wire N__20503;
    wire N__20502;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20489;
    wire N__20488;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20453;
    wire N__20450;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20423;
    wire N__20418;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20403;
    wire N__20402;
    wire N__20399;
    wire N__20396;
    wire N__20395;
    wire N__20394;
    wire N__20387;
    wire N__20384;
    wire N__20379;
    wire N__20376;
    wire N__20375;
    wire N__20372;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20345;
    wire N__20342;
    wire N__20337;
    wire N__20332;
    wire N__20325;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20321;
    wire N__20320;
    wire N__20319;
    wire N__20318;
    wire N__20311;
    wire N__20310;
    wire N__20301;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20284;
    wire N__20283;
    wire N__20282;
    wire N__20279;
    wire N__20274;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20264;
    wire N__20259;
    wire N__20256;
    wire N__20251;
    wire N__20246;
    wire N__20241;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20222;
    wire N__20221;
    wire N__20220;
    wire N__20219;
    wire N__20218;
    wire N__20217;
    wire N__20216;
    wire N__20215;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20207;
    wire N__20206;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20198;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20191;
    wire N__20186;
    wire N__20183;
    wire N__20178;
    wire N__20169;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20152;
    wire N__20149;
    wire N__20144;
    wire N__20143;
    wire N__20140;
    wire N__20135;
    wire N__20130;
    wire N__20123;
    wire N__20116;
    wire N__20113;
    wire N__20104;
    wire N__20099;
    wire N__20094;
    wire N__20093;
    wire N__20092;
    wire N__20091;
    wire N__20090;
    wire N__20087;
    wire N__20086;
    wire N__20083;
    wire N__20082;
    wire N__20079;
    wire N__20078;
    wire N__20077;
    wire N__20076;
    wire N__20075;
    wire N__20072;
    wire N__20071;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20055;
    wire N__20050;
    wire N__20049;
    wire N__20046;
    wire N__20045;
    wire N__20040;
    wire N__20035;
    wire N__20032;
    wire N__20031;
    wire N__20028;
    wire N__20023;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19987;
    wire N__19982;
    wire N__19979;
    wire N__19974;
    wire N__19971;
    wire N__19962;
    wire N__19961;
    wire N__19960;
    wire N__19959;
    wire N__19958;
    wire N__19957;
    wire N__19956;
    wire N__19955;
    wire N__19954;
    wire N__19953;
    wire N__19952;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19926;
    wire N__19921;
    wire N__19918;
    wire N__19917;
    wire N__19914;
    wire N__19909;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19893;
    wire N__19890;
    wire N__19885;
    wire N__19880;
    wire N__19875;
    wire N__19872;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19850;
    wire N__19845;
    wire N__19844;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19833;
    wire N__19832;
    wire N__19831;
    wire N__19830;
    wire N__19825;
    wire N__19824;
    wire N__19823;
    wire N__19822;
    wire N__19821;
    wire N__19820;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19810;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19788;
    wire N__19783;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19775;
    wire N__19768;
    wire N__19767;
    wire N__19762;
    wire N__19757;
    wire N__19752;
    wire N__19749;
    wire N__19740;
    wire N__19737;
    wire N__19736;
    wire N__19735;
    wire N__19734;
    wire N__19731;
    wire N__19730;
    wire N__19729;
    wire N__19726;
    wire N__19725;
    wire N__19724;
    wire N__19721;
    wire N__19720;
    wire N__19717;
    wire N__19716;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19712;
    wire N__19711;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19685;
    wire N__19682;
    wire N__19679;
    wire N__19672;
    wire N__19667;
    wire N__19666;
    wire N__19665;
    wire N__19662;
    wire N__19655;
    wire N__19652;
    wire N__19645;
    wire N__19642;
    wire N__19639;
    wire N__19632;
    wire N__19629;
    wire N__19624;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19615;
    wire N__19610;
    wire N__19607;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19585;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19538;
    wire N__19535;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19529;
    wire N__19528;
    wire N__19527;
    wire N__19524;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19502;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19478;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19448;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19440;
    wire N__19439;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19424;
    wire N__19423;
    wire N__19422;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19404;
    wire N__19399;
    wire N__19396;
    wire N__19385;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19367;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19357;
    wire N__19352;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19335;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19321;
    wire N__19318;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19314;
    wire N__19313;
    wire N__19312;
    wire N__19311;
    wire N__19310;
    wire N__19307;
    wire N__19306;
    wire N__19305;
    wire N__19298;
    wire N__19295;
    wire N__19290;
    wire N__19285;
    wire N__19280;
    wire N__19275;
    wire N__19272;
    wire N__19271;
    wire N__19264;
    wire N__19261;
    wire N__19256;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19230;
    wire N__19227;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19215;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19197;
    wire N__19194;
    wire N__19193;
    wire N__19192;
    wire N__19191;
    wire N__19190;
    wire N__19185;
    wire N__19182;
    wire N__19177;
    wire N__19172;
    wire N__19165;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19157;
    wire N__19154;
    wire N__19151;
    wire N__19150;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19129;
    wire N__19124;
    wire N__19121;
    wire N__19118;
    wire N__19117;
    wire N__19116;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19101;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19085;
    wire N__19076;
    wire N__19059;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19049;
    wire N__19048;
    wire N__19047;
    wire N__19042;
    wire N__19041;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19023;
    wire N__19020;
    wire N__19019;
    wire N__19018;
    wire N__19017;
    wire N__19014;
    wire N__19009;
    wire N__19006;
    wire N__18999;
    wire N__18998;
    wire N__18997;
    wire N__18996;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18971;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18935;
    wire N__18934;
    wire N__18933;
    wire N__18932;
    wire N__18931;
    wire N__18928;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18920;
    wire N__18919;
    wire N__18914;
    wire N__18911;
    wire N__18910;
    wire N__18909;
    wire N__18906;
    wire N__18901;
    wire N__18898;
    wire N__18893;
    wire N__18892;
    wire N__18891;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18876;
    wire N__18875;
    wire N__18872;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18854;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18839;
    wire N__18834;
    wire N__18831;
    wire N__18822;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18804;
    wire N__18797;
    wire N__18792;
    wire N__18787;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18760;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18740;
    wire N__18737;
    wire N__18734;
    wire N__18731;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18725;
    wire N__18724;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18701;
    wire N__18698;
    wire N__18695;
    wire N__18692;
    wire N__18689;
    wire N__18686;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18665;
    wire N__18662;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18646;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18630;
    wire N__18627;
    wire N__18626;
    wire N__18625;
    wire N__18622;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18606;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18595;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18587;
    wire N__18586;
    wire N__18585;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18570;
    wire N__18569;
    wire N__18566;
    wire N__18563;
    wire N__18560;
    wire N__18559;
    wire N__18556;
    wire N__18553;
    wire N__18548;
    wire N__18545;
    wire N__18542;
    wire N__18537;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18512;
    wire N__18509;
    wire N__18506;
    wire N__18503;
    wire N__18496;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18480;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18399;
    wire N__18396;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18382;
    wire N__18375;
    wire N__18372;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18342;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18337;
    wire N__18328;
    wire N__18325;
    wire N__18324;
    wire N__18323;
    wire N__18322;
    wire N__18321;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18287;
    wire N__18284;
    wire N__18275;
    wire N__18272;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18233;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18203;
    wire N__18200;
    wire N__18199;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18171;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18159;
    wire N__18158;
    wire N__18157;
    wire N__18156;
    wire N__18155;
    wire N__18154;
    wire N__18153;
    wire N__18152;
    wire N__18151;
    wire N__18150;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18138;
    wire N__18137;
    wire N__18130;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18087;
    wire N__18084;
    wire N__18079;
    wire N__18076;
    wire N__18071;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18055;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18003;
    wire N__18000;
    wire N__17999;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17954;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17940;
    wire N__17939;
    wire N__17938;
    wire N__17937;
    wire N__17936;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17920;
    wire N__17913;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17903;
    wire N__17902;
    wire N__17901;
    wire N__17900;
    wire N__17899;
    wire N__17896;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17846;
    wire N__17845;
    wire N__17842;
    wire N__17837;
    wire N__17832;
    wire N__17829;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17805;
    wire N__17802;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17797;
    wire N__17794;
    wire N__17791;
    wire N__17782;
    wire N__17777;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17714;
    wire N__17713;
    wire N__17712;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17700;
    wire N__17695;
    wire N__17688;
    wire N__17687;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17654;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17630;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17558;
    wire N__17557;
    wire N__17556;
    wire N__17555;
    wire N__17552;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17540;
    wire N__17535;
    wire N__17532;
    wire N__17523;
    wire N__17522;
    wire N__17519;
    wire N__17518;
    wire N__17515;
    wire N__17514;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17502;
    wire N__17499;
    wire N__17496;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17457;
    wire N__17454;
    wire N__17451;
    wire N__17448;
    wire N__17445;
    wire N__17442;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17420;
    wire N__17419;
    wire N__17416;
    wire N__17415;
    wire N__17414;
    wire N__17413;
    wire N__17410;
    wire N__17409;
    wire N__17402;
    wire N__17393;
    wire N__17390;
    wire N__17385;
    wire N__17382;
    wire N__17381;
    wire N__17378;
    wire N__17377;
    wire N__17376;
    wire N__17375;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17367;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17353;
    wire N__17350;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17334;
    wire N__17331;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17165;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17145;
    wire N__17144;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17117;
    wire N__17114;
    wire N__17113;
    wire N__17112;
    wire N__17111;
    wire N__17108;
    wire N__17107;
    wire N__17104;
    wire N__17097;
    wire N__17096;
    wire N__17095;
    wire N__17094;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17082;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17061;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17045;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17037;
    wire N__17036;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17015;
    wire N__17014;
    wire N__17013;
    wire N__17012;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16989;
    wire N__16988;
    wire N__16987;
    wire N__16984;
    wire N__16983;
    wire N__16980;
    wire N__16979;
    wire N__16978;
    wire N__16965;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16955;
    wire N__16952;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16944;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16895;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16863;
    wire N__16862;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16856;
    wire N__16853;
    wire N__16850;
    wire N__16839;
    wire N__16836;
    wire N__16835;
    wire N__16834;
    wire N__16833;
    wire N__16832;
    wire N__16831;
    wire N__16830;
    wire N__16829;
    wire N__16822;
    wire N__16819;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16801;
    wire N__16798;
    wire N__16797;
    wire N__16796;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16779;
    wire N__16770;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16726;
    wire N__16721;
    wire N__16720;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16697;
    wire N__16694;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16684;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16644;
    wire N__16643;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16601;
    wire N__16600;
    wire N__16599;
    wire N__16594;
    wire N__16593;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16578;
    wire N__16575;
    wire N__16570;
    wire N__16567;
    wire N__16562;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16535;
    wire N__16534;
    wire N__16533;
    wire N__16532;
    wire N__16531;
    wire N__16530;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16490;
    wire N__16489;
    wire N__16486;
    wire N__16481;
    wire N__16476;
    wire N__16475;
    wire N__16472;
    wire N__16471;
    wire N__16468;
    wire N__16465;
    wire N__16462;
    wire N__16457;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16424;
    wire N__16423;
    wire N__16422;
    wire N__16419;
    wire N__16418;
    wire N__16415;
    wire N__16412;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16391;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16379;
    wire N__16378;
    wire N__16377;
    wire N__16376;
    wire N__16375;
    wire N__16374;
    wire N__16371;
    wire N__16358;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16337;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16307;
    wire N__16304;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16287;
    wire N__16286;
    wire N__16283;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16254;
    wire N__16253;
    wire N__16252;
    wire N__16251;
    wire N__16250;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16242;
    wire N__16241;
    wire N__16240;
    wire N__16239;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16226;
    wire N__16223;
    wire N__16214;
    wire N__16209;
    wire N__16198;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16181;
    wire N__16178;
    wire N__16175;
    wire N__16174;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16130;
    wire N__16129;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16117;
    wire N__16114;
    wire N__16109;
    wire N__16104;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16089;
    wire N__16086;
    wire N__16085;
    wire N__16082;
    wire N__16081;
    wire N__16078;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15985;
    wire N__15980;
    wire N__15975;
    wire N__15972;
    wire N__15971;
    wire N__15968;
    wire N__15965;
    wire N__15964;
    wire N__15963;
    wire N__15962;
    wire N__15961;
    wire N__15960;
    wire N__15957;
    wire N__15950;
    wire N__15943;
    wire N__15940;
    wire N__15935;
    wire N__15930;
    wire N__15929;
    wire N__15926;
    wire N__15925;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15919;
    wire N__15918;
    wire N__15915;
    wire N__15908;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15885;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15878;
    wire N__15875;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15851;
    wire N__15844;
    wire N__15839;
    wire N__15836;
    wire N__15831;
    wire N__15828;
    wire N__15827;
    wire N__15826;
    wire N__15825;
    wire N__15824;
    wire N__15823;
    wire N__15822;
    wire N__15819;
    wire N__15812;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15776;
    wire N__15775;
    wire N__15774;
    wire N__15773;
    wire N__15772;
    wire N__15771;
    wire N__15770;
    wire N__15769;
    wire N__15768;
    wire N__15757;
    wire N__15750;
    wire N__15745;
    wire N__15742;
    wire N__15737;
    wire N__15732;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15720;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15701;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15693;
    wire N__15692;
    wire N__15689;
    wire N__15684;
    wire N__15681;
    wire N__15676;
    wire N__15673;
    wire N__15666;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15630;
    wire N__15629;
    wire N__15628;
    wire N__15627;
    wire N__15626;
    wire N__15625;
    wire N__15624;
    wire N__15623;
    wire N__15620;
    wire N__15615;
    wire N__15608;
    wire N__15607;
    wire N__15606;
    wire N__15603;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15553;
    wire N__15548;
    wire N__15543;
    wire N__15540;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15515;
    wire N__15514;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15506;
    wire N__15505;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15482;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15422;
    wire N__15421;
    wire N__15418;
    wire N__15415;
    wire N__15414;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15410;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15390;
    wire N__15387;
    wire N__15382;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15366;
    wire N__15365;
    wire N__15364;
    wire N__15361;
    wire N__15356;
    wire N__15353;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15341;
    wire N__15340;
    wire N__15337;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15325;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15257;
    wire N__15254;
    wire N__15253;
    wire N__15250;
    wire N__15249;
    wire N__15248;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15182;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15155;
    wire N__15154;
    wire N__15153;
    wire N__15152;
    wire N__15151;
    wire N__15138;
    wire N__15135;
    wire N__15134;
    wire N__15133;
    wire N__15132;
    wire N__15131;
    wire N__15130;
    wire N__15125;
    wire N__15116;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15069;
    wire N__15068;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15047;
    wire N__15046;
    wire N__15045;
    wire N__15044;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14960;
    wire N__14959;
    wire N__14958;
    wire N__14957;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14914;
    wire N__14907;
    wire N__14898;
    wire N__14895;
    wire N__14894;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14883;
    wire N__14882;
    wire N__14879;
    wire N__14874;
    wire N__14869;
    wire N__14866;
    wire N__14863;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14834;
    wire N__14833;
    wire N__14832;
    wire N__14829;
    wire N__14828;
    wire N__14827;
    wire N__14826;
    wire N__14825;
    wire N__14824;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14803;
    wire N__14798;
    wire N__14793;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14756;
    wire N__14755;
    wire N__14752;
    wire N__14747;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14697;
    wire N__14696;
    wire N__14691;
    wire N__14688;
    wire N__14685;
    wire N__14684;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14667;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14567;
    wire N__14564;
    wire N__14563;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14522;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14421;
    wire N__14420;
    wire N__14417;
    wire N__14416;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14402;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14388;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14372;
    wire N__14371;
    wire N__14370;
    wire N__14369;
    wire N__14368;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14352;
    wire N__14351;
    wire N__14350;
    wire N__14347;
    wire N__14342;
    wire N__14339;
    wire N__14334;
    wire N__14333;
    wire N__14332;
    wire N__14331;
    wire N__14330;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14318;
    wire N__14315;
    wire N__14306;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14280;
    wire N__14279;
    wire N__14278;
    wire N__14277;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14244;
    wire N__14243;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14193;
    wire N__14190;
    wire N__14187;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14160;
    wire N__14157;
    wire N__14154;
    wire N__14153;
    wire N__14152;
    wire N__14151;
    wire N__14150;
    wire N__14149;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14129;
    wire N__14124;
    wire N__14123;
    wire N__14122;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14108;
    wire N__14107;
    wire N__14098;
    wire N__14095;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14061;
    wire N__14060;
    wire N__14059;
    wire N__14058;
    wire N__14057;
    wire N__14056;
    wire N__14047;
    wire N__14046;
    wire N__14045;
    wire N__14042;
    wire N__14039;
    wire N__14036;
    wire N__14031;
    wire N__14026;
    wire N__14023;
    wire N__14018;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13995;
    wire N__13992;
    wire N__13991;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13960;
    wire N__13959;
    wire N__13958;
    wire N__13957;
    wire N__13956;
    wire N__13955;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13936;
    wire N__13931;
    wire N__13928;
    wire N__13927;
    wire N__13926;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13886;
    wire N__13885;
    wire N__13884;
    wire N__13883;
    wire N__13882;
    wire N__13881;
    wire N__13878;
    wire N__13877;
    wire N__13876;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13840;
    wire N__13839;
    wire N__13838;
    wire N__13835;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13816;
    wire N__13811;
    wire N__13804;
    wire N__13797;
    wire N__13794;
    wire N__13791;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13778;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13703;
    wire N__13702;
    wire N__13701;
    wire N__13700;
    wire N__13699;
    wire N__13692;
    wire N__13689;
    wire N__13688;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13680;
    wire N__13679;
    wire N__13678;
    wire N__13673;
    wire N__13672;
    wire N__13671;
    wire N__13668;
    wire N__13663;
    wire N__13658;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13642;
    wire N__13639;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13574;
    wire N__13573;
    wire N__13572;
    wire N__13571;
    wire N__13570;
    wire N__13569;
    wire N__13568;
    wire N__13563;
    wire N__13556;
    wire N__13555;
    wire N__13550;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13540;
    wire N__13539;
    wire N__13538;
    wire N__13537;
    wire N__13536;
    wire N__13535;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13477;
    wire N__13474;
    wire N__13455;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13451;
    wire N__13448;
    wire N__13447;
    wire N__13444;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13434;
    wire N__13433;
    wire N__13426;
    wire N__13423;
    wire N__13416;
    wire N__13415;
    wire N__13414;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13409;
    wire N__13408;
    wire N__13405;
    wire N__13404;
    wire N__13403;
    wire N__13400;
    wire N__13395;
    wire N__13390;
    wire N__13387;
    wire N__13382;
    wire N__13375;
    wire N__13370;
    wire N__13367;
    wire N__13360;
    wire N__13357;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13335;
    wire N__13332;
    wire N__13329;
    wire N__13326;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13298;
    wire N__13297;
    wire N__13290;
    wire N__13287;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13276;
    wire N__13271;
    wire N__13266;
    wire N__13265;
    wire N__13262;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13250;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13238;
    wire N__13235;
    wire N__13234;
    wire N__13231;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13193;
    wire N__13192;
    wire N__13189;
    wire N__13184;
    wire N__13179;
    wire N__13176;
    wire N__13175;
    wire N__13174;
    wire N__13171;
    wire N__13166;
    wire N__13161;
    wire N__13158;
    wire N__13157;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13127;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13066;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12997;
    wire N__12996;
    wire N__12995;
    wire N__12994;
    wire N__12989;
    wire N__12986;
    wire N__12979;
    wire N__12976;
    wire N__12969;
    wire N__12968;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12929;
    wire N__12926;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12890;
    wire N__12889;
    wire N__12888;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12833;
    wire N__12830;
    wire N__12829;
    wire N__12828;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12811;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12782;
    wire N__12781;
    wire N__12780;
    wire N__12779;
    wire N__12770;
    wire N__12767;
    wire N__12762;
    wire N__12761;
    wire N__12758;
    wire N__12755;
    wire N__12754;
    wire N__12753;
    wire N__12752;
    wire N__12743;
    wire N__12740;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12725;
    wire N__12722;
    wire N__12721;
    wire N__12718;
    wire N__12713;
    wire N__12712;
    wire N__12711;
    wire N__12710;
    wire N__12709;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12691;
    wire N__12684;
    wire N__12683;
    wire N__12682;
    wire N__12679;
    wire N__12678;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12670;
    wire N__12669;
    wire N__12668;
    wire N__12661;
    wire N__12650;
    wire N__12647;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12614;
    wire N__12613;
    wire N__12612;
    wire N__12611;
    wire N__12610;
    wire N__12609;
    wire N__12608;
    wire N__12599;
    wire N__12590;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12528;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12491;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12473;
    wire N__12470;
    wire N__12469;
    wire N__12468;
    wire N__12467;
    wire N__12464;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12452;
    wire N__12451;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12432;
    wire N__12423;
    wire N__12422;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12406;
    wire N__12403;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12384;
    wire N__12375;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12354;
    wire N__12351;
    wire N__12350;
    wire N__12347;
    wire N__12346;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12334;
    wire N__12331;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12257;
    wire N__12254;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12237;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12214;
    wire N__12207;
    wire N__12206;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12192;
    wire N__12191;
    wire N__12186;
    wire N__12179;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12162;
    wire N__12159;
    wire N__12154;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12126;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12099;
    wire N__12098;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12056;
    wire N__12051;
    wire N__12048;
    wire N__12047;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12041;
    wire N__12040;
    wire N__12039;
    wire N__12028;
    wire N__12023;
    wire N__12018;
    wire N__12015;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12007;
    wire N__12006;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11991;
    wire N__11982;
    wire N__11979;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11965;
    wire N__11958;
    wire N__11957;
    wire N__11956;
    wire N__11955;
    wire N__11954;
    wire N__11951;
    wire N__11942;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11930;
    wire N__11929;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11855;
    wire N__11852;
    wire N__11849;
    wire N__11844;
    wire N__11841;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11737;
    wire N__11736;
    wire N__11735;
    wire N__11730;
    wire N__11727;
    wire N__11722;
    wire N__11719;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11681;
    wire N__11680;
    wire N__11677;
    wire N__11672;
    wire N__11669;
    wire N__11664;
    wire N__11663;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11649;
    wire N__11646;
    wire N__11645;
    wire N__11644;
    wire N__11643;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11629;
    wire N__11626;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11616;
    wire N__11615;
    wire N__11604;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11588;
    wire N__11587;
    wire N__11586;
    wire N__11585;
    wire N__11584;
    wire N__11583;
    wire N__11578;
    wire N__11573;
    wire N__11570;
    wire N__11563;
    wire N__11558;
    wire N__11555;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11528;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11504;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11477;
    wire N__11474;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11459;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11415;
    wire N__11412;
    wire N__11411;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11405;
    wire N__11400;
    wire N__11393;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11383;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11358;
    wire N__11351;
    wire N__11346;
    wire N__11345;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11330;
    wire N__11319;
    wire N__11316;
    wire N__11315;
    wire N__11314;
    wire N__11309;
    wire N__11306;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11294;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11260;
    wire N__11255;
    wire N__11252;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11240;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11216;
    wire N__11215;
    wire N__11214;
    wire N__11211;
    wire N__11204;
    wire N__11199;
    wire N__11198;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11180;
    wire N__11175;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11167;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11155;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11138;
    wire N__11135;
    wire N__11130;
    wire N__11125;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11101;
    wire N__11100;
    wire N__11099;
    wire N__11098;
    wire N__11095;
    wire N__11088;
    wire N__11083;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11025;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11017;
    wire N__11014;
    wire N__11009;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10928;
    wire N__10923;
    wire N__10920;
    wire N__10919;
    wire N__10914;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10906;
    wire N__10905;
    wire N__10904;
    wire N__10903;
    wire N__10898;
    wire N__10891;
    wire N__10888;
    wire N__10881;
    wire N__10880;
    wire N__10879;
    wire N__10876;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10868;
    wire N__10863;
    wire N__10856;
    wire N__10851;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10843;
    wire N__10838;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10785;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10773;
    wire N__10772;
    wire N__10771;
    wire N__10770;
    wire N__10767;
    wire N__10760;
    wire N__10757;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10745;
    wire N__10744;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10723;
    wire N__10716;
    wire N__10715;
    wire N__10714;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10686;
    wire N__10679;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10659;
    wire N__10656;
    wire N__10651;
    wire N__10648;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10636;
    wire N__10631;
    wire N__10626;
    wire N__10625;
    wire N__10624;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10591;
    wire N__10586;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10558;
    wire N__10553;
    wire N__10548;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10495;
    wire N__10494;
    wire N__10489;
    wire N__10488;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10480;
    wire N__10477;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10457;
    wire N__10446;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10391;
    wire N__10388;
    wire N__10383;
    wire N__10382;
    wire N__10381;
    wire N__10378;
    wire N__10377;
    wire N__10370;
    wire N__10367;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10355;
    wire N__10354;
    wire N__10353;
    wire N__10350;
    wire N__10345;
    wire N__10342;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10329;
    wire N__10328;
    wire N__10323;
    wire N__10318;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10296;
    wire N__10295;
    wire N__10294;
    wire N__10293;
    wire N__10292;
    wire N__10287;
    wire N__10280;
    wire N__10275;
    wire N__10274;
    wire N__10273;
    wire N__10270;
    wire N__10263;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10255;
    wire N__10248;
    wire N__10245;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10235;
    wire N__10232;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10109;
    wire N__10108;
    wire N__10105;
    wire N__10100;
    wire N__10095;
    wire N__10092;
    wire N__10091;
    wire N__10090;
    wire N__10089;
    wire N__10086;
    wire N__10079;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10069;
    wire N__10064;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10035;
    wire N__10032;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9990;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9935;
    wire N__9932;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9904;
    wire N__9897;
    wire N__9896;
    wire N__9895;
    wire N__9892;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9849;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9834;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9765;
    wire N__9758;
    wire N__9753;
    wire N__9750;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9744;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9710;
    wire N__9705;
    wire N__9702;
    wire N__9701;
    wire N__9696;
    wire N__9693;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9681;
    wire N__9678;
    wire N__9677;
    wire N__9672;
    wire N__9669;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9644;
    wire N__9643;
    wire N__9640;
    wire N__9635;
    wire N__9630;
    wire N__9627;
    wire N__9626;
    wire N__9625;
    wire N__9624;
    wire N__9623;
    wire N__9622;
    wire N__9615;
    wire N__9610;
    wire N__9607;
    wire N__9602;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9588;
    wire N__9587;
    wire N__9586;
    wire N__9585;
    wire N__9576;
    wire N__9573;
    wire N__9572;
    wire N__9571;
    wire N__9568;
    wire N__9561;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9543;
    wire N__9540;
    wire N__9539;
    wire N__9538;
    wire N__9537;
    wire N__9536;
    wire N__9525;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9516;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_15 ;
    wire bfn_1_5_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire resetGen_reset_count_2_2_cascade_;
    wire resetGen_reset_count_2;
    wire bfn_1_9_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire Lab_UT_dispString_m103_ns_1_cascade_;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire buart__rx_N_27_0_i_cascade_;
    wire N_179;
    wire uart_RXD;
    wire \Lab_UT.dispString.N_115_mux ;
    wire \Lab_UT.dispString.N_115_mux_cascade_ ;
    wire buart__rx_bitcount_1;
    wire buart__rx_bitcount_4;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \Lab_UT.dispString.N_177 ;
    wire buart__rx_ser_clk_cascade_;
    wire buart__rx_bitcount_0;
    wire buart__rx_sample;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_1_13_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire buart__rx_ser_clk;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \uu0.un44_ci_cascade_ ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un44_ci ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un66_ci ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un220_ci ;
    wire \uu0.un143_ci_0 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un4_l_count_11 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un4_l_count_16_cascade_ ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.un110_ci ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.un11_l_count_i_g ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un165_ci_0 ;
    wire resetGen_reset_count_1;
    wire N_107;
    wire m72_cascade_;
    wire N_105;
    wire \resetGen.reset_countZ0Z_3 ;
    wire resetGen_reset_count_4;
    wire resetGen_reset_count_0;
    wire buart__rx_hh_0;
    wire \Lab_UT.dictrl.g0_69_1_cascade_ ;
    wire \Lab_UT.dictrl.g1_0_3_1 ;
    wire \Lab_UT.dictrl.g1_5_1_cascade_ ;
    wire \Lab_UT.dictrl.N_61_1 ;
    wire \Lab_UT.dictrl.g1_7_0 ;
    wire \Lab_UT.dictrl.N_1792_1_cascade_ ;
    wire \Lab_UT.dictrl.N_1451_0 ;
    wire \Lab_UT.dictrl.g0_i_a5_2_4_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_a5_2_5 ;
    wire \Lab_UT.dictrl.g0_5_3 ;
    wire \Lab_UT.dictrl.g0_5_4 ;
    wire \Lab_UT.dictrl.g1_6_0 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.un404_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.trig_rd_is_det_cascade_ ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.un306_ci_cascade_ ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.vbuf_count.un328_ci_3_cascade_ ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.un1_l_count_2_2 ;
    wire \uu2.un306_ci ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.un350_ci ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un11_l_count_i ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \buart.Z_tx.un1_bitcount_c3_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0 ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \Lab_UT.dictrl.g0_12_o6_2_2 ;
    wire \Lab_UT.dictrl.N_13_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_10Z0Z_3 ;
    wire \Lab_UT.dictrl.m34_4Z0Z_2 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_ ;
    wire buart__rx_hh_1;
    wire \Lab_UT.dictrl.m40Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.N_10_3 ;
    wire \Lab_UT.dictrl.N_5_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_9Z0Z_3 ;
    wire \Lab_UT.dictrl.g1_4 ;
    wire \Lab_UT.dictrl.N_97_mux_0_cascade_ ;
    wire \Lab_UT.dictrl.N_2435_0 ;
    wire \Lab_UT.dictrl.g1_5_0 ;
    wire \Lab_UT.dictrl.N_97_mux_0 ;
    wire \Lab_UT.dictrl.g0_16_2_cascade_ ;
    wire \Lab_UT.dictrl.N_2446_1 ;
    wire \uu2.mem0.w_addr_0 ;
    wire clk;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.w_addr_1 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \INVuu2.w_addr_user_1C_net ;
    wire \uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.un426_ci_3_cascade_ ;
    wire \INVuu2.w_addr_user_nesr_8C_net ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu2.un284_ci ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.un1_l_count_1_0 ;
    wire vbuf_tx_data_rdy;
    wire \uu0.un88_ci_3 ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un99_ci_0 ;
    wire \Lab_UT.dispString.dOutP_0_iv_2_tz_1 ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_1_1 ;
    wire \Lab_UT.dispString.m74_ns_1 ;
    wire \Lab_UT.dispString.m77_ns_1 ;
    wire \Lab_UT.dispString.N_30_i ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_1 ;
    wire \uu0.sec_clkDZ0 ;
    wire \Lab_UT.alarmstate_1_0_i_1_cascade_ ;
    wire G_215_cascade_;
    wire G_214;
    wire G_216;
    wire G_214_cascade_;
    wire \Lab_UT.m57 ;
    wire G_213;
    wire G_215;
    wire G_213_cascade_;
    wire \Lab_UT.dictrl.m71Z0Z_0 ;
    wire N_105_mux;
    wire \Lab_UT.dispString.N_186 ;
    wire \Lab_UT.dictrl.g0_12_a6_3Z0Z_7 ;
    wire \Lab_UT.dictrl.g0_12_a6_3_8_cascade_ ;
    wire \Lab_UT.dictrl.N_16 ;
    wire N_10_2;
    wire \Lab_UT.dictrl.N_97_mux_0_0_0 ;
    wire \Lab_UT.dictrl.g0_10_1_cascade_ ;
    wire \Lab_UT.dictrl.m63_d_0_ns_1_1 ;
    wire \Lab_UT.dispString.N_112_mux ;
    wire \Lab_UT.dictrl.m27_d_1 ;
    wire \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_ ;
    wire \Lab_UT.dictrl.G_17_i_a5_0_0 ;
    wire \buart.Z_rx.G_17_i_a5_2_5 ;
    wire \buart.Z_rx.G_17_i_a5_2_4 ;
    wire G_17_i_a5_2_6_cascade_;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_fast_2;
    wire \Lab_UT.dictrl.g2_0_3_0_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_4_0 ;
    wire bu_rx_data_1_rep1;
    wire bu_rx_data_2_rep1;
    wire \Lab_UT.dispString.m107_eZ0Z_3 ;
    wire bu_rx_data_fast_5;
    wire \Lab_UT.dictrl.N_10_1_cascade_ ;
    wire \Lab_UT.dictrl.N_17_0 ;
    wire \Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_ ;
    wire N_22;
    wire \Lab_UT.dictrl.N_1105_0 ;
    wire bu_rx_data_fast_7;
    wire \Lab_UT.dictrl.N_10_1 ;
    wire \Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_m2_1_1 ;
    wire \Lab_UT.dictrl.g0_i_m2_1_a6_3_2 ;
    wire bu_rx_data_fast_3;
    wire \Lab_UT.dictrl.N_7_0 ;
    wire \Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_ ;
    wire \Lab_UT.dictrl.G_17_i_a5_1 ;
    wire \uu2.mem0.N_66_i ;
    wire \uu2.mem0.N_56_i ;
    wire \uu2.N_95_mux ;
    wire \uu2.N_96_mux_cascade_ ;
    wire \uu2.mem0.N_63_i ;
    wire \uu2.mem0.N_69_i ;
    wire \uu2.N_96_mux ;
    wire \uu2.mem0.N_71_i ;
    wire \uu2.mem0.N_91_mux ;
    wire \uu2.mem0.N_50_i ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_ ;
    wire \INVuu2.w_addr_displaying_4C_net ;
    wire \uu2.un1_w_user_lf_0_cascade_ ;
    wire \uu2.un1_w_user_lfZ0Z_4 ;
    wire \uu2.un1_w_user_lf_0 ;
    wire L3_tx_data_5;
    wire L3_tx_data_1;
    wire L3_tx_data_4;
    wire \uu2.m35Z0Z_4_cascade_ ;
    wire \uu2.un1_w_user_cr_0_cascade_ ;
    wire \uu2.mem0.w_data_2 ;
    wire \Lab_UT.dispString.N_145 ;
    wire \Lab_UT.dispString.N_146_cascade_ ;
    wire L3_tx_data_2;
    wire L3_tx_data_0;
    wire L3_tx_data_6;
    wire \Lab_UT.dispString.m82_ns_1_cascade_ ;
    wire \Lab_UT.dispString.N_156_cascade_ ;
    wire L3_tx_data_3;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire \Lab_UT.dispString.b1_m_1 ;
    wire \Lab_UT.dispString.m67_ns_1_cascade_ ;
    wire \Lab_UT.dispString.N_143 ;
    wire \Lab_UT.dispString.N_23_0 ;
    wire \Lab_UT.dispString.N_158 ;
    wire \Lab_UT.dispString.m90_ns_1_cascade_ ;
    wire \Lab_UT.dispString.N_164 ;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.dispString.N_166 ;
    wire \Lab_UT.dispString.N_167 ;
    wire Lab_UT_dictrl_g1_0_3;
    wire \Lab_UT.dictrl.g0_12_a6_3_6 ;
    wire \Lab_UT.dictrl.N_10 ;
    wire \Lab_UT.dictrl.g0_12_1 ;
    wire \Lab_UT.dictrl.m15Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.N_8_0 ;
    wire \Lab_UT.dictrl.N_93_cascade_ ;
    wire \Lab_UT.dictrl.N_10_0 ;
    wire \Lab_UT.dictrl.g0_i_a4_0_1 ;
    wire \Lab_UT.dictrl.g0_i_a4_0_3 ;
    wire \Lab_UT.dictrl.m15Z0Z_1 ;
    wire \Lab_UT.dictrl.N_88_mux ;
    wire \Lab_UT.dictrl.g2_0_4_1_cascade_ ;
    wire \Lab_UT.dictrl.m53_d_1_2_cascade_ ;
    wire \Lab_UT.dictrl.N_45_cascade_ ;
    wire bu_rx_data_1_rep2;
    wire \Lab_UT.dictrl.g2_0_3_1 ;
    wire bu_rx_data_2_rep2;
    wire Lab_UT_dictrl_m59_1;
    wire \Lab_UT.dictrl.m59_3_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_3_4 ;
    wire \Lab_UT.dictrl.g2_0_4_4_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_3_2 ;
    wire \Lab_UT.dictrl.g2_0_4_2_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_3 ;
    wire \Lab_UT.dictrl.g2_0_4_cascade_ ;
    wire bu_rx_data_fast_0;
    wire bu_rx_data_fast_4;
    wire bu_rx_data_3_rep1;
    wire \Lab_UT.dictrl.g2_0_3_3 ;
    wire \Lab_UT.dictrl.g2_0_4_3_cascade_ ;
    wire \Lab_UT.dictrl.m12Z0Z_1 ;
    wire \Lab_UT.dictrl.N_11_1_cascade_ ;
    wire \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0 ;
    wire \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_ ;
    wire bu_rx_data_fast_6;
    wire \buart.Z_rx.sample_g ;
    wire \Lab_UT.dictrl.N_100 ;
    wire \Lab_UT.dictrl.next_state_RNO_8Z0Z_0 ;
    wire \Lab_UT.dictrl.m63_d_0_ns_1 ;
    wire \Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ;
    wire \Lab_UT.dictrl.next_state_RNO_3Z0Z_0 ;
    wire \Lab_UT.dictrl.m67_am_1_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ;
    wire \Lab_UT.dictrl.G_17_i_a5_0 ;
    wire \Lab_UT.dictrl.N_65 ;
    wire \Lab_UT.dictrl.N_65_cascade_ ;
    wire \Lab_UT.dictrl.N_101 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.N_91 ;
    wire \uu2.N_28_cascade_ ;
    wire \uu2.bitmap_pmux_26_i_m2_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.N_55_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i7_mux_0 ;
    wire \uu2.N_406_cascade_ ;
    wire \uu2.bitmap_pmux ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.N_207 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.N_195 ;
    wire \INVuu2.bitmap_296C_net ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \uu2.bitmap_pmux_15_ns_1 ;
    wire \INVuu2.bitmap_66C_net ;
    wire o_One_Sec_Pulse;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \INVuu2.bitmap_111C_net ;
    wire \Lab_UT.didp.regrce4.LdAMtens_0 ;
    wire \Lab_UT.didp.countrce4.q_5_3_cascade_ ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.didp.countrce4.un20_qPone ;
    wire \Lab_UT.dictrl.g0_12_a6_0_1 ;
    wire \Lab_UT.dictrl.state_2_rep1 ;
    wire \Lab_UT.dictrl.N_62_1 ;
    wire \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ;
    wire \Lab_UT.dictrl.N_79 ;
    wire \Lab_UT.dictrl.state_i_4_1 ;
    wire \Lab_UT.dictrl.N_99 ;
    wire buart__rx_bitcount_3;
    wire buart__rx_valid_3;
    wire \Lab_UT.dictrl.g0_0_2_1_cascade_ ;
    wire \Lab_UT.dictrl.g2_1_0 ;
    wire \Lab_UT.dictrl.g0_0_2_cascade_ ;
    wire \Lab_UT.dictrl.m27_1 ;
    wire \Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83 ;
    wire \Lab_UT.dictrl.N_61 ;
    wire \Lab_UT.dictrl.N_62_cascade_ ;
    wire \Lab_UT.dictrl.N_9_0 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1 ;
    wire \Lab_UT.dictrl.state_fast_1 ;
    wire \Lab_UT.dictrl.N_1110_1 ;
    wire \Lab_UT.dictrl.N_1459_1 ;
    wire \Lab_UT.dictrl.N_40_8 ;
    wire \Lab_UT.dictrl.N_40_3_cascade_ ;
    wire \Lab_UT.dictrl.N_1102_2 ;
    wire \Lab_UT.dictrl.g2_1_2 ;
    wire \Lab_UT.dictrl.N_1462_2_cascade_ ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4 ;
    wire \Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3 ;
    wire \Lab_UT.dictrl.N_11_0_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1 ;
    wire \Lab_UT.dictrl.next_state_0_0 ;
    wire \Lab_UT.dictrl.N_8 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_ ;
    wire \Lab_UT.dictrl.N_20_0 ;
    wire \Lab_UT.dictrl.N_18_0_cascade_ ;
    wire \Lab_UT.dictrl.state_fast_3 ;
    wire \Lab_UT.dictrl.state_fast_2 ;
    wire \Lab_UT.dictrl.state_1_rep1 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_3_2 ;
    wire \Lab_UT.dictrl.N_11_1 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_4_6 ;
    wire \Lab_UT.dictrl.N_22_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_4_7 ;
    wire \Lab_UT.dictrl.m53_d_1_3 ;
    wire \Lab_UT.dictrl.N_97_mux_5_cascade_ ;
    wire \Lab_UT.dictrl.N_40 ;
    wire \Lab_UT.dictrl.N_62 ;
    wire \Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNO_1Z0Z_2 ;
    wire \Lab_UT.dictrl.next_state_RNO_0Z0Z_2 ;
    wire \Lab_UT.dictrl.state_3_rep1 ;
    wire \Lab_UT.dictrl.next_state_0_2 ;
    wire \Lab_UT.dictrl.next_state_RNINV3PZ0Z_2 ;
    wire \Lab_UT.min2_3 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \INVuu2.bitmap_203C_net ;
    wire \uu2.bitmap_pmux_sn_N_65 ;
    wire \uu2.N_54 ;
    wire \uu2.N_53 ;
    wire \uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_ ;
    wire \INVuu2.w_addr_displaying_1C_net ;
    wire \Lab_UT.min1_2 ;
    wire \Lab_UT.min1_1 ;
    wire \Lab_UT.min1_3 ;
    wire \Lab_UT.min1_0 ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0 ;
    wire \INVuu2.bitmap_197C_net ;
    wire buart__rx_startbit;
    wire buart__rx_N_27_0_i;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire buart__rx_bitcount_2;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.min2_1 ;
    wire \Lab_UT.min2_2 ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.didp.regrce2.LdAStens_0 ;
    wire \Lab_UT.didp.countrce4.q_5_2_cascade_ ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.dispString.m49Z0Z_0 ;
    wire \Lab_UT.dispString.m49Z0Z_1 ;
    wire \Lab_UT.dispString.m49Z0Z_3_cascade_ ;
    wire \Lab_UT.loadalarm_0_cascade_ ;
    wire \Lab_UT.min2_0 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.dictrl.g0_12_a6_1_3_cascade_ ;
    wire \Lab_UT.dictrl.N_18 ;
    wire \Lab_UT.dictrl.m35_0 ;
    wire \Lab_UT.didp.countrce4.un13_qPone ;
    wire \Lab_UT.LdAMtens ;
    wire \Lab_UT.LdAMones ;
    wire \Lab_UT.LdAStens ;
    wire \Lab_UT.dictrl.N_1460_2 ;
    wire \Lab_UT.dictrl.state_fast_0 ;
    wire \Lab_UT.dictrl.N_23_1 ;
    wire G_17_i_0;
    wire \Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_latmux_2_1 ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.dictrl.next_state_0_3 ;
    wire \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ;
    wire \Lab_UT.dictrl.G_17_i_a5_1_1 ;
    wire \Lab_UT.dictrl.state_1_rep2 ;
    wire \Lab_UT.dictrl.N_15_0 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_1 ;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_m2_0_2 ;
    wire \Lab_UT.dictrl.next_state_0_0_2_cascade_ ;
    wire rst;
    wire \Lab_UT.dictrl.g0_12_a6_2_2 ;
    wire \Lab_UT.dictrl.N_19 ;
    wire \Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_ ;
    wire \Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2 ;
    wire \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.N_1792_0_0_0 ;
    wire \Lab_UT.dictrl.m53_d_1_5 ;
    wire bu_rx_data_4_rep1;
    wire \Lab_UT.dictrl.N_40_0 ;
    wire \Lab_UT.dictrl.N_6 ;
    wire \Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_i_m2_i_1 ;
    wire \Lab_UT.dictrl.N_97_mux_1 ;
    wire \Lab_UT.dictrl.g0_i_a5_0_2 ;
    wire \Lab_UT.dictrl.g2_2 ;
    wire \Lab_UT.dictrl.g2_3_cascade_ ;
    wire \Lab_UT.dictrl.next_state_3_1 ;
    wire \Lab_UT.dictrl.g1_1 ;
    wire \Lab_UT.dictrl.N_5 ;
    wire \Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_ ;
    wire \Lab_UT.dictrl.N_9 ;
    wire \Lab_UT.dictrl.g2_1_3 ;
    wire \Lab_UT.dictrl.N_1462_3_cascade_ ;
    wire \Lab_UT.dictrl.N_1102_3 ;
    wire \Lab_UT.dictrl.N_1460_3 ;
    wire \Lab_UT.dictrl.m53_d_1_1 ;
    wire \Lab_UT.dictrl.N_97_mux_3_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.un3_w_addr_user_4_cascade_ ;
    wire \uu2.un3_w_addr_user_5 ;
    wire \uu2.un3_w_addr_user ;
    wire \INVuu2.w_addr_displaying_nesr_5C_net ;
    wire \uu2.un21_w_addr_displaying_0_0 ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.w_addr_displayingZ1Z_4 ;
    wire \uu2.bitmap_pmux_sn_N_33_cascade_ ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.bitmap_pmux_sn_m15_0_1 ;
    wire \uu2.w_addr_displaying_0_rep1_RNIDASJZ0 ;
    wire \uu2.w_addr_displaying_RNIR2PLZ0Z_8 ;
    wire \uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1 ;
    wire \uu2.bitmap_pmux_29_0 ;
    wire \uu2.N_24_0 ;
    wire \uu2.w_addr_displaying_RNIU1AF7Z0Z_0 ;
    wire \INVuu2.w_addr_displaying_3C_net ;
    wire \Lab_UT.dictrl.m12Z0Z_2 ;
    wire \INVuu2.bitmap_215C_net ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.N_198_cascade_ ;
    wire \uu2.N_199 ;
    wire \uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_ ;
    wire \uu2.N_196 ;
    wire \uu2.bitmap_pmux_27_i_m2_ns_1 ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.N_15 ;
    wire \uu2.N_17 ;
    wire \uu2.bitmap_pmux_25_i_m2_ns_1_cascade_ ;
    wire \uu2.N_49 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.N_13 ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_3_cascade_ ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.didp.countrce1.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_2_cascade_ ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.dispString.m49Z0Z_12 ;
    wire \Lab_UT.dispString.m49Z0Z_4_cascade_ ;
    wire \Lab_UT.dispString.N_128_mux ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.didp.countrce1.q_5_1 ;
    wire \Lab_UT.LdASones ;
    wire \Lab_UT.didp.regrce1.LdASones_0 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.dispString.N_180 ;
    wire \Lab_UT.dispString.m49Z0Z_7 ;
    wire \Lab_UT.dispString.m49Z0Z_11 ;
    wire \Lab_UT.didp.countrce1.q_5_0_cascade_ ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.LdMtens_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_5_0_cascade_ ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdMtens_0 ;
    wire \Lab_UT.dictrl.state_0_rep1 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0 ;
    wire \Lab_UT.state_i_4_0 ;
    wire \Lab_UT.dicRun_2 ;
    wire bu_rx_data_7;
    wire bu_rx_data_6;
    wire \Lab_UT.dictrl.g0_i_a4_1_5 ;
    wire \Lab_UT.dictrl.g0_i_a4_1_4_cascade_ ;
    wire bu_rx_data_5;
    wire \Lab_UT.dictrl.N_12 ;
    wire \Lab_UT.dictrl.N_4 ;
    wire bu_rx_data_4;
    wire \Lab_UT.dictrl.N_7 ;
    wire bu_rx_data_3_rep2;
    wire \Lab_UT.N_115 ;
    wire \Lab_UT.dictrl.N_39 ;
    wire bu_rx_data_6_rep1;
    wire \Lab_UT.dictrl.m53_d_1_0 ;
    wire \Lab_UT.dictrl.N_97_mux_2_cascade_ ;
    wire \Lab_UT.dictrl.g2_1 ;
    wire \Lab_UT.dictrl.N_1462_0 ;
    wire \Lab_UT.dictrl.N_1102_0_cascade_ ;
    wire \Lab_UT.dictrl.N_97_mux_7 ;
    wire \Lab_UT.dictrl.N_1106_1_cascade_ ;
    wire \Lab_UT.dictrl.g1_1_1_0 ;
    wire bu_rx_data_7_rep1;
    wire \Lab_UT.dictrl.N_59 ;
    wire \Lab_UT.dictrl.N_97_mux ;
    wire \Lab_UT.dictrl.N_59_cascade_ ;
    wire \Lab_UT.dictrl.state_0_rep2 ;
    wire \Lab_UT.dictrl.N_40_5_cascade_ ;
    wire \Lab_UT.dictrl.N_40_4 ;
    wire \Lab_UT.dictrl.N_40_2_cascade_ ;
    wire \Lab_UT.dictrl.m23_aZ0Z0 ;
    wire \Lab_UT.dictrl.N_40_7 ;
    wire \Lab_UT.dictrl.N_40_7_cascade_ ;
    wire \Lab_UT.dictrl.g2_1_5 ;
    wire \Lab_UT.dictrl.N_1462_5_cascade_ ;
    wire \Lab_UT.dictrl.N_1102_5 ;
    wire bu_rx_data_0_rep1;
    wire bu_rx_data_5_rep1;
    wire bu_rx_data_4_rep2;
    wire \Lab_UT.dictrl.g0_i_m2_0_a7_4_8 ;
    wire \Lab_UT.dictrl.N_19_0 ;
    wire bu_rx_data_6_rep2;
    wire \Lab_UT.dictrl.m40Z0Z_1 ;
    wire \Lab_UT.dictrl.m53_d_1_4 ;
    wire \Lab_UT.dictrl.state_2_rep2 ;
    wire \Lab_UT.dictrl.N_97_mux_6_cascade_ ;
    wire \Lab_UT.dictrl.state_3_rep2 ;
    wire \Lab_UT.dictrl.g2_1_4 ;
    wire \Lab_UT.dictrl.N_1462_4 ;
    wire \Lab_UT.dictrl.N_1102_4_cascade_ ;
    wire \Lab_UT.dictrl.N_6_0 ;
    wire \Lab_UT.dictrl.next_state_2_1 ;
    wire \Lab_UT.dictrl.g0_i_0 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.un28_w_addr_user_i ;
    wire \uu2.un404_ci ;
    wire \uu2.un426_ci_3 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \INVuu2.w_addr_user_5C_net ;
    wire \uu2.w_addr_user_RNI43E87Z0Z_2 ;
    wire \uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_ ;
    wire \uu2.N_397 ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \uu2.w_addr_displayingZ1Z_3 ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.N_32 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.N_20 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.bitmap_RNIE7RKZ0Z_58_cascade_ ;
    wire \uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.bitmap_RNI020QZ0Z_186 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \Lab_UT.sec2_1 ;
    wire \Lab_UT.sec2_3 ;
    wire \Lab_UT.sec2_2 ;
    wire \Lab_UT.sec2_0 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \INVuu2.bitmap_87C_net ;
    wire \Lab_UT.didp.countrce2.q_5_0_cascade_ ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.loadalarm_0 ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.dispString.m49Z0Z_5 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.didp.regrce3.LdAMones_0 ;
    wire bu_rx_data_0;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.didp.un1_dicLdMones_0_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_1 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.dispString.m49Z0Z_2 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.un24_ce_2 ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.didp.ce_12_3_cascade_ ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.un18_ce ;
    wire oneSecStrb;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.didp.reset_12_1_3 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.LdStens_i_4 ;
    wire \Lab_UT.dictrl.stateZ0Z_2 ;
    wire \Lab_UT.dictrl.N_1460_4 ;
    wire \Lab_UT.dictrl.g2_4 ;
    wire \Lab_UT.dictrl.next_state_4_1_cascade_ ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.LdSones_i_4 ;
    wire \Lab_UT.didp.un1_dicLdSones_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3 ;
    wire \Lab_UT.LdSones ;
    wire bu_rx_data_rdy_0_g;
    wire \Lab_UT.dictrl.g2_5 ;
    wire \Lab_UT.dictrl.g1_3 ;
    wire \Lab_UT.dictrl.g2_5_cascade_ ;
    wire \Lab_UT.dictrl.N_1460_5 ;
    wire \Lab_UT.dictrl.state_ret_12and_0_ns_sn ;
    wire \Lab_UT.dictrl.state_ret_12and_0_ns_rn_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0 ;
    wire \Lab_UT.dictrl.g2_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_2_0_1 ;
    wire \Lab_UT.dictrl.stateZ0Z_1 ;
    wire \Lab_UT.dictrl.N_1460_0 ;
    wire \Lab_UT.dictrl.g2_cascade_ ;
    wire \Lab_UT.dictrl.next_state_0_1 ;
    wire \Lab_UT.dictrl.N_40_3 ;
    wire \Lab_UT.dictrl.N_1105_1_cascade_ ;
    wire \Lab_UT.dictrl.state_i_3_2 ;
    wire \Lab_UT.dictrl.N_79_0 ;
    wire \Lab_UT.dictrl.N_40_5 ;
    wire \Lab_UT.dictrl.g1_2 ;
    wire \Lab_UT.dictrl.N_40_2 ;
    wire \Lab_UT.dictrl.g1_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0 ;
    wire \Lab_UT.state_3 ;
    wire \Lab_UT.dictrl.N_40_1 ;
    wire \Lab_UT.dictrl.g1 ;
    wire \Lab_UT.dictrl.N_97_mux_4 ;
    wire \Lab_UT.dictrl.stateZ0Z_0 ;
    wire \Lab_UT.dictrl.g1_1_1 ;
    wire \Lab_UT.dictrl.m34_4 ;
    wire \Lab_UT.dictrl.N_1106_0 ;
    wire \Lab_UT.dictrl.N_1462_1 ;
    wire \Lab_UT.dictrl.N_1102_1 ;
    wire \Lab_UT.dictrl.g2_1_1 ;
    wire \Lab_UT.dictrl.un1_next_state66_0 ;
    wire \Lab_UT.dictrl.N_1460_1 ;
    wire L3_tx_data_rdy;
    wire \uu2.un1_w_user_cr_0 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.N_75_mux ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.N_14_i_cascade_ ;
    wire \uu2.N_15_i ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ;
    wire \uu2.N_33_cascade_ ;
    wire \uu2.N_14_i ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \INVuu2.w_addr_displaying_0C_net ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \INVuu2.bitmap_212C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.N_194 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.N_197 ;
    wire \Lab_UT.sec1_2 ;
    wire \Lab_UT.sec1_1 ;
    wire \Lab_UT.sec1_3 ;
    wire \Lab_UT.sec1_0 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \INVuu2.bitmap_84C_net ;
    wire \Lab_UT.didp.countrce2.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce2.q_5_2_cascade_ ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.di_Stens_0 ;
    wire bu_rx_data_1;
    wire \Lab_UT.didp.un1_dicLdStens_0 ;
    wire \Lab_UT.didp.countrce2.q_5_1_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.didp.countrce2.un20_qPone ;
    wire \Lab_UT.LdStens ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.didp.countrce2.q_5_3 ;
    wire \Lab_UT.didp.countrce3.ce_12_2_3 ;
    wire \Lab_UT.didp.countrce3.un13_qPone_cascade_ ;
    wire bu_rx_data_2;
    wire \Lab_UT.didp.countrce3.q_5_2_cascade_ ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire bu_rx_data_3;
    wire \Lab_UT.didp.un1_dicLdMones_0 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_3_cascade_ ;
    wire \Lab_UT.di_Mones_3 ;
    wire clk_g;
    wire bu_rx_data_rdy;
    wire rst_g;
    wire bu_rx_data_rdy_0;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__9504),
            .RESETB(N__16951),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__11040,N__11025,N__11220,N__11937,N__12015,N__11199,N__11175,N__11148,N__11109}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__23511,N__14397,N__14439,N__14451,N__13041,N__13059,N__11811,N__11823,N__11874}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__13101,dangling_wire_31,N__12942,dangling_wire_32,N__12915,dangling_wire_33,N__12951,dangling_wire_34,N__13320,dangling_wire_35,N__13137,dangling_wire_36,N__13119}),
            .RCLKE(),
            .RCLK(N__26198),
            .RE(N__16944),
            .WCLKE(N__11840),
            .WCLK(N__26197),
            .WE(N__11844));
    IO_PAD led_obuft_3_iopad (
            .OE(N__26842),
            .DIN(N__26841),
            .DOUT(N__26840),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__26842),
            .PADOUT(N__26841),
            .PADIN(N__26840),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__26833),
            .DIN(N__26832),
            .DOUT(N__26831),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__26833),
            .PADOUT(N__26832),
            .PADIN(N__26831),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__26824),
            .DIN(N__26823),
            .DOUT(N__26822),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__26824),
            .PADOUT(N__26823),
            .PADIN(N__26822),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__26142),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__26815),
            .DIN(N__26814),
            .DOUT(N__26813),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__26815),
            .PADOUT(N__26814),
            .PADIN(N__26813),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__26806),
            .DIN(N__26805),
            .DOUT(N__26804),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__26806),
            .PADOUT(N__26805),
            .PADIN(N__26804),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__26797),
            .DIN(N__26796),
            .DOUT(N__26795),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__26797),
            .PADOUT(N__26796),
            .PADIN(N__26795),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__26788),
            .DIN(N__26787),
            .DOUT(N__26786),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__26788),
            .PADOUT(N__26787),
            .PADIN(N__26786),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__26779),
            .DIN(N__26778),
            .DOUT(N__26777),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__26779),
            .PADOUT(N__26778),
            .PADIN(N__26777),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__26770),
            .DIN(N__26769),
            .DOUT(N__26768),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__26770),
            .PADOUT(N__26769),
            .PADIN(N__26768),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__26761),
            .DIN(N__26760),
            .DOUT(N__26759),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__26761),
            .PADOUT(N__26760),
            .PADIN(N__26759),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__6553 (
            .O(N__26742),
            .I(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ));
    InMux I__6552 (
            .O(N__26739),
            .I(N__26735));
    InMux I__6551 (
            .O(N__26738),
            .I(N__26732));
    LocalMux I__6550 (
            .O(N__26735),
            .I(N__26725));
    LocalMux I__6549 (
            .O(N__26732),
            .I(N__26725));
    InMux I__6548 (
            .O(N__26731),
            .I(N__26719));
    InMux I__6547 (
            .O(N__26730),
            .I(N__26716));
    Span4Mux_v I__6546 (
            .O(N__26725),
            .I(N__26712));
    InMux I__6545 (
            .O(N__26724),
            .I(N__26709));
    InMux I__6544 (
            .O(N__26723),
            .I(N__26706));
    InMux I__6543 (
            .O(N__26722),
            .I(N__26703));
    LocalMux I__6542 (
            .O(N__26719),
            .I(N__26700));
    LocalMux I__6541 (
            .O(N__26716),
            .I(N__26697));
    InMux I__6540 (
            .O(N__26715),
            .I(N__26694));
    IoSpan4Mux I__6539 (
            .O(N__26712),
            .I(N__26690));
    LocalMux I__6538 (
            .O(N__26709),
            .I(N__26681));
    LocalMux I__6537 (
            .O(N__26706),
            .I(N__26681));
    LocalMux I__6536 (
            .O(N__26703),
            .I(N__26672));
    Span4Mux_s2_h I__6535 (
            .O(N__26700),
            .I(N__26672));
    Span4Mux_v I__6534 (
            .O(N__26697),
            .I(N__26672));
    LocalMux I__6533 (
            .O(N__26694),
            .I(N__26672));
    InMux I__6532 (
            .O(N__26693),
            .I(N__26669));
    IoSpan4Mux I__6531 (
            .O(N__26690),
            .I(N__26664));
    InMux I__6530 (
            .O(N__26689),
            .I(N__26655));
    InMux I__6529 (
            .O(N__26688),
            .I(N__26655));
    InMux I__6528 (
            .O(N__26687),
            .I(N__26655));
    InMux I__6527 (
            .O(N__26686),
            .I(N__26655));
    Span4Mux_v I__6526 (
            .O(N__26681),
            .I(N__26652));
    Span4Mux_h I__6525 (
            .O(N__26672),
            .I(N__26644));
    LocalMux I__6524 (
            .O(N__26669),
            .I(N__26644));
    InMux I__6523 (
            .O(N__26668),
            .I(N__26639));
    InMux I__6522 (
            .O(N__26667),
            .I(N__26639));
    Span4Mux_s2_h I__6521 (
            .O(N__26664),
            .I(N__26634));
    LocalMux I__6520 (
            .O(N__26655),
            .I(N__26634));
    Sp12to4 I__6519 (
            .O(N__26652),
            .I(N__26631));
    InMux I__6518 (
            .O(N__26651),
            .I(N__26628));
    InMux I__6517 (
            .O(N__26650),
            .I(N__26623));
    InMux I__6516 (
            .O(N__26649),
            .I(N__26623));
    Span4Mux_v I__6515 (
            .O(N__26644),
            .I(N__26618));
    LocalMux I__6514 (
            .O(N__26639),
            .I(N__26618));
    Span4Mux_h I__6513 (
            .O(N__26634),
            .I(N__26612));
    Span12Mux_s10_h I__6512 (
            .O(N__26631),
            .I(N__26607));
    LocalMux I__6511 (
            .O(N__26628),
            .I(N__26607));
    LocalMux I__6510 (
            .O(N__26623),
            .I(N__26604));
    Span4Mux_h I__6509 (
            .O(N__26618),
            .I(N__26601));
    InMux I__6508 (
            .O(N__26617),
            .I(N__26594));
    InMux I__6507 (
            .O(N__26616),
            .I(N__26594));
    InMux I__6506 (
            .O(N__26615),
            .I(N__26594));
    Span4Mux_h I__6505 (
            .O(N__26612),
            .I(N__26591));
    Odrv12 I__6504 (
            .O(N__26607),
            .I(bu_rx_data_2));
    Odrv4 I__6503 (
            .O(N__26604),
            .I(bu_rx_data_2));
    Odrv4 I__6502 (
            .O(N__26601),
            .I(bu_rx_data_2));
    LocalMux I__6501 (
            .O(N__26594),
            .I(bu_rx_data_2));
    Odrv4 I__6500 (
            .O(N__26591),
            .I(bu_rx_data_2));
    CascadeMux I__6499 (
            .O(N__26580),
            .I(\Lab_UT.didp.countrce3.q_5_2_cascade_ ));
    InMux I__6498 (
            .O(N__26577),
            .I(N__26574));
    LocalMux I__6497 (
            .O(N__26574),
            .I(N__26567));
    CascadeMux I__6496 (
            .O(N__26573),
            .I(N__26563));
    InMux I__6495 (
            .O(N__26572),
            .I(N__26555));
    InMux I__6494 (
            .O(N__26571),
            .I(N__26555));
    InMux I__6493 (
            .O(N__26570),
            .I(N__26555));
    Span4Mux_v I__6492 (
            .O(N__26567),
            .I(N__26552));
    InMux I__6491 (
            .O(N__26566),
            .I(N__26545));
    InMux I__6490 (
            .O(N__26563),
            .I(N__26545));
    InMux I__6489 (
            .O(N__26562),
            .I(N__26545));
    LocalMux I__6488 (
            .O(N__26555),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv4 I__6487 (
            .O(N__26552),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__6486 (
            .O(N__26545),
            .I(\Lab_UT.di_Mones_1 ));
    InMux I__6485 (
            .O(N__26538),
            .I(N__26532));
    InMux I__6484 (
            .O(N__26537),
            .I(N__26532));
    LocalMux I__6483 (
            .O(N__26532),
            .I(N__26524));
    InMux I__6482 (
            .O(N__26531),
            .I(N__26521));
    InMux I__6481 (
            .O(N__26530),
            .I(N__26518));
    InMux I__6480 (
            .O(N__26529),
            .I(N__26511));
    InMux I__6479 (
            .O(N__26528),
            .I(N__26511));
    InMux I__6478 (
            .O(N__26527),
            .I(N__26511));
    Span4Mux_h I__6477 (
            .O(N__26524),
            .I(N__26508));
    LocalMux I__6476 (
            .O(N__26521),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__6475 (
            .O(N__26518),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__6474 (
            .O(N__26511),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__6473 (
            .O(N__26508),
            .I(\Lab_UT.di_Mones_0 ));
    InMux I__6472 (
            .O(N__26499),
            .I(N__26494));
    CascadeMux I__6471 (
            .O(N__26498),
            .I(N__26489));
    CascadeMux I__6470 (
            .O(N__26497),
            .I(N__26486));
    LocalMux I__6469 (
            .O(N__26494),
            .I(N__26483));
    InMux I__6468 (
            .O(N__26493),
            .I(N__26473));
    InMux I__6467 (
            .O(N__26492),
            .I(N__26473));
    InMux I__6466 (
            .O(N__26489),
            .I(N__26473));
    InMux I__6465 (
            .O(N__26486),
            .I(N__26473));
    Span4Mux_h I__6464 (
            .O(N__26483),
            .I(N__26470));
    InMux I__6463 (
            .O(N__26482),
            .I(N__26467));
    LocalMux I__6462 (
            .O(N__26473),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__6461 (
            .O(N__26470),
            .I(\Lab_UT.di_Mones_2 ));
    LocalMux I__6460 (
            .O(N__26467),
            .I(\Lab_UT.di_Mones_2 ));
    InMux I__6459 (
            .O(N__26460),
            .I(N__26452));
    InMux I__6458 (
            .O(N__26459),
            .I(N__26449));
    InMux I__6457 (
            .O(N__26458),
            .I(N__26440));
    InMux I__6456 (
            .O(N__26457),
            .I(N__26440));
    InMux I__6455 (
            .O(N__26456),
            .I(N__26440));
    InMux I__6454 (
            .O(N__26455),
            .I(N__26440));
    LocalMux I__6453 (
            .O(N__26452),
            .I(N__26435));
    LocalMux I__6452 (
            .O(N__26449),
            .I(N__26435));
    LocalMux I__6451 (
            .O(N__26440),
            .I(N__26432));
    Odrv4 I__6450 (
            .O(N__26435),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__6449 (
            .O(N__26432),
            .I(\Lab_UT.LdMones ));
    CascadeMux I__6448 (
            .O(N__26427),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    InMux I__6447 (
            .O(N__26424),
            .I(N__26417));
    InMux I__6446 (
            .O(N__26423),
            .I(N__26414));
    InMux I__6445 (
            .O(N__26422),
            .I(N__26409));
    InMux I__6444 (
            .O(N__26421),
            .I(N__26406));
    InMux I__6443 (
            .O(N__26420),
            .I(N__26403));
    LocalMux I__6442 (
            .O(N__26417),
            .I(N__26398));
    LocalMux I__6441 (
            .O(N__26414),
            .I(N__26398));
    InMux I__6440 (
            .O(N__26413),
            .I(N__26395));
    InMux I__6439 (
            .O(N__26412),
            .I(N__26392));
    LocalMux I__6438 (
            .O(N__26409),
            .I(N__26381));
    LocalMux I__6437 (
            .O(N__26406),
            .I(N__26381));
    LocalMux I__6436 (
            .O(N__26403),
            .I(N__26381));
    Span4Mux_v I__6435 (
            .O(N__26398),
            .I(N__26378));
    LocalMux I__6434 (
            .O(N__26395),
            .I(N__26373));
    LocalMux I__6433 (
            .O(N__26392),
            .I(N__26373));
    CascadeMux I__6432 (
            .O(N__26391),
            .I(N__26367));
    CascadeMux I__6431 (
            .O(N__26390),
            .I(N__26364));
    InMux I__6430 (
            .O(N__26389),
            .I(N__26361));
    InMux I__6429 (
            .O(N__26388),
            .I(N__26355));
    Span4Mux_v I__6428 (
            .O(N__26381),
            .I(N__26350));
    Span4Mux_h I__6427 (
            .O(N__26378),
            .I(N__26350));
    Span4Mux_v I__6426 (
            .O(N__26373),
            .I(N__26345));
    InMux I__6425 (
            .O(N__26372),
            .I(N__26342));
    InMux I__6424 (
            .O(N__26371),
            .I(N__26339));
    InMux I__6423 (
            .O(N__26370),
            .I(N__26332));
    InMux I__6422 (
            .O(N__26367),
            .I(N__26332));
    InMux I__6421 (
            .O(N__26364),
            .I(N__26332));
    LocalMux I__6420 (
            .O(N__26361),
            .I(N__26327));
    InMux I__6419 (
            .O(N__26360),
            .I(N__26320));
    InMux I__6418 (
            .O(N__26359),
            .I(N__26320));
    InMux I__6417 (
            .O(N__26358),
            .I(N__26320));
    LocalMux I__6416 (
            .O(N__26355),
            .I(N__26317));
    Span4Mux_h I__6415 (
            .O(N__26350),
            .I(N__26314));
    InMux I__6414 (
            .O(N__26349),
            .I(N__26309));
    InMux I__6413 (
            .O(N__26348),
            .I(N__26309));
    Span4Mux_h I__6412 (
            .O(N__26345),
            .I(N__26302));
    LocalMux I__6411 (
            .O(N__26342),
            .I(N__26302));
    LocalMux I__6410 (
            .O(N__26339),
            .I(N__26302));
    LocalMux I__6409 (
            .O(N__26332),
            .I(N__26299));
    InMux I__6408 (
            .O(N__26331),
            .I(N__26294));
    InMux I__6407 (
            .O(N__26330),
            .I(N__26294));
    Span4Mux_v I__6406 (
            .O(N__26327),
            .I(N__26289));
    LocalMux I__6405 (
            .O(N__26320),
            .I(N__26289));
    Span12Mux_s8_h I__6404 (
            .O(N__26317),
            .I(N__26282));
    Sp12to4 I__6403 (
            .O(N__26314),
            .I(N__26282));
    LocalMux I__6402 (
            .O(N__26309),
            .I(N__26282));
    Span4Mux_v I__6401 (
            .O(N__26302),
            .I(N__26277));
    Span4Mux_h I__6400 (
            .O(N__26299),
            .I(N__26277));
    LocalMux I__6399 (
            .O(N__26294),
            .I(bu_rx_data_3));
    Odrv4 I__6398 (
            .O(N__26289),
            .I(bu_rx_data_3));
    Odrv12 I__6397 (
            .O(N__26282),
            .I(bu_rx_data_3));
    Odrv4 I__6396 (
            .O(N__26277),
            .I(bu_rx_data_3));
    InMux I__6395 (
            .O(N__26268),
            .I(N__26262));
    InMux I__6394 (
            .O(N__26267),
            .I(N__26262));
    LocalMux I__6393 (
            .O(N__26262),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    CascadeMux I__6392 (
            .O(N__26259),
            .I(N__26253));
    InMux I__6391 (
            .O(N__26258),
            .I(N__26248));
    InMux I__6390 (
            .O(N__26257),
            .I(N__26248));
    InMux I__6389 (
            .O(N__26256),
            .I(N__26243));
    InMux I__6388 (
            .O(N__26253),
            .I(N__26243));
    LocalMux I__6387 (
            .O(N__26248),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    LocalMux I__6386 (
            .O(N__26243),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    CascadeMux I__6385 (
            .O(N__26238),
            .I(\Lab_UT.didp.countrce3.q_5_3_cascade_ ));
    CascadeMux I__6384 (
            .O(N__26235),
            .I(N__26232));
    InMux I__6383 (
            .O(N__26232),
            .I(N__26223));
    InMux I__6382 (
            .O(N__26231),
            .I(N__26223));
    InMux I__6381 (
            .O(N__26230),
            .I(N__26216));
    InMux I__6380 (
            .O(N__26229),
            .I(N__26216));
    InMux I__6379 (
            .O(N__26228),
            .I(N__26216));
    LocalMux I__6378 (
            .O(N__26223),
            .I(N__26213));
    LocalMux I__6377 (
            .O(N__26216),
            .I(N__26208));
    Span4Mux_h I__6376 (
            .O(N__26213),
            .I(N__26208));
    Odrv4 I__6375 (
            .O(N__26208),
            .I(\Lab_UT.di_Mones_3 ));
    ClkMux I__6374 (
            .O(N__26205),
            .I(N__25932));
    ClkMux I__6373 (
            .O(N__26204),
            .I(N__25932));
    ClkMux I__6372 (
            .O(N__26203),
            .I(N__25932));
    ClkMux I__6371 (
            .O(N__26202),
            .I(N__25932));
    ClkMux I__6370 (
            .O(N__26201),
            .I(N__25932));
    ClkMux I__6369 (
            .O(N__26200),
            .I(N__25932));
    ClkMux I__6368 (
            .O(N__26199),
            .I(N__25932));
    ClkMux I__6367 (
            .O(N__26198),
            .I(N__25932));
    ClkMux I__6366 (
            .O(N__26197),
            .I(N__25932));
    ClkMux I__6365 (
            .O(N__26196),
            .I(N__25932));
    ClkMux I__6364 (
            .O(N__26195),
            .I(N__25932));
    ClkMux I__6363 (
            .O(N__26194),
            .I(N__25932));
    ClkMux I__6362 (
            .O(N__26193),
            .I(N__25932));
    ClkMux I__6361 (
            .O(N__26192),
            .I(N__25932));
    ClkMux I__6360 (
            .O(N__26191),
            .I(N__25932));
    ClkMux I__6359 (
            .O(N__26190),
            .I(N__25932));
    ClkMux I__6358 (
            .O(N__26189),
            .I(N__25932));
    ClkMux I__6357 (
            .O(N__26188),
            .I(N__25932));
    ClkMux I__6356 (
            .O(N__26187),
            .I(N__25932));
    ClkMux I__6355 (
            .O(N__26186),
            .I(N__25932));
    ClkMux I__6354 (
            .O(N__26185),
            .I(N__25932));
    ClkMux I__6353 (
            .O(N__26184),
            .I(N__25932));
    ClkMux I__6352 (
            .O(N__26183),
            .I(N__25932));
    ClkMux I__6351 (
            .O(N__26182),
            .I(N__25932));
    ClkMux I__6350 (
            .O(N__26181),
            .I(N__25932));
    ClkMux I__6349 (
            .O(N__26180),
            .I(N__25932));
    ClkMux I__6348 (
            .O(N__26179),
            .I(N__25932));
    ClkMux I__6347 (
            .O(N__26178),
            .I(N__25932));
    ClkMux I__6346 (
            .O(N__26177),
            .I(N__25932));
    ClkMux I__6345 (
            .O(N__26176),
            .I(N__25932));
    ClkMux I__6344 (
            .O(N__26175),
            .I(N__25932));
    ClkMux I__6343 (
            .O(N__26174),
            .I(N__25932));
    ClkMux I__6342 (
            .O(N__26173),
            .I(N__25932));
    ClkMux I__6341 (
            .O(N__26172),
            .I(N__25932));
    ClkMux I__6340 (
            .O(N__26171),
            .I(N__25932));
    ClkMux I__6339 (
            .O(N__26170),
            .I(N__25932));
    ClkMux I__6338 (
            .O(N__26169),
            .I(N__25932));
    ClkMux I__6337 (
            .O(N__26168),
            .I(N__25932));
    ClkMux I__6336 (
            .O(N__26167),
            .I(N__25932));
    ClkMux I__6335 (
            .O(N__26166),
            .I(N__25932));
    ClkMux I__6334 (
            .O(N__26165),
            .I(N__25932));
    ClkMux I__6333 (
            .O(N__26164),
            .I(N__25932));
    ClkMux I__6332 (
            .O(N__26163),
            .I(N__25932));
    ClkMux I__6331 (
            .O(N__26162),
            .I(N__25932));
    ClkMux I__6330 (
            .O(N__26161),
            .I(N__25932));
    ClkMux I__6329 (
            .O(N__26160),
            .I(N__25932));
    ClkMux I__6328 (
            .O(N__26159),
            .I(N__25932));
    ClkMux I__6327 (
            .O(N__26158),
            .I(N__25932));
    ClkMux I__6326 (
            .O(N__26157),
            .I(N__25932));
    ClkMux I__6325 (
            .O(N__26156),
            .I(N__25932));
    ClkMux I__6324 (
            .O(N__26155),
            .I(N__25932));
    ClkMux I__6323 (
            .O(N__26154),
            .I(N__25932));
    ClkMux I__6322 (
            .O(N__26153),
            .I(N__25932));
    ClkMux I__6321 (
            .O(N__26152),
            .I(N__25932));
    ClkMux I__6320 (
            .O(N__26151),
            .I(N__25932));
    ClkMux I__6319 (
            .O(N__26150),
            .I(N__25932));
    ClkMux I__6318 (
            .O(N__26149),
            .I(N__25932));
    ClkMux I__6317 (
            .O(N__26148),
            .I(N__25932));
    ClkMux I__6316 (
            .O(N__26147),
            .I(N__25932));
    ClkMux I__6315 (
            .O(N__26146),
            .I(N__25932));
    ClkMux I__6314 (
            .O(N__26145),
            .I(N__25932));
    ClkMux I__6313 (
            .O(N__26144),
            .I(N__25932));
    ClkMux I__6312 (
            .O(N__26143),
            .I(N__25932));
    ClkMux I__6311 (
            .O(N__26142),
            .I(N__25932));
    ClkMux I__6310 (
            .O(N__26141),
            .I(N__25932));
    ClkMux I__6309 (
            .O(N__26140),
            .I(N__25932));
    ClkMux I__6308 (
            .O(N__26139),
            .I(N__25932));
    ClkMux I__6307 (
            .O(N__26138),
            .I(N__25932));
    ClkMux I__6306 (
            .O(N__26137),
            .I(N__25932));
    ClkMux I__6305 (
            .O(N__26136),
            .I(N__25932));
    ClkMux I__6304 (
            .O(N__26135),
            .I(N__25932));
    ClkMux I__6303 (
            .O(N__26134),
            .I(N__25932));
    ClkMux I__6302 (
            .O(N__26133),
            .I(N__25932));
    ClkMux I__6301 (
            .O(N__26132),
            .I(N__25932));
    ClkMux I__6300 (
            .O(N__26131),
            .I(N__25932));
    ClkMux I__6299 (
            .O(N__26130),
            .I(N__25932));
    ClkMux I__6298 (
            .O(N__26129),
            .I(N__25932));
    ClkMux I__6297 (
            .O(N__26128),
            .I(N__25932));
    ClkMux I__6296 (
            .O(N__26127),
            .I(N__25932));
    ClkMux I__6295 (
            .O(N__26126),
            .I(N__25932));
    ClkMux I__6294 (
            .O(N__26125),
            .I(N__25932));
    ClkMux I__6293 (
            .O(N__26124),
            .I(N__25932));
    ClkMux I__6292 (
            .O(N__26123),
            .I(N__25932));
    ClkMux I__6291 (
            .O(N__26122),
            .I(N__25932));
    ClkMux I__6290 (
            .O(N__26121),
            .I(N__25932));
    ClkMux I__6289 (
            .O(N__26120),
            .I(N__25932));
    ClkMux I__6288 (
            .O(N__26119),
            .I(N__25932));
    ClkMux I__6287 (
            .O(N__26118),
            .I(N__25932));
    ClkMux I__6286 (
            .O(N__26117),
            .I(N__25932));
    ClkMux I__6285 (
            .O(N__26116),
            .I(N__25932));
    ClkMux I__6284 (
            .O(N__26115),
            .I(N__25932));
    GlobalMux I__6283 (
            .O(N__25932),
            .I(N__25929));
    gio2CtrlBuf I__6282 (
            .O(N__25929),
            .I(clk_g));
    InMux I__6281 (
            .O(N__25926),
            .I(N__25919));
    InMux I__6280 (
            .O(N__25925),
            .I(N__25919));
    InMux I__6279 (
            .O(N__25924),
            .I(N__25915));
    LocalMux I__6278 (
            .O(N__25919),
            .I(N__25912));
    InMux I__6277 (
            .O(N__25918),
            .I(N__25909));
    LocalMux I__6276 (
            .O(N__25915),
            .I(N__25906));
    Span4Mux_v I__6275 (
            .O(N__25912),
            .I(N__25903));
    LocalMux I__6274 (
            .O(N__25909),
            .I(N__25900));
    Span4Mux_s3_h I__6273 (
            .O(N__25906),
            .I(N__25896));
    Sp12to4 I__6272 (
            .O(N__25903),
            .I(N__25891));
    Span12Mux_s1_h I__6271 (
            .O(N__25900),
            .I(N__25891));
    InMux I__6270 (
            .O(N__25899),
            .I(N__25888));
    Odrv4 I__6269 (
            .O(N__25896),
            .I(bu_rx_data_rdy));
    Odrv12 I__6268 (
            .O(N__25891),
            .I(bu_rx_data_rdy));
    LocalMux I__6267 (
            .O(N__25888),
            .I(bu_rx_data_rdy));
    InMux I__6266 (
            .O(N__25881),
            .I(N__25869));
    InMux I__6265 (
            .O(N__25880),
            .I(N__25866));
    InMux I__6264 (
            .O(N__25879),
            .I(N__25863));
    InMux I__6263 (
            .O(N__25878),
            .I(N__25860));
    InMux I__6262 (
            .O(N__25877),
            .I(N__25855));
    InMux I__6261 (
            .O(N__25876),
            .I(N__25855));
    InMux I__6260 (
            .O(N__25875),
            .I(N__25852));
    InMux I__6259 (
            .O(N__25874),
            .I(N__25849));
    InMux I__6258 (
            .O(N__25873),
            .I(N__25846));
    InMux I__6257 (
            .O(N__25872),
            .I(N__25843));
    LocalMux I__6256 (
            .O(N__25869),
            .I(N__25796));
    LocalMux I__6255 (
            .O(N__25866),
            .I(N__25793));
    LocalMux I__6254 (
            .O(N__25863),
            .I(N__25790));
    LocalMux I__6253 (
            .O(N__25860),
            .I(N__25787));
    LocalMux I__6252 (
            .O(N__25855),
            .I(N__25784));
    LocalMux I__6251 (
            .O(N__25852),
            .I(N__25781));
    LocalMux I__6250 (
            .O(N__25849),
            .I(N__25762));
    LocalMux I__6249 (
            .O(N__25846),
            .I(N__25759));
    LocalMux I__6248 (
            .O(N__25843),
            .I(N__25756));
    SRMux I__6247 (
            .O(N__25842),
            .I(N__25617));
    SRMux I__6246 (
            .O(N__25841),
            .I(N__25617));
    SRMux I__6245 (
            .O(N__25840),
            .I(N__25617));
    SRMux I__6244 (
            .O(N__25839),
            .I(N__25617));
    SRMux I__6243 (
            .O(N__25838),
            .I(N__25617));
    SRMux I__6242 (
            .O(N__25837),
            .I(N__25617));
    SRMux I__6241 (
            .O(N__25836),
            .I(N__25617));
    SRMux I__6240 (
            .O(N__25835),
            .I(N__25617));
    SRMux I__6239 (
            .O(N__25834),
            .I(N__25617));
    SRMux I__6238 (
            .O(N__25833),
            .I(N__25617));
    SRMux I__6237 (
            .O(N__25832),
            .I(N__25617));
    SRMux I__6236 (
            .O(N__25831),
            .I(N__25617));
    SRMux I__6235 (
            .O(N__25830),
            .I(N__25617));
    SRMux I__6234 (
            .O(N__25829),
            .I(N__25617));
    SRMux I__6233 (
            .O(N__25828),
            .I(N__25617));
    SRMux I__6232 (
            .O(N__25827),
            .I(N__25617));
    SRMux I__6231 (
            .O(N__25826),
            .I(N__25617));
    SRMux I__6230 (
            .O(N__25825),
            .I(N__25617));
    SRMux I__6229 (
            .O(N__25824),
            .I(N__25617));
    SRMux I__6228 (
            .O(N__25823),
            .I(N__25617));
    SRMux I__6227 (
            .O(N__25822),
            .I(N__25617));
    SRMux I__6226 (
            .O(N__25821),
            .I(N__25617));
    SRMux I__6225 (
            .O(N__25820),
            .I(N__25617));
    SRMux I__6224 (
            .O(N__25819),
            .I(N__25617));
    SRMux I__6223 (
            .O(N__25818),
            .I(N__25617));
    SRMux I__6222 (
            .O(N__25817),
            .I(N__25617));
    SRMux I__6221 (
            .O(N__25816),
            .I(N__25617));
    SRMux I__6220 (
            .O(N__25815),
            .I(N__25617));
    SRMux I__6219 (
            .O(N__25814),
            .I(N__25617));
    SRMux I__6218 (
            .O(N__25813),
            .I(N__25617));
    SRMux I__6217 (
            .O(N__25812),
            .I(N__25617));
    SRMux I__6216 (
            .O(N__25811),
            .I(N__25617));
    SRMux I__6215 (
            .O(N__25810),
            .I(N__25617));
    SRMux I__6214 (
            .O(N__25809),
            .I(N__25617));
    SRMux I__6213 (
            .O(N__25808),
            .I(N__25617));
    SRMux I__6212 (
            .O(N__25807),
            .I(N__25617));
    SRMux I__6211 (
            .O(N__25806),
            .I(N__25617));
    SRMux I__6210 (
            .O(N__25805),
            .I(N__25617));
    SRMux I__6209 (
            .O(N__25804),
            .I(N__25617));
    SRMux I__6208 (
            .O(N__25803),
            .I(N__25617));
    SRMux I__6207 (
            .O(N__25802),
            .I(N__25617));
    SRMux I__6206 (
            .O(N__25801),
            .I(N__25617));
    SRMux I__6205 (
            .O(N__25800),
            .I(N__25617));
    SRMux I__6204 (
            .O(N__25799),
            .I(N__25617));
    Glb2LocalMux I__6203 (
            .O(N__25796),
            .I(N__25617));
    Glb2LocalMux I__6202 (
            .O(N__25793),
            .I(N__25617));
    Glb2LocalMux I__6201 (
            .O(N__25790),
            .I(N__25617));
    Glb2LocalMux I__6200 (
            .O(N__25787),
            .I(N__25617));
    Glb2LocalMux I__6199 (
            .O(N__25784),
            .I(N__25617));
    Glb2LocalMux I__6198 (
            .O(N__25781),
            .I(N__25617));
    SRMux I__6197 (
            .O(N__25780),
            .I(N__25617));
    SRMux I__6196 (
            .O(N__25779),
            .I(N__25617));
    SRMux I__6195 (
            .O(N__25778),
            .I(N__25617));
    SRMux I__6194 (
            .O(N__25777),
            .I(N__25617));
    SRMux I__6193 (
            .O(N__25776),
            .I(N__25617));
    SRMux I__6192 (
            .O(N__25775),
            .I(N__25617));
    SRMux I__6191 (
            .O(N__25774),
            .I(N__25617));
    SRMux I__6190 (
            .O(N__25773),
            .I(N__25617));
    SRMux I__6189 (
            .O(N__25772),
            .I(N__25617));
    SRMux I__6188 (
            .O(N__25771),
            .I(N__25617));
    SRMux I__6187 (
            .O(N__25770),
            .I(N__25617));
    SRMux I__6186 (
            .O(N__25769),
            .I(N__25617));
    SRMux I__6185 (
            .O(N__25768),
            .I(N__25617));
    SRMux I__6184 (
            .O(N__25767),
            .I(N__25617));
    SRMux I__6183 (
            .O(N__25766),
            .I(N__25617));
    SRMux I__6182 (
            .O(N__25765),
            .I(N__25617));
    Glb2LocalMux I__6181 (
            .O(N__25762),
            .I(N__25617));
    Glb2LocalMux I__6180 (
            .O(N__25759),
            .I(N__25617));
    Glb2LocalMux I__6179 (
            .O(N__25756),
            .I(N__25617));
    GlobalMux I__6178 (
            .O(N__25617),
            .I(N__25614));
    gio2CtrlBuf I__6177 (
            .O(N__25614),
            .I(rst_g));
    IoInMux I__6176 (
            .O(N__25611),
            .I(N__25608));
    LocalMux I__6175 (
            .O(N__25608),
            .I(bu_rx_data_rdy_0));
    CascadeMux I__6174 (
            .O(N__25605),
            .I(\Lab_UT.didp.countrce2.un13_qPone_cascade_ ));
    CascadeMux I__6173 (
            .O(N__25602),
            .I(\Lab_UT.didp.countrce2.q_5_2_cascade_ ));
    CascadeMux I__6172 (
            .O(N__25599),
            .I(N__25595));
    InMux I__6171 (
            .O(N__25598),
            .I(N__25590));
    InMux I__6170 (
            .O(N__25595),
            .I(N__25590));
    LocalMux I__6169 (
            .O(N__25590),
            .I(N__25583));
    InMux I__6168 (
            .O(N__25589),
            .I(N__25580));
    InMux I__6167 (
            .O(N__25588),
            .I(N__25577));
    InMux I__6166 (
            .O(N__25587),
            .I(N__25572));
    InMux I__6165 (
            .O(N__25586),
            .I(N__25572));
    Span4Mux_h I__6164 (
            .O(N__25583),
            .I(N__25569));
    LocalMux I__6163 (
            .O(N__25580),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__6162 (
            .O(N__25577),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__6161 (
            .O(N__25572),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv4 I__6160 (
            .O(N__25569),
            .I(\Lab_UT.di_Stens_2 ));
    InMux I__6159 (
            .O(N__25560),
            .I(N__25550));
    InMux I__6158 (
            .O(N__25559),
            .I(N__25543));
    InMux I__6157 (
            .O(N__25558),
            .I(N__25543));
    InMux I__6156 (
            .O(N__25557),
            .I(N__25543));
    InMux I__6155 (
            .O(N__25556),
            .I(N__25534));
    InMux I__6154 (
            .O(N__25555),
            .I(N__25534));
    InMux I__6153 (
            .O(N__25554),
            .I(N__25534));
    InMux I__6152 (
            .O(N__25553),
            .I(N__25534));
    LocalMux I__6151 (
            .O(N__25550),
            .I(N__25531));
    LocalMux I__6150 (
            .O(N__25543),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__6149 (
            .O(N__25534),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv4 I__6148 (
            .O(N__25531),
            .I(\Lab_UT.di_Stens_0 ));
    InMux I__6147 (
            .O(N__25524),
            .I(N__25516));
    InMux I__6146 (
            .O(N__25523),
            .I(N__25513));
    InMux I__6145 (
            .O(N__25522),
            .I(N__25510));
    InMux I__6144 (
            .O(N__25521),
            .I(N__25507));
    InMux I__6143 (
            .O(N__25520),
            .I(N__25504));
    InMux I__6142 (
            .O(N__25519),
            .I(N__25498));
    LocalMux I__6141 (
            .O(N__25516),
            .I(N__25490));
    LocalMux I__6140 (
            .O(N__25513),
            .I(N__25485));
    LocalMux I__6139 (
            .O(N__25510),
            .I(N__25485));
    LocalMux I__6138 (
            .O(N__25507),
            .I(N__25482));
    LocalMux I__6137 (
            .O(N__25504),
            .I(N__25478));
    InMux I__6136 (
            .O(N__25503),
            .I(N__25475));
    InMux I__6135 (
            .O(N__25502),
            .I(N__25470));
    InMux I__6134 (
            .O(N__25501),
            .I(N__25470));
    LocalMux I__6133 (
            .O(N__25498),
            .I(N__25467));
    InMux I__6132 (
            .O(N__25497),
            .I(N__25458));
    InMux I__6131 (
            .O(N__25496),
            .I(N__25458));
    InMux I__6130 (
            .O(N__25495),
            .I(N__25458));
    InMux I__6129 (
            .O(N__25494),
            .I(N__25458));
    InMux I__6128 (
            .O(N__25493),
            .I(N__25453));
    Span4Mux_v I__6127 (
            .O(N__25490),
            .I(N__25450));
    Span4Mux_v I__6126 (
            .O(N__25485),
            .I(N__25447));
    Span4Mux_v I__6125 (
            .O(N__25482),
            .I(N__25444));
    InMux I__6124 (
            .O(N__25481),
            .I(N__25441));
    Span4Mux_h I__6123 (
            .O(N__25478),
            .I(N__25434));
    LocalMux I__6122 (
            .O(N__25475),
            .I(N__25434));
    LocalMux I__6121 (
            .O(N__25470),
            .I(N__25431));
    Span4Mux_v I__6120 (
            .O(N__25467),
            .I(N__25426));
    LocalMux I__6119 (
            .O(N__25458),
            .I(N__25426));
    InMux I__6118 (
            .O(N__25457),
            .I(N__25421));
    InMux I__6117 (
            .O(N__25456),
            .I(N__25421));
    LocalMux I__6116 (
            .O(N__25453),
            .I(N__25418));
    Sp12to4 I__6115 (
            .O(N__25450),
            .I(N__25409));
    Sp12to4 I__6114 (
            .O(N__25447),
            .I(N__25409));
    Sp12to4 I__6113 (
            .O(N__25444),
            .I(N__25409));
    LocalMux I__6112 (
            .O(N__25441),
            .I(N__25409));
    CascadeMux I__6111 (
            .O(N__25440),
            .I(N__25405));
    CascadeMux I__6110 (
            .O(N__25439),
            .I(N__25402));
    Span4Mux_h I__6109 (
            .O(N__25434),
            .I(N__25399));
    Span4Mux_v I__6108 (
            .O(N__25431),
            .I(N__25394));
    Span4Mux_h I__6107 (
            .O(N__25426),
            .I(N__25394));
    LocalMux I__6106 (
            .O(N__25421),
            .I(N__25389));
    Span12Mux_v I__6105 (
            .O(N__25418),
            .I(N__25389));
    Span12Mux_s10_h I__6104 (
            .O(N__25409),
            .I(N__25386));
    InMux I__6103 (
            .O(N__25408),
            .I(N__25379));
    InMux I__6102 (
            .O(N__25405),
            .I(N__25379));
    InMux I__6101 (
            .O(N__25402),
            .I(N__25379));
    Span4Mux_v I__6100 (
            .O(N__25399),
            .I(N__25374));
    Span4Mux_h I__6099 (
            .O(N__25394),
            .I(N__25374));
    Odrv12 I__6098 (
            .O(N__25389),
            .I(bu_rx_data_1));
    Odrv12 I__6097 (
            .O(N__25386),
            .I(bu_rx_data_1));
    LocalMux I__6096 (
            .O(N__25379),
            .I(bu_rx_data_1));
    Odrv4 I__6095 (
            .O(N__25374),
            .I(bu_rx_data_1));
    InMux I__6094 (
            .O(N__25365),
            .I(N__25357));
    InMux I__6093 (
            .O(N__25364),
            .I(N__25357));
    InMux I__6092 (
            .O(N__25363),
            .I(N__25354));
    InMux I__6091 (
            .O(N__25362),
            .I(N__25351));
    LocalMux I__6090 (
            .O(N__25357),
            .I(N__25344));
    LocalMux I__6089 (
            .O(N__25354),
            .I(N__25344));
    LocalMux I__6088 (
            .O(N__25351),
            .I(N__25344));
    Span4Mux_s1_h I__6087 (
            .O(N__25344),
            .I(N__25341));
    Odrv4 I__6086 (
            .O(N__25341),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    CascadeMux I__6085 (
            .O(N__25338),
            .I(\Lab_UT.didp.countrce2.q_5_1_cascade_ ));
    CascadeMux I__6084 (
            .O(N__25335),
            .I(N__25332));
    InMux I__6083 (
            .O(N__25332),
            .I(N__25324));
    InMux I__6082 (
            .O(N__25331),
            .I(N__25324));
    InMux I__6081 (
            .O(N__25330),
            .I(N__25321));
    InMux I__6080 (
            .O(N__25329),
            .I(N__25318));
    LocalMux I__6079 (
            .O(N__25324),
            .I(N__25313));
    LocalMux I__6078 (
            .O(N__25321),
            .I(N__25313));
    LocalMux I__6077 (
            .O(N__25318),
            .I(N__25310));
    Span4Mux_s1_h I__6076 (
            .O(N__25313),
            .I(N__25307));
    Odrv4 I__6075 (
            .O(N__25310),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    Odrv4 I__6074 (
            .O(N__25307),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    CascadeMux I__6073 (
            .O(N__25302),
            .I(N__25293));
    InMux I__6072 (
            .O(N__25301),
            .I(N__25284));
    InMux I__6071 (
            .O(N__25300),
            .I(N__25284));
    InMux I__6070 (
            .O(N__25299),
            .I(N__25284));
    InMux I__6069 (
            .O(N__25298),
            .I(N__25284));
    InMux I__6068 (
            .O(N__25297),
            .I(N__25277));
    InMux I__6067 (
            .O(N__25296),
            .I(N__25277));
    InMux I__6066 (
            .O(N__25293),
            .I(N__25277));
    LocalMux I__6065 (
            .O(N__25284),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__6064 (
            .O(N__25277),
            .I(\Lab_UT.di_Stens_1 ));
    InMux I__6063 (
            .O(N__25272),
            .I(N__25269));
    LocalMux I__6062 (
            .O(N__25269),
            .I(\Lab_UT.didp.countrce2.un20_qPone ));
    CascadeMux I__6061 (
            .O(N__25266),
            .I(N__25261));
    CascadeMux I__6060 (
            .O(N__25265),
            .I(N__25257));
    InMux I__6059 (
            .O(N__25264),
            .I(N__25252));
    InMux I__6058 (
            .O(N__25261),
            .I(N__25252));
    InMux I__6057 (
            .O(N__25260),
            .I(N__25249));
    InMux I__6056 (
            .O(N__25257),
            .I(N__25246));
    LocalMux I__6055 (
            .O(N__25252),
            .I(N__25241));
    LocalMux I__6054 (
            .O(N__25249),
            .I(N__25241));
    LocalMux I__6053 (
            .O(N__25246),
            .I(N__25238));
    Span4Mux_v I__6052 (
            .O(N__25241),
            .I(N__25235));
    Span4Mux_s0_h I__6051 (
            .O(N__25238),
            .I(N__25232));
    Odrv4 I__6050 (
            .O(N__25235),
            .I(\Lab_UT.LdStens ));
    Odrv4 I__6049 (
            .O(N__25232),
            .I(\Lab_UT.LdStens ));
    CascadeMux I__6048 (
            .O(N__25227),
            .I(N__25223));
    CascadeMux I__6047 (
            .O(N__25226),
            .I(N__25217));
    InMux I__6046 (
            .O(N__25223),
            .I(N__25212));
    InMux I__6045 (
            .O(N__25222),
            .I(N__25212));
    InMux I__6044 (
            .O(N__25221),
            .I(N__25209));
    InMux I__6043 (
            .O(N__25220),
            .I(N__25206));
    InMux I__6042 (
            .O(N__25217),
            .I(N__25203));
    LocalMux I__6041 (
            .O(N__25212),
            .I(N__25200));
    LocalMux I__6040 (
            .O(N__25209),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__6039 (
            .O(N__25206),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__6038 (
            .O(N__25203),
            .I(\Lab_UT.di_Stens_3 ));
    Odrv12 I__6037 (
            .O(N__25200),
            .I(\Lab_UT.di_Stens_3 ));
    InMux I__6036 (
            .O(N__25191),
            .I(N__25188));
    LocalMux I__6035 (
            .O(N__25188),
            .I(\Lab_UT.didp.countrce2.q_5_3 ));
    InMux I__6034 (
            .O(N__25185),
            .I(N__25176));
    InMux I__6033 (
            .O(N__25184),
            .I(N__25176));
    InMux I__6032 (
            .O(N__25183),
            .I(N__25176));
    LocalMux I__6031 (
            .O(N__25176),
            .I(\Lab_UT.didp.countrce3.ce_12_2_3 ));
    CascadeMux I__6030 (
            .O(N__25173),
            .I(N__25164));
    InMux I__6029 (
            .O(N__25172),
            .I(N__25157));
    InMux I__6028 (
            .O(N__25171),
            .I(N__25157));
    InMux I__6027 (
            .O(N__25170),
            .I(N__25154));
    CascadeMux I__6026 (
            .O(N__25169),
            .I(N__25151));
    CascadeMux I__6025 (
            .O(N__25168),
            .I(N__25148));
    InMux I__6024 (
            .O(N__25167),
            .I(N__25143));
    InMux I__6023 (
            .O(N__25164),
            .I(N__25143));
    CascadeMux I__6022 (
            .O(N__25163),
            .I(N__25140));
    CascadeMux I__6021 (
            .O(N__25162),
            .I(N__25137));
    LocalMux I__6020 (
            .O(N__25157),
            .I(N__25131));
    LocalMux I__6019 (
            .O(N__25154),
            .I(N__25131));
    InMux I__6018 (
            .O(N__25151),
            .I(N__25126));
    InMux I__6017 (
            .O(N__25148),
            .I(N__25126));
    LocalMux I__6016 (
            .O(N__25143),
            .I(N__25123));
    InMux I__6015 (
            .O(N__25140),
            .I(N__25116));
    InMux I__6014 (
            .O(N__25137),
            .I(N__25116));
    InMux I__6013 (
            .O(N__25136),
            .I(N__25116));
    Span4Mux_s3_h I__6012 (
            .O(N__25131),
            .I(N__25113));
    LocalMux I__6011 (
            .O(N__25126),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__6010 (
            .O(N__25123),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__6009 (
            .O(N__25116),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__6008 (
            .O(N__25113),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CascadeMux I__6007 (
            .O(N__25104),
            .I(N__25097));
    InMux I__6006 (
            .O(N__25103),
            .I(N__25094));
    InMux I__6005 (
            .O(N__25102),
            .I(N__25091));
    InMux I__6004 (
            .O(N__25101),
            .I(N__25080));
    InMux I__6003 (
            .O(N__25100),
            .I(N__25080));
    InMux I__6002 (
            .O(N__25097),
            .I(N__25080));
    LocalMux I__6001 (
            .O(N__25094),
            .I(N__25071));
    LocalMux I__6000 (
            .O(N__25091),
            .I(N__25071));
    InMux I__5999 (
            .O(N__25090),
            .I(N__25068));
    InMux I__5998 (
            .O(N__25089),
            .I(N__25061));
    InMux I__5997 (
            .O(N__25088),
            .I(N__25061));
    InMux I__5996 (
            .O(N__25087),
            .I(N__25061));
    LocalMux I__5995 (
            .O(N__25080),
            .I(N__25058));
    InMux I__5994 (
            .O(N__25079),
            .I(N__25053));
    InMux I__5993 (
            .O(N__25078),
            .I(N__25053));
    InMux I__5992 (
            .O(N__25077),
            .I(N__25048));
    InMux I__5991 (
            .O(N__25076),
            .I(N__25048));
    Span4Mux_s3_h I__5990 (
            .O(N__25071),
            .I(N__25043));
    LocalMux I__5989 (
            .O(N__25068),
            .I(N__25043));
    LocalMux I__5988 (
            .O(N__25061),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__5987 (
            .O(N__25058),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__5986 (
            .O(N__25053),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__5985 (
            .O(N__25048),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__5984 (
            .O(N__25043),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__5983 (
            .O(N__25032),
            .I(N__25021));
    InMux I__5982 (
            .O(N__25031),
            .I(N__25021));
    InMux I__5981 (
            .O(N__25030),
            .I(N__25021));
    InMux I__5980 (
            .O(N__25029),
            .I(N__25014));
    InMux I__5979 (
            .O(N__25028),
            .I(N__25014));
    LocalMux I__5978 (
            .O(N__25021),
            .I(N__25011));
    InMux I__5977 (
            .O(N__25020),
            .I(N__25008));
    InMux I__5976 (
            .O(N__25019),
            .I(N__25005));
    LocalMux I__5975 (
            .O(N__25014),
            .I(N__25002));
    Span4Mux_s3_h I__5974 (
            .O(N__25011),
            .I(N__24995));
    LocalMux I__5973 (
            .O(N__25008),
            .I(N__24992));
    LocalMux I__5972 (
            .O(N__25005),
            .I(N__24989));
    Span4Mux_s2_v I__5971 (
            .O(N__25002),
            .I(N__24986));
    InMux I__5970 (
            .O(N__25001),
            .I(N__24977));
    InMux I__5969 (
            .O(N__25000),
            .I(N__24977));
    InMux I__5968 (
            .O(N__24999),
            .I(N__24977));
    InMux I__5967 (
            .O(N__24998),
            .I(N__24977));
    Odrv4 I__5966 (
            .O(N__24995),
            .I(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ));
    Odrv4 I__5965 (
            .O(N__24992),
            .I(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ));
    Odrv4 I__5964 (
            .O(N__24989),
            .I(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ));
    Odrv4 I__5963 (
            .O(N__24986),
            .I(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ));
    LocalMux I__5962 (
            .O(N__24977),
            .I(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ));
    CascadeMux I__5961 (
            .O(N__24966),
            .I(\uu2.N_33_cascade_ ));
    InMux I__5960 (
            .O(N__24963),
            .I(N__24960));
    LocalMux I__5959 (
            .O(N__24960),
            .I(\uu2.N_14_i ));
    InMux I__5958 (
            .O(N__24957),
            .I(N__24947));
    InMux I__5957 (
            .O(N__24956),
            .I(N__24947));
    InMux I__5956 (
            .O(N__24955),
            .I(N__24947));
    CascadeMux I__5955 (
            .O(N__24954),
            .I(N__24944));
    LocalMux I__5954 (
            .O(N__24947),
            .I(N__24941));
    InMux I__5953 (
            .O(N__24944),
            .I(N__24938));
    Span4Mux_s0_v I__5952 (
            .O(N__24941),
            .I(N__24933));
    LocalMux I__5951 (
            .O(N__24938),
            .I(N__24930));
    InMux I__5950 (
            .O(N__24937),
            .I(N__24927));
    InMux I__5949 (
            .O(N__24936),
            .I(N__24924));
    Span4Mux_h I__5948 (
            .O(N__24933),
            .I(N__24921));
    Span4Mux_s1_v I__5947 (
            .O(N__24930),
            .I(N__24918));
    LocalMux I__5946 (
            .O(N__24927),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__5945 (
            .O(N__24924),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__5944 (
            .O(N__24921),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__5943 (
            .O(N__24918),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__5942 (
            .O(N__24909),
            .I(N__24906));
    LocalMux I__5941 (
            .O(N__24906),
            .I(N__24903));
    Odrv12 I__5940 (
            .O(N__24903),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__5939 (
            .O(N__24900),
            .I(N__24897));
    LocalMux I__5938 (
            .O(N__24897),
            .I(\uu2.bitmapZ0Z_180 ));
    InMux I__5937 (
            .O(N__24894),
            .I(N__24886));
    InMux I__5936 (
            .O(N__24893),
            .I(N__24883));
    InMux I__5935 (
            .O(N__24892),
            .I(N__24878));
    InMux I__5934 (
            .O(N__24891),
            .I(N__24878));
    InMux I__5933 (
            .O(N__24890),
            .I(N__24875));
    InMux I__5932 (
            .O(N__24889),
            .I(N__24872));
    LocalMux I__5931 (
            .O(N__24886),
            .I(N__24869));
    LocalMux I__5930 (
            .O(N__24883),
            .I(N__24864));
    LocalMux I__5929 (
            .O(N__24878),
            .I(N__24864));
    LocalMux I__5928 (
            .O(N__24875),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__5927 (
            .O(N__24872),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__5926 (
            .O(N__24869),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv12 I__5925 (
            .O(N__24864),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    InMux I__5924 (
            .O(N__24855),
            .I(N__24852));
    LocalMux I__5923 (
            .O(N__24852),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__5922 (
            .O(N__24849),
            .I(N__24846));
    LocalMux I__5921 (
            .O(N__24846),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__5920 (
            .O(N__24843),
            .I(N__24840));
    LocalMux I__5919 (
            .O(N__24840),
            .I(\uu2.N_194 ));
    InMux I__5918 (
            .O(N__24837),
            .I(N__24834));
    LocalMux I__5917 (
            .O(N__24834),
            .I(N__24831));
    Odrv4 I__5916 (
            .O(N__24831),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__5915 (
            .O(N__24828),
            .I(N__24825));
    LocalMux I__5914 (
            .O(N__24825),
            .I(N__24821));
    InMux I__5913 (
            .O(N__24824),
            .I(N__24817));
    Span4Mux_v I__5912 (
            .O(N__24821),
            .I(N__24814));
    InMux I__5911 (
            .O(N__24820),
            .I(N__24811));
    LocalMux I__5910 (
            .O(N__24817),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__5909 (
            .O(N__24814),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__5908 (
            .O(N__24811),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__5907 (
            .O(N__24804),
            .I(N__24801));
    LocalMux I__5906 (
            .O(N__24801),
            .I(N__24798));
    Odrv4 I__5905 (
            .O(N__24798),
            .I(\uu2.N_197 ));
    CascadeMux I__5904 (
            .O(N__24795),
            .I(N__24791));
    CascadeMux I__5903 (
            .O(N__24794),
            .I(N__24788));
    InMux I__5902 (
            .O(N__24791),
            .I(N__24779));
    InMux I__5901 (
            .O(N__24788),
            .I(N__24779));
    InMux I__5900 (
            .O(N__24787),
            .I(N__24776));
    InMux I__5899 (
            .O(N__24786),
            .I(N__24769));
    InMux I__5898 (
            .O(N__24785),
            .I(N__24769));
    InMux I__5897 (
            .O(N__24784),
            .I(N__24769));
    LocalMux I__5896 (
            .O(N__24779),
            .I(N__24765));
    LocalMux I__5895 (
            .O(N__24776),
            .I(N__24760));
    LocalMux I__5894 (
            .O(N__24769),
            .I(N__24760));
    InMux I__5893 (
            .O(N__24768),
            .I(N__24757));
    Span4Mux_s2_h I__5892 (
            .O(N__24765),
            .I(N__24754));
    Span4Mux_s2_h I__5891 (
            .O(N__24760),
            .I(N__24751));
    LocalMux I__5890 (
            .O(N__24757),
            .I(N__24748));
    Odrv4 I__5889 (
            .O(N__24754),
            .I(\Lab_UT.sec1_2 ));
    Odrv4 I__5888 (
            .O(N__24751),
            .I(\Lab_UT.sec1_2 ));
    Odrv12 I__5887 (
            .O(N__24748),
            .I(\Lab_UT.sec1_2 ));
    InMux I__5886 (
            .O(N__24741),
            .I(N__24736));
    InMux I__5885 (
            .O(N__24740),
            .I(N__24731));
    InMux I__5884 (
            .O(N__24739),
            .I(N__24731));
    LocalMux I__5883 (
            .O(N__24736),
            .I(N__24727));
    LocalMux I__5882 (
            .O(N__24731),
            .I(N__24724));
    CascadeMux I__5881 (
            .O(N__24730),
            .I(N__24720));
    Span4Mux_h I__5880 (
            .O(N__24727),
            .I(N__24713));
    Span4Mux_s0_h I__5879 (
            .O(N__24724),
            .I(N__24713));
    InMux I__5878 (
            .O(N__24723),
            .I(N__24710));
    InMux I__5877 (
            .O(N__24720),
            .I(N__24703));
    InMux I__5876 (
            .O(N__24719),
            .I(N__24703));
    InMux I__5875 (
            .O(N__24718),
            .I(N__24703));
    Odrv4 I__5874 (
            .O(N__24713),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__5873 (
            .O(N__24710),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__5872 (
            .O(N__24703),
            .I(\Lab_UT.sec1_1 ));
    CascadeMux I__5871 (
            .O(N__24696),
            .I(N__24688));
    CascadeMux I__5870 (
            .O(N__24695),
            .I(N__24684));
    CascadeMux I__5869 (
            .O(N__24694),
            .I(N__24681));
    CascadeMux I__5868 (
            .O(N__24693),
            .I(N__24678));
    InMux I__5867 (
            .O(N__24692),
            .I(N__24673));
    InMux I__5866 (
            .O(N__24691),
            .I(N__24673));
    InMux I__5865 (
            .O(N__24688),
            .I(N__24670));
    InMux I__5864 (
            .O(N__24687),
            .I(N__24663));
    InMux I__5863 (
            .O(N__24684),
            .I(N__24663));
    InMux I__5862 (
            .O(N__24681),
            .I(N__24663));
    InMux I__5861 (
            .O(N__24678),
            .I(N__24660));
    LocalMux I__5860 (
            .O(N__24673),
            .I(N__24657));
    LocalMux I__5859 (
            .O(N__24670),
            .I(N__24652));
    LocalMux I__5858 (
            .O(N__24663),
            .I(N__24652));
    LocalMux I__5857 (
            .O(N__24660),
            .I(N__24649));
    Span12Mux_s4_h I__5856 (
            .O(N__24657),
            .I(N__24646));
    Span4Mux_s3_h I__5855 (
            .O(N__24652),
            .I(N__24641));
    Span4Mux_s3_v I__5854 (
            .O(N__24649),
            .I(N__24641));
    Odrv12 I__5853 (
            .O(N__24646),
            .I(\Lab_UT.sec1_3 ));
    Odrv4 I__5852 (
            .O(N__24641),
            .I(\Lab_UT.sec1_3 ));
    InMux I__5851 (
            .O(N__24636),
            .I(N__24633));
    LocalMux I__5850 (
            .O(N__24633),
            .I(N__24628));
    InMux I__5849 (
            .O(N__24632),
            .I(N__24623));
    InMux I__5848 (
            .O(N__24631),
            .I(N__24623));
    Span4Mux_v I__5847 (
            .O(N__24628),
            .I(N__24616));
    LocalMux I__5846 (
            .O(N__24623),
            .I(N__24613));
    InMux I__5845 (
            .O(N__24622),
            .I(N__24610));
    InMux I__5844 (
            .O(N__24621),
            .I(N__24603));
    InMux I__5843 (
            .O(N__24620),
            .I(N__24603));
    InMux I__5842 (
            .O(N__24619),
            .I(N__24603));
    Odrv4 I__5841 (
            .O(N__24616),
            .I(\Lab_UT.sec1_0 ));
    Odrv4 I__5840 (
            .O(N__24613),
            .I(\Lab_UT.sec1_0 ));
    LocalMux I__5839 (
            .O(N__24610),
            .I(\Lab_UT.sec1_0 ));
    LocalMux I__5838 (
            .O(N__24603),
            .I(\Lab_UT.sec1_0 ));
    InMux I__5837 (
            .O(N__24594),
            .I(N__24591));
    LocalMux I__5836 (
            .O(N__24591),
            .I(\uu2.bitmapZ0Z_84 ));
    InMux I__5835 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__5834 (
            .O(N__24585),
            .I(N__24579));
    InMux I__5833 (
            .O(N__24584),
            .I(N__24571));
    InMux I__5832 (
            .O(N__24583),
            .I(N__24571));
    InMux I__5831 (
            .O(N__24582),
            .I(N__24571));
    Span4Mux_s3_v I__5830 (
            .O(N__24579),
            .I(N__24568));
    InMux I__5829 (
            .O(N__24578),
            .I(N__24565));
    LocalMux I__5828 (
            .O(N__24571),
            .I(N__24562));
    Odrv4 I__5827 (
            .O(N__24568),
            .I(\Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0 ));
    LocalMux I__5826 (
            .O(N__24565),
            .I(\Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0 ));
    Odrv4 I__5825 (
            .O(N__24562),
            .I(\Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0 ));
    CascadeMux I__5824 (
            .O(N__24555),
            .I(N__24548));
    CascadeMux I__5823 (
            .O(N__24554),
            .I(N__24540));
    CascadeMux I__5822 (
            .O(N__24553),
            .I(N__24537));
    InMux I__5821 (
            .O(N__24552),
            .I(N__24528));
    InMux I__5820 (
            .O(N__24551),
            .I(N__24528));
    InMux I__5819 (
            .O(N__24548),
            .I(N__24525));
    CascadeMux I__5818 (
            .O(N__24547),
            .I(N__24518));
    InMux I__5817 (
            .O(N__24546),
            .I(N__24515));
    InMux I__5816 (
            .O(N__24545),
            .I(N__24512));
    InMux I__5815 (
            .O(N__24544),
            .I(N__24509));
    InMux I__5814 (
            .O(N__24543),
            .I(N__24504));
    InMux I__5813 (
            .O(N__24540),
            .I(N__24504));
    InMux I__5812 (
            .O(N__24537),
            .I(N__24501));
    InMux I__5811 (
            .O(N__24536),
            .I(N__24498));
    InMux I__5810 (
            .O(N__24535),
            .I(N__24495));
    InMux I__5809 (
            .O(N__24534),
            .I(N__24492));
    CascadeMux I__5808 (
            .O(N__24533),
            .I(N__24486));
    LocalMux I__5807 (
            .O(N__24528),
            .I(N__24481));
    LocalMux I__5806 (
            .O(N__24525),
            .I(N__24478));
    InMux I__5805 (
            .O(N__24524),
            .I(N__24469));
    InMux I__5804 (
            .O(N__24523),
            .I(N__24469));
    InMux I__5803 (
            .O(N__24522),
            .I(N__24469));
    InMux I__5802 (
            .O(N__24521),
            .I(N__24469));
    InMux I__5801 (
            .O(N__24518),
            .I(N__24466));
    LocalMux I__5800 (
            .O(N__24515),
            .I(N__24463));
    LocalMux I__5799 (
            .O(N__24512),
            .I(N__24460));
    LocalMux I__5798 (
            .O(N__24509),
            .I(N__24451));
    LocalMux I__5797 (
            .O(N__24504),
            .I(N__24451));
    LocalMux I__5796 (
            .O(N__24501),
            .I(N__24451));
    LocalMux I__5795 (
            .O(N__24498),
            .I(N__24446));
    LocalMux I__5794 (
            .O(N__24495),
            .I(N__24446));
    LocalMux I__5793 (
            .O(N__24492),
            .I(N__24443));
    InMux I__5792 (
            .O(N__24491),
            .I(N__24438));
    InMux I__5791 (
            .O(N__24490),
            .I(N__24438));
    InMux I__5790 (
            .O(N__24489),
            .I(N__24433));
    InMux I__5789 (
            .O(N__24486),
            .I(N__24433));
    InMux I__5788 (
            .O(N__24485),
            .I(N__24430));
    InMux I__5787 (
            .O(N__24484),
            .I(N__24427));
    Span4Mux_s2_v I__5786 (
            .O(N__24481),
            .I(N__24420));
    Span4Mux_h I__5785 (
            .O(N__24478),
            .I(N__24420));
    LocalMux I__5784 (
            .O(N__24469),
            .I(N__24420));
    LocalMux I__5783 (
            .O(N__24466),
            .I(N__24417));
    Span4Mux_s2_v I__5782 (
            .O(N__24463),
            .I(N__24414));
    Span4Mux_h I__5781 (
            .O(N__24460),
            .I(N__24411));
    InMux I__5780 (
            .O(N__24459),
            .I(N__24406));
    InMux I__5779 (
            .O(N__24458),
            .I(N__24406));
    Span4Mux_h I__5778 (
            .O(N__24451),
            .I(N__24401));
    Span4Mux_h I__5777 (
            .O(N__24446),
            .I(N__24401));
    Span4Mux_s3_v I__5776 (
            .O(N__24443),
            .I(N__24394));
    LocalMux I__5775 (
            .O(N__24438),
            .I(N__24394));
    LocalMux I__5774 (
            .O(N__24433),
            .I(N__24394));
    LocalMux I__5773 (
            .O(N__24430),
            .I(N__24383));
    LocalMux I__5772 (
            .O(N__24427),
            .I(N__24383));
    Span4Mux_v I__5771 (
            .O(N__24420),
            .I(N__24383));
    Span4Mux_v I__5770 (
            .O(N__24417),
            .I(N__24383));
    Span4Mux_v I__5769 (
            .O(N__24414),
            .I(N__24383));
    Odrv4 I__5768 (
            .O(N__24411),
            .I(\Lab_UT.state_3 ));
    LocalMux I__5767 (
            .O(N__24406),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5766 (
            .O(N__24401),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5765 (
            .O(N__24394),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5764 (
            .O(N__24383),
            .I(\Lab_UT.state_3 ));
    InMux I__5763 (
            .O(N__24372),
            .I(N__24369));
    LocalMux I__5762 (
            .O(N__24369),
            .I(N__24365));
    InMux I__5761 (
            .O(N__24368),
            .I(N__24362));
    Span4Mux_v I__5760 (
            .O(N__24365),
            .I(N__24357));
    LocalMux I__5759 (
            .O(N__24362),
            .I(N__24357));
    Span4Mux_h I__5758 (
            .O(N__24357),
            .I(N__24354));
    Odrv4 I__5757 (
            .O(N__24354),
            .I(\Lab_UT.dictrl.N_40_1 ));
    InMux I__5756 (
            .O(N__24351),
            .I(N__24348));
    LocalMux I__5755 (
            .O(N__24348),
            .I(\Lab_UT.dictrl.g1 ));
    InMux I__5754 (
            .O(N__24345),
            .I(N__24342));
    LocalMux I__5753 (
            .O(N__24342),
            .I(N__24338));
    InMux I__5752 (
            .O(N__24341),
            .I(N__24335));
    Span4Mux_h I__5751 (
            .O(N__24338),
            .I(N__24332));
    LocalMux I__5750 (
            .O(N__24335),
            .I(N__24329));
    Odrv4 I__5749 (
            .O(N__24332),
            .I(\Lab_UT.dictrl.N_97_mux_4 ));
    Odrv4 I__5748 (
            .O(N__24329),
            .I(\Lab_UT.dictrl.N_97_mux_4 ));
    InMux I__5747 (
            .O(N__24324),
            .I(N__24313));
    CascadeMux I__5746 (
            .O(N__24323),
            .I(N__24310));
    InMux I__5745 (
            .O(N__24322),
            .I(N__24300));
    InMux I__5744 (
            .O(N__24321),
            .I(N__24295));
    InMux I__5743 (
            .O(N__24320),
            .I(N__24295));
    InMux I__5742 (
            .O(N__24319),
            .I(N__24283));
    InMux I__5741 (
            .O(N__24318),
            .I(N__24283));
    InMux I__5740 (
            .O(N__24317),
            .I(N__24283));
    InMux I__5739 (
            .O(N__24316),
            .I(N__24283));
    LocalMux I__5738 (
            .O(N__24313),
            .I(N__24280));
    InMux I__5737 (
            .O(N__24310),
            .I(N__24272));
    InMux I__5736 (
            .O(N__24309),
            .I(N__24272));
    InMux I__5735 (
            .O(N__24308),
            .I(N__24268));
    InMux I__5734 (
            .O(N__24307),
            .I(N__24265));
    InMux I__5733 (
            .O(N__24306),
            .I(N__24262));
    InMux I__5732 (
            .O(N__24305),
            .I(N__24259));
    InMux I__5731 (
            .O(N__24304),
            .I(N__24254));
    InMux I__5730 (
            .O(N__24303),
            .I(N__24254));
    LocalMux I__5729 (
            .O(N__24300),
            .I(N__24249));
    LocalMux I__5728 (
            .O(N__24295),
            .I(N__24249));
    InMux I__5727 (
            .O(N__24294),
            .I(N__24246));
    InMux I__5726 (
            .O(N__24293),
            .I(N__24243));
    InMux I__5725 (
            .O(N__24292),
            .I(N__24240));
    LocalMux I__5724 (
            .O(N__24283),
            .I(N__24237));
    Span4Mux_s2_v I__5723 (
            .O(N__24280),
            .I(N__24234));
    InMux I__5722 (
            .O(N__24279),
            .I(N__24229));
    InMux I__5721 (
            .O(N__24278),
            .I(N__24229));
    InMux I__5720 (
            .O(N__24277),
            .I(N__24226));
    LocalMux I__5719 (
            .O(N__24272),
            .I(N__24223));
    InMux I__5718 (
            .O(N__24271),
            .I(N__24220));
    LocalMux I__5717 (
            .O(N__24268),
            .I(N__24217));
    LocalMux I__5716 (
            .O(N__24265),
            .I(N__24210));
    LocalMux I__5715 (
            .O(N__24262),
            .I(N__24210));
    LocalMux I__5714 (
            .O(N__24259),
            .I(N__24210));
    LocalMux I__5713 (
            .O(N__24254),
            .I(N__24201));
    Span4Mux_h I__5712 (
            .O(N__24249),
            .I(N__24201));
    LocalMux I__5711 (
            .O(N__24246),
            .I(N__24201));
    LocalMux I__5710 (
            .O(N__24243),
            .I(N__24201));
    LocalMux I__5709 (
            .O(N__24240),
            .I(N__24196));
    Span4Mux_s3_h I__5708 (
            .O(N__24237),
            .I(N__24196));
    Span4Mux_v I__5707 (
            .O(N__24234),
            .I(N__24191));
    LocalMux I__5706 (
            .O(N__24229),
            .I(N__24191));
    LocalMux I__5705 (
            .O(N__24226),
            .I(N__24186));
    Span4Mux_s3_h I__5704 (
            .O(N__24223),
            .I(N__24186));
    LocalMux I__5703 (
            .O(N__24220),
            .I(N__24183));
    Span4Mux_v I__5702 (
            .O(N__24217),
            .I(N__24178));
    Span4Mux_v I__5701 (
            .O(N__24210),
            .I(N__24178));
    Span4Mux_v I__5700 (
            .O(N__24201),
            .I(N__24173));
    Span4Mux_h I__5699 (
            .O(N__24196),
            .I(N__24173));
    Odrv4 I__5698 (
            .O(N__24191),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5697 (
            .O(N__24186),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv12 I__5696 (
            .O(N__24183),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5695 (
            .O(N__24178),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5694 (
            .O(N__24173),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    CascadeMux I__5693 (
            .O(N__24162),
            .I(N__24159));
    InMux I__5692 (
            .O(N__24159),
            .I(N__24156));
    LocalMux I__5691 (
            .O(N__24156),
            .I(N__24153));
    Span4Mux_v I__5690 (
            .O(N__24153),
            .I(N__24150));
    Odrv4 I__5689 (
            .O(N__24150),
            .I(\Lab_UT.dictrl.g1_1_1 ));
    InMux I__5688 (
            .O(N__24147),
            .I(N__24141));
    InMux I__5687 (
            .O(N__24146),
            .I(N__24136));
    InMux I__5686 (
            .O(N__24145),
            .I(N__24136));
    InMux I__5685 (
            .O(N__24144),
            .I(N__24133));
    LocalMux I__5684 (
            .O(N__24141),
            .I(N__24130));
    LocalMux I__5683 (
            .O(N__24136),
            .I(N__24127));
    LocalMux I__5682 (
            .O(N__24133),
            .I(N__24122));
    Span4Mux_v I__5681 (
            .O(N__24130),
            .I(N__24122));
    Span4Mux_s3_h I__5680 (
            .O(N__24127),
            .I(N__24119));
    Span4Mux_h I__5679 (
            .O(N__24122),
            .I(N__24116));
    Span4Mux_h I__5678 (
            .O(N__24119),
            .I(N__24113));
    Odrv4 I__5677 (
            .O(N__24116),
            .I(\Lab_UT.dictrl.m34_4 ));
    Odrv4 I__5676 (
            .O(N__24113),
            .I(\Lab_UT.dictrl.m34_4 ));
    InMux I__5675 (
            .O(N__24108),
            .I(N__24105));
    LocalMux I__5674 (
            .O(N__24105),
            .I(N__24102));
    Odrv4 I__5673 (
            .O(N__24102),
            .I(\Lab_UT.dictrl.N_1106_0 ));
    InMux I__5672 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__5671 (
            .O(N__24096),
            .I(N__24093));
    Span4Mux_s2_v I__5670 (
            .O(N__24093),
            .I(N__24090));
    Odrv4 I__5669 (
            .O(N__24090),
            .I(\Lab_UT.dictrl.N_1462_1 ));
    InMux I__5668 (
            .O(N__24087),
            .I(N__24084));
    LocalMux I__5667 (
            .O(N__24084),
            .I(N__24081));
    Span4Mux_s3_h I__5666 (
            .O(N__24081),
            .I(N__24078));
    Odrv4 I__5665 (
            .O(N__24078),
            .I(\Lab_UT.dictrl.N_1102_1 ));
    CascadeMux I__5664 (
            .O(N__24075),
            .I(N__24072));
    InMux I__5663 (
            .O(N__24072),
            .I(N__24069));
    LocalMux I__5662 (
            .O(N__24069),
            .I(N__24066));
    Odrv4 I__5661 (
            .O(N__24066),
            .I(\Lab_UT.dictrl.g2_1_1 ));
    InMux I__5660 (
            .O(N__24063),
            .I(N__24059));
    InMux I__5659 (
            .O(N__24062),
            .I(N__24045));
    LocalMux I__5658 (
            .O(N__24059),
            .I(N__24042));
    CascadeMux I__5657 (
            .O(N__24058),
            .I(N__24027));
    CascadeMux I__5656 (
            .O(N__24057),
            .I(N__24024));
    InMux I__5655 (
            .O(N__24056),
            .I(N__24021));
    InMux I__5654 (
            .O(N__24055),
            .I(N__24018));
    CascadeMux I__5653 (
            .O(N__24054),
            .I(N__24008));
    CascadeMux I__5652 (
            .O(N__24053),
            .I(N__24005));
    CascadeMux I__5651 (
            .O(N__24052),
            .I(N__23994));
    CascadeMux I__5650 (
            .O(N__24051),
            .I(N__23991));
    CascadeMux I__5649 (
            .O(N__24050),
            .I(N__23988));
    CascadeMux I__5648 (
            .O(N__24049),
            .I(N__23985));
    InMux I__5647 (
            .O(N__24048),
            .I(N__23978));
    LocalMux I__5646 (
            .O(N__24045),
            .I(N__23975));
    Span4Mux_h I__5645 (
            .O(N__24042),
            .I(N__23972));
    InMux I__5644 (
            .O(N__24041),
            .I(N__23969));
    InMux I__5643 (
            .O(N__24040),
            .I(N__23959));
    InMux I__5642 (
            .O(N__24039),
            .I(N__23955));
    InMux I__5641 (
            .O(N__24038),
            .I(N__23940));
    InMux I__5640 (
            .O(N__24037),
            .I(N__23940));
    InMux I__5639 (
            .O(N__24036),
            .I(N__23940));
    InMux I__5638 (
            .O(N__24035),
            .I(N__23940));
    InMux I__5637 (
            .O(N__24034),
            .I(N__23940));
    InMux I__5636 (
            .O(N__24033),
            .I(N__23940));
    InMux I__5635 (
            .O(N__24032),
            .I(N__23940));
    InMux I__5634 (
            .O(N__24031),
            .I(N__23935));
    InMux I__5633 (
            .O(N__24030),
            .I(N__23935));
    InMux I__5632 (
            .O(N__24027),
            .I(N__23930));
    InMux I__5631 (
            .O(N__24024),
            .I(N__23930));
    LocalMux I__5630 (
            .O(N__24021),
            .I(N__23925));
    LocalMux I__5629 (
            .O(N__24018),
            .I(N__23925));
    InMux I__5628 (
            .O(N__24017),
            .I(N__23922));
    InMux I__5627 (
            .O(N__24016),
            .I(N__23919));
    InMux I__5626 (
            .O(N__24015),
            .I(N__23912));
    InMux I__5625 (
            .O(N__24014),
            .I(N__23912));
    InMux I__5624 (
            .O(N__24013),
            .I(N__23912));
    CascadeMux I__5623 (
            .O(N__24012),
            .I(N__23906));
    InMux I__5622 (
            .O(N__24011),
            .I(N__23902));
    InMux I__5621 (
            .O(N__24008),
            .I(N__23893));
    InMux I__5620 (
            .O(N__24005),
            .I(N__23893));
    InMux I__5619 (
            .O(N__24004),
            .I(N__23893));
    InMux I__5618 (
            .O(N__24003),
            .I(N__23893));
    InMux I__5617 (
            .O(N__24002),
            .I(N__23890));
    InMux I__5616 (
            .O(N__24001),
            .I(N__23883));
    InMux I__5615 (
            .O(N__24000),
            .I(N__23883));
    InMux I__5614 (
            .O(N__23999),
            .I(N__23883));
    InMux I__5613 (
            .O(N__23998),
            .I(N__23876));
    InMux I__5612 (
            .O(N__23997),
            .I(N__23876));
    InMux I__5611 (
            .O(N__23994),
            .I(N__23876));
    InMux I__5610 (
            .O(N__23991),
            .I(N__23869));
    InMux I__5609 (
            .O(N__23988),
            .I(N__23869));
    InMux I__5608 (
            .O(N__23985),
            .I(N__23869));
    InMux I__5607 (
            .O(N__23984),
            .I(N__23866));
    InMux I__5606 (
            .O(N__23983),
            .I(N__23859));
    InMux I__5605 (
            .O(N__23982),
            .I(N__23859));
    InMux I__5604 (
            .O(N__23981),
            .I(N__23859));
    LocalMux I__5603 (
            .O(N__23978),
            .I(N__23854));
    Span4Mux_v I__5602 (
            .O(N__23975),
            .I(N__23854));
    IoSpan4Mux I__5601 (
            .O(N__23972),
            .I(N__23849));
    LocalMux I__5600 (
            .O(N__23969),
            .I(N__23849));
    InMux I__5599 (
            .O(N__23968),
            .I(N__23840));
    InMux I__5598 (
            .O(N__23967),
            .I(N__23840));
    InMux I__5597 (
            .O(N__23966),
            .I(N__23840));
    InMux I__5596 (
            .O(N__23965),
            .I(N__23840));
    InMux I__5595 (
            .O(N__23964),
            .I(N__23833));
    InMux I__5594 (
            .O(N__23963),
            .I(N__23833));
    InMux I__5593 (
            .O(N__23962),
            .I(N__23833));
    LocalMux I__5592 (
            .O(N__23959),
            .I(N__23830));
    InMux I__5591 (
            .O(N__23958),
            .I(N__23824));
    LocalMux I__5590 (
            .O(N__23955),
            .I(N__23821));
    LocalMux I__5589 (
            .O(N__23940),
            .I(N__23818));
    LocalMux I__5588 (
            .O(N__23935),
            .I(N__23805));
    LocalMux I__5587 (
            .O(N__23930),
            .I(N__23805));
    Span4Mux_h I__5586 (
            .O(N__23925),
            .I(N__23805));
    LocalMux I__5585 (
            .O(N__23922),
            .I(N__23805));
    LocalMux I__5584 (
            .O(N__23919),
            .I(N__23805));
    LocalMux I__5583 (
            .O(N__23912),
            .I(N__23805));
    InMux I__5582 (
            .O(N__23911),
            .I(N__23802));
    InMux I__5581 (
            .O(N__23910),
            .I(N__23793));
    InMux I__5580 (
            .O(N__23909),
            .I(N__23793));
    InMux I__5579 (
            .O(N__23906),
            .I(N__23793));
    InMux I__5578 (
            .O(N__23905),
            .I(N__23793));
    LocalMux I__5577 (
            .O(N__23902),
            .I(N__23790));
    LocalMux I__5576 (
            .O(N__23893),
            .I(N__23783));
    LocalMux I__5575 (
            .O(N__23890),
            .I(N__23783));
    LocalMux I__5574 (
            .O(N__23883),
            .I(N__23783));
    LocalMux I__5573 (
            .O(N__23876),
            .I(N__23776));
    LocalMux I__5572 (
            .O(N__23869),
            .I(N__23776));
    LocalMux I__5571 (
            .O(N__23866),
            .I(N__23776));
    LocalMux I__5570 (
            .O(N__23859),
            .I(N__23769));
    Span4Mux_h I__5569 (
            .O(N__23854),
            .I(N__23769));
    Span4Mux_s2_v I__5568 (
            .O(N__23849),
            .I(N__23769));
    LocalMux I__5567 (
            .O(N__23840),
            .I(N__23762));
    LocalMux I__5566 (
            .O(N__23833),
            .I(N__23762));
    Span4Mux_s2_v I__5565 (
            .O(N__23830),
            .I(N__23762));
    InMux I__5564 (
            .O(N__23829),
            .I(N__23759));
    InMux I__5563 (
            .O(N__23828),
            .I(N__23754));
    InMux I__5562 (
            .O(N__23827),
            .I(N__23754));
    LocalMux I__5561 (
            .O(N__23824),
            .I(N__23749));
    Span4Mux_h I__5560 (
            .O(N__23821),
            .I(N__23749));
    Span4Mux_v I__5559 (
            .O(N__23818),
            .I(N__23744));
    Span4Mux_v I__5558 (
            .O(N__23805),
            .I(N__23744));
    LocalMux I__5557 (
            .O(N__23802),
            .I(N__23735));
    LocalMux I__5556 (
            .O(N__23793),
            .I(N__23735));
    Span12Mux_s4_h I__5555 (
            .O(N__23790),
            .I(N__23735));
    Span12Mux_s5_v I__5554 (
            .O(N__23783),
            .I(N__23735));
    Span4Mux_h I__5553 (
            .O(N__23776),
            .I(N__23728));
    Span4Mux_h I__5552 (
            .O(N__23769),
            .I(N__23728));
    Span4Mux_h I__5551 (
            .O(N__23762),
            .I(N__23728));
    LocalMux I__5550 (
            .O(N__23759),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__5549 (
            .O(N__23754),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5548 (
            .O(N__23749),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5547 (
            .O(N__23744),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv12 I__5546 (
            .O(N__23735),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5545 (
            .O(N__23728),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    InMux I__5544 (
            .O(N__23715),
            .I(N__23712));
    LocalMux I__5543 (
            .O(N__23712),
            .I(N__23709));
    Odrv12 I__5542 (
            .O(N__23709),
            .I(\Lab_UT.dictrl.N_1460_1 ));
    CascadeMux I__5541 (
            .O(N__23706),
            .I(N__23701));
    CascadeMux I__5540 (
            .O(N__23705),
            .I(N__23698));
    InMux I__5539 (
            .O(N__23704),
            .I(N__23694));
    InMux I__5538 (
            .O(N__23701),
            .I(N__23684));
    InMux I__5537 (
            .O(N__23698),
            .I(N__23684));
    InMux I__5536 (
            .O(N__23697),
            .I(N__23684));
    LocalMux I__5535 (
            .O(N__23694),
            .I(N__23681));
    CascadeMux I__5534 (
            .O(N__23693),
            .I(N__23677));
    CascadeMux I__5533 (
            .O(N__23692),
            .I(N__23673));
    CascadeMux I__5532 (
            .O(N__23691),
            .I(N__23670));
    LocalMux I__5531 (
            .O(N__23684),
            .I(N__23663));
    Span4Mux_s2_h I__5530 (
            .O(N__23681),
            .I(N__23663));
    InMux I__5529 (
            .O(N__23680),
            .I(N__23655));
    InMux I__5528 (
            .O(N__23677),
            .I(N__23655));
    InMux I__5527 (
            .O(N__23676),
            .I(N__23655));
    InMux I__5526 (
            .O(N__23673),
            .I(N__23646));
    InMux I__5525 (
            .O(N__23670),
            .I(N__23646));
    InMux I__5524 (
            .O(N__23669),
            .I(N__23646));
    InMux I__5523 (
            .O(N__23668),
            .I(N__23646));
    Span4Mux_h I__5522 (
            .O(N__23663),
            .I(N__23643));
    InMux I__5521 (
            .O(N__23662),
            .I(N__23638));
    LocalMux I__5520 (
            .O(N__23655),
            .I(N__23635));
    LocalMux I__5519 (
            .O(N__23646),
            .I(N__23630));
    IoSpan4Mux I__5518 (
            .O(N__23643),
            .I(N__23630));
    InMux I__5517 (
            .O(N__23642),
            .I(N__23625));
    InMux I__5516 (
            .O(N__23641),
            .I(N__23625));
    LocalMux I__5515 (
            .O(N__23638),
            .I(L3_tx_data_rdy));
    Odrv4 I__5514 (
            .O(N__23635),
            .I(L3_tx_data_rdy));
    Odrv4 I__5513 (
            .O(N__23630),
            .I(L3_tx_data_rdy));
    LocalMux I__5512 (
            .O(N__23625),
            .I(L3_tx_data_rdy));
    InMux I__5511 (
            .O(N__23616),
            .I(N__23613));
    LocalMux I__5510 (
            .O(N__23613),
            .I(N__23610));
    Span4Mux_s1_h I__5509 (
            .O(N__23610),
            .I(N__23600));
    InMux I__5508 (
            .O(N__23609),
            .I(N__23593));
    InMux I__5507 (
            .O(N__23608),
            .I(N__23593));
    InMux I__5506 (
            .O(N__23607),
            .I(N__23593));
    InMux I__5505 (
            .O(N__23606),
            .I(N__23581));
    InMux I__5504 (
            .O(N__23605),
            .I(N__23581));
    InMux I__5503 (
            .O(N__23604),
            .I(N__23581));
    InMux I__5502 (
            .O(N__23603),
            .I(N__23581));
    Span4Mux_h I__5501 (
            .O(N__23600),
            .I(N__23575));
    LocalMux I__5500 (
            .O(N__23593),
            .I(N__23572));
    InMux I__5499 (
            .O(N__23592),
            .I(N__23565));
    InMux I__5498 (
            .O(N__23591),
            .I(N__23565));
    InMux I__5497 (
            .O(N__23590),
            .I(N__23565));
    LocalMux I__5496 (
            .O(N__23581),
            .I(N__23562));
    InMux I__5495 (
            .O(N__23580),
            .I(N__23555));
    InMux I__5494 (
            .O(N__23579),
            .I(N__23555));
    InMux I__5493 (
            .O(N__23578),
            .I(N__23555));
    Odrv4 I__5492 (
            .O(N__23575),
            .I(\uu2.un1_w_user_cr_0 ));
    Odrv4 I__5491 (
            .O(N__23572),
            .I(\uu2.un1_w_user_cr_0 ));
    LocalMux I__5490 (
            .O(N__23565),
            .I(\uu2.un1_w_user_cr_0 ));
    Odrv4 I__5489 (
            .O(N__23562),
            .I(\uu2.un1_w_user_cr_0 ));
    LocalMux I__5488 (
            .O(N__23555),
            .I(\uu2.un1_w_user_cr_0 ));
    CascadeMux I__5487 (
            .O(N__23544),
            .I(N__23540));
    InMux I__5486 (
            .O(N__23543),
            .I(N__23537));
    InMux I__5485 (
            .O(N__23540),
            .I(N__23534));
    LocalMux I__5484 (
            .O(N__23537),
            .I(N__23530));
    LocalMux I__5483 (
            .O(N__23534),
            .I(N__23527));
    InMux I__5482 (
            .O(N__23533),
            .I(N__23524));
    Span4Mux_s1_v I__5481 (
            .O(N__23530),
            .I(N__23521));
    Span12Mux_s1_h I__5480 (
            .O(N__23527),
            .I(N__23518));
    LocalMux I__5479 (
            .O(N__23524),
            .I(\uu2.w_addr_userZ0Z_8 ));
    Odrv4 I__5478 (
            .O(N__23521),
            .I(\uu2.w_addr_userZ0Z_8 ));
    Odrv12 I__5477 (
            .O(N__23518),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CascadeMux I__5476 (
            .O(N__23511),
            .I(N__23508));
    InMux I__5475 (
            .O(N__23508),
            .I(N__23505));
    LocalMux I__5474 (
            .O(N__23505),
            .I(N__23502));
    Span4Mux_s1_v I__5473 (
            .O(N__23502),
            .I(N__23499));
    Span4Mux_h I__5472 (
            .O(N__23499),
            .I(N__23496));
    Span4Mux_h I__5471 (
            .O(N__23496),
            .I(N__23493));
    Odrv4 I__5470 (
            .O(N__23493),
            .I(\uu2.mem0.w_addr_8 ));
    InMux I__5469 (
            .O(N__23490),
            .I(N__23482));
    InMux I__5468 (
            .O(N__23489),
            .I(N__23475));
    InMux I__5467 (
            .O(N__23488),
            .I(N__23475));
    InMux I__5466 (
            .O(N__23487),
            .I(N__23475));
    InMux I__5465 (
            .O(N__23486),
            .I(N__23468));
    CascadeMux I__5464 (
            .O(N__23485),
            .I(N__23465));
    LocalMux I__5463 (
            .O(N__23482),
            .I(N__23457));
    LocalMux I__5462 (
            .O(N__23475),
            .I(N__23457));
    InMux I__5461 (
            .O(N__23474),
            .I(N__23450));
    InMux I__5460 (
            .O(N__23473),
            .I(N__23450));
    InMux I__5459 (
            .O(N__23472),
            .I(N__23450));
    InMux I__5458 (
            .O(N__23471),
            .I(N__23447));
    LocalMux I__5457 (
            .O(N__23468),
            .I(N__23444));
    InMux I__5456 (
            .O(N__23465),
            .I(N__23435));
    InMux I__5455 (
            .O(N__23464),
            .I(N__23435));
    InMux I__5454 (
            .O(N__23463),
            .I(N__23435));
    InMux I__5453 (
            .O(N__23462),
            .I(N__23435));
    Span4Mux_h I__5452 (
            .O(N__23457),
            .I(N__23432));
    LocalMux I__5451 (
            .O(N__23450),
            .I(N__23429));
    LocalMux I__5450 (
            .O(N__23447),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv12 I__5449 (
            .O(N__23444),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__5448 (
            .O(N__23435),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__5447 (
            .O(N__23432),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__5446 (
            .O(N__23429),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    InMux I__5445 (
            .O(N__23418),
            .I(N__23414));
    InMux I__5444 (
            .O(N__23417),
            .I(N__23411));
    LocalMux I__5443 (
            .O(N__23414),
            .I(N__23408));
    LocalMux I__5442 (
            .O(N__23411),
            .I(N__23405));
    Span4Mux_s1_v I__5441 (
            .O(N__23408),
            .I(N__23397));
    Span4Mux_s2_h I__5440 (
            .O(N__23405),
            .I(N__23397));
    InMux I__5439 (
            .O(N__23404),
            .I(N__23390));
    InMux I__5438 (
            .O(N__23403),
            .I(N__23390));
    InMux I__5437 (
            .O(N__23402),
            .I(N__23390));
    Odrv4 I__5436 (
            .O(N__23397),
            .I(\uu2.N_75_mux ));
    LocalMux I__5435 (
            .O(N__23390),
            .I(\uu2.N_75_mux ));
    CascadeMux I__5434 (
            .O(N__23385),
            .I(N__23382));
    InMux I__5433 (
            .O(N__23382),
            .I(N__23377));
    InMux I__5432 (
            .O(N__23381),
            .I(N__23374));
    CascadeMux I__5431 (
            .O(N__23380),
            .I(N__23369));
    LocalMux I__5430 (
            .O(N__23377),
            .I(N__23366));
    LocalMux I__5429 (
            .O(N__23374),
            .I(N__23363));
    CascadeMux I__5428 (
            .O(N__23373),
            .I(N__23359));
    InMux I__5427 (
            .O(N__23372),
            .I(N__23354));
    InMux I__5426 (
            .O(N__23369),
            .I(N__23354));
    Span4Mux_h I__5425 (
            .O(N__23366),
            .I(N__23349));
    Span4Mux_h I__5424 (
            .O(N__23363),
            .I(N__23349));
    InMux I__5423 (
            .O(N__23362),
            .I(N__23344));
    InMux I__5422 (
            .O(N__23359),
            .I(N__23344));
    LocalMux I__5421 (
            .O(N__23354),
            .I(N__23335));
    IoSpan4Mux I__5420 (
            .O(N__23349),
            .I(N__23335));
    LocalMux I__5419 (
            .O(N__23344),
            .I(N__23335));
    CascadeMux I__5418 (
            .O(N__23343),
            .I(N__23331));
    CascadeMux I__5417 (
            .O(N__23342),
            .I(N__23324));
    Sp12to4 I__5416 (
            .O(N__23335),
            .I(N__23321));
    InMux I__5415 (
            .O(N__23334),
            .I(N__23310));
    InMux I__5414 (
            .O(N__23331),
            .I(N__23310));
    InMux I__5413 (
            .O(N__23330),
            .I(N__23310));
    InMux I__5412 (
            .O(N__23329),
            .I(N__23310));
    InMux I__5411 (
            .O(N__23328),
            .I(N__23310));
    InMux I__5410 (
            .O(N__23327),
            .I(N__23305));
    InMux I__5409 (
            .O(N__23324),
            .I(N__23305));
    Span12Mux_s1_v I__5408 (
            .O(N__23321),
            .I(N__23300));
    LocalMux I__5407 (
            .O(N__23310),
            .I(N__23300));
    LocalMux I__5406 (
            .O(N__23305),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv12 I__5405 (
            .O(N__23300),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__5404 (
            .O(N__23295),
            .I(N__23292));
    LocalMux I__5403 (
            .O(N__23292),
            .I(N__23286));
    InMux I__5402 (
            .O(N__23291),
            .I(N__23279));
    InMux I__5401 (
            .O(N__23290),
            .I(N__23279));
    InMux I__5400 (
            .O(N__23289),
            .I(N__23279));
    Span4Mux_s2_h I__5399 (
            .O(N__23286),
            .I(N__23274));
    LocalMux I__5398 (
            .O(N__23279),
            .I(N__23271));
    InMux I__5397 (
            .O(N__23278),
            .I(N__23266));
    InMux I__5396 (
            .O(N__23277),
            .I(N__23266));
    Odrv4 I__5395 (
            .O(N__23274),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__5394 (
            .O(N__23271),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__5393 (
            .O(N__23266),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    CascadeMux I__5392 (
            .O(N__23259),
            .I(\uu2.N_14_i_cascade_ ));
    CascadeMux I__5391 (
            .O(N__23256),
            .I(N__23253));
    InMux I__5390 (
            .O(N__23253),
            .I(N__23238));
    InMux I__5389 (
            .O(N__23252),
            .I(N__23238));
    InMux I__5388 (
            .O(N__23251),
            .I(N__23238));
    InMux I__5387 (
            .O(N__23250),
            .I(N__23238));
    InMux I__5386 (
            .O(N__23249),
            .I(N__23238));
    LocalMux I__5385 (
            .O(N__23238),
            .I(N__23235));
    Span4Mux_v I__5384 (
            .O(N__23235),
            .I(N__23232));
    Odrv4 I__5383 (
            .O(N__23232),
            .I(\uu2.N_15_i ));
    InMux I__5382 (
            .O(N__23229),
            .I(N__23226));
    LocalMux I__5381 (
            .O(N__23226),
            .I(N__23223));
    Odrv4 I__5380 (
            .O(N__23223),
            .I(\Lab_UT.dictrl.state_ret_12and_0_ns_sn ));
    InMux I__5379 (
            .O(N__23220),
            .I(N__23217));
    LocalMux I__5378 (
            .O(N__23217),
            .I(N__23214));
    Odrv12 I__5377 (
            .O(N__23214),
            .I(\Lab_UT.dictrl.state_ret_12and_0_ns_rn_0 ));
    CascadeMux I__5376 (
            .O(N__23211),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ));
    InMux I__5375 (
            .O(N__23208),
            .I(N__23205));
    LocalMux I__5374 (
            .O(N__23205),
            .I(N__23199));
    InMux I__5373 (
            .O(N__23204),
            .I(N__23192));
    InMux I__5372 (
            .O(N__23203),
            .I(N__23192));
    InMux I__5371 (
            .O(N__23202),
            .I(N__23192));
    Span4Mux_s3_h I__5370 (
            .O(N__23199),
            .I(N__23188));
    LocalMux I__5369 (
            .O(N__23192),
            .I(N__23185));
    InMux I__5368 (
            .O(N__23191),
            .I(N__23182));
    Odrv4 I__5367 (
            .O(N__23188),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    Odrv12 I__5366 (
            .O(N__23185),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    LocalMux I__5365 (
            .O(N__23182),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    CascadeMux I__5364 (
            .O(N__23175),
            .I(\Lab_UT.dictrl.g2_0_cascade_ ));
    InMux I__5363 (
            .O(N__23172),
            .I(N__23169));
    LocalMux I__5362 (
            .O(N__23169),
            .I(\Lab_UT.dictrl.next_state_2_0_1 ));
    CascadeMux I__5361 (
            .O(N__23166),
            .I(N__23156));
    CascadeMux I__5360 (
            .O(N__23165),
            .I(N__23149));
    CascadeMux I__5359 (
            .O(N__23164),
            .I(N__23145));
    CascadeMux I__5358 (
            .O(N__23163),
            .I(N__23142));
    CascadeMux I__5357 (
            .O(N__23162),
            .I(N__23139));
    CascadeMux I__5356 (
            .O(N__23161),
            .I(N__23134));
    CascadeMux I__5355 (
            .O(N__23160),
            .I(N__23129));
    InMux I__5354 (
            .O(N__23159),
            .I(N__23124));
    InMux I__5353 (
            .O(N__23156),
            .I(N__23124));
    CascadeMux I__5352 (
            .O(N__23155),
            .I(N__23120));
    InMux I__5351 (
            .O(N__23154),
            .I(N__23104));
    InMux I__5350 (
            .O(N__23153),
            .I(N__23104));
    InMux I__5349 (
            .O(N__23152),
            .I(N__23104));
    InMux I__5348 (
            .O(N__23149),
            .I(N__23104));
    InMux I__5347 (
            .O(N__23148),
            .I(N__23104));
    InMux I__5346 (
            .O(N__23145),
            .I(N__23104));
    InMux I__5345 (
            .O(N__23142),
            .I(N__23104));
    InMux I__5344 (
            .O(N__23139),
            .I(N__23101));
    InMux I__5343 (
            .O(N__23138),
            .I(N__23098));
    InMux I__5342 (
            .O(N__23137),
            .I(N__23095));
    InMux I__5341 (
            .O(N__23134),
            .I(N__23090));
    InMux I__5340 (
            .O(N__23133),
            .I(N__23090));
    InMux I__5339 (
            .O(N__23132),
            .I(N__23085));
    InMux I__5338 (
            .O(N__23129),
            .I(N__23085));
    LocalMux I__5337 (
            .O(N__23124),
            .I(N__23079));
    InMux I__5336 (
            .O(N__23123),
            .I(N__23074));
    InMux I__5335 (
            .O(N__23120),
            .I(N__23074));
    InMux I__5334 (
            .O(N__23119),
            .I(N__23071));
    LocalMux I__5333 (
            .O(N__23104),
            .I(N__23066));
    LocalMux I__5332 (
            .O(N__23101),
            .I(N__23066));
    LocalMux I__5331 (
            .O(N__23098),
            .I(N__23063));
    LocalMux I__5330 (
            .O(N__23095),
            .I(N__23060));
    LocalMux I__5329 (
            .O(N__23090),
            .I(N__23055));
    LocalMux I__5328 (
            .O(N__23085),
            .I(N__23055));
    InMux I__5327 (
            .O(N__23084),
            .I(N__23052));
    InMux I__5326 (
            .O(N__23083),
            .I(N__23049));
    InMux I__5325 (
            .O(N__23082),
            .I(N__23046));
    Span4Mux_s2_v I__5324 (
            .O(N__23079),
            .I(N__23041));
    LocalMux I__5323 (
            .O(N__23074),
            .I(N__23041));
    LocalMux I__5322 (
            .O(N__23071),
            .I(N__23036));
    Span4Mux_h I__5321 (
            .O(N__23066),
            .I(N__23036));
    Span4Mux_v I__5320 (
            .O(N__23063),
            .I(N__23029));
    Span4Mux_v I__5319 (
            .O(N__23060),
            .I(N__23029));
    Span4Mux_v I__5318 (
            .O(N__23055),
            .I(N__23029));
    LocalMux I__5317 (
            .O(N__23052),
            .I(N__23026));
    LocalMux I__5316 (
            .O(N__23049),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5315 (
            .O(N__23046),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5314 (
            .O(N__23041),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5313 (
            .O(N__23036),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5312 (
            .O(N__23029),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv12 I__5311 (
            .O(N__23026),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    InMux I__5310 (
            .O(N__23013),
            .I(N__23010));
    LocalMux I__5309 (
            .O(N__23010),
            .I(N__23007));
    Odrv4 I__5308 (
            .O(N__23007),
            .I(\Lab_UT.dictrl.N_1460_0 ));
    CascadeMux I__5307 (
            .O(N__23004),
            .I(\Lab_UT.dictrl.g2_cascade_ ));
    InMux I__5306 (
            .O(N__23001),
            .I(N__22998));
    LocalMux I__5305 (
            .O(N__22998),
            .I(N__22995));
    Odrv4 I__5304 (
            .O(N__22995),
            .I(\Lab_UT.dictrl.next_state_0_1 ));
    InMux I__5303 (
            .O(N__22992),
            .I(N__22989));
    LocalMux I__5302 (
            .O(N__22989),
            .I(N__22986));
    Odrv12 I__5301 (
            .O(N__22986),
            .I(\Lab_UT.dictrl.N_40_3 ));
    CascadeMux I__5300 (
            .O(N__22983),
            .I(\Lab_UT.dictrl.N_1105_1_cascade_ ));
    InMux I__5299 (
            .O(N__22980),
            .I(N__22974));
    InMux I__5298 (
            .O(N__22979),
            .I(N__22969));
    InMux I__5297 (
            .O(N__22978),
            .I(N__22963));
    InMux I__5296 (
            .O(N__22977),
            .I(N__22960));
    LocalMux I__5295 (
            .O(N__22974),
            .I(N__22957));
    InMux I__5294 (
            .O(N__22973),
            .I(N__22952));
    InMux I__5293 (
            .O(N__22972),
            .I(N__22952));
    LocalMux I__5292 (
            .O(N__22969),
            .I(N__22949));
    InMux I__5291 (
            .O(N__22968),
            .I(N__22940));
    InMux I__5290 (
            .O(N__22967),
            .I(N__22937));
    InMux I__5289 (
            .O(N__22966),
            .I(N__22934));
    LocalMux I__5288 (
            .O(N__22963),
            .I(N__22931));
    LocalMux I__5287 (
            .O(N__22960),
            .I(N__22928));
    Span4Mux_v I__5286 (
            .O(N__22957),
            .I(N__22921));
    LocalMux I__5285 (
            .O(N__22952),
            .I(N__22921));
    Span4Mux_v I__5284 (
            .O(N__22949),
            .I(N__22921));
    InMux I__5283 (
            .O(N__22948),
            .I(N__22914));
    InMux I__5282 (
            .O(N__22947),
            .I(N__22914));
    InMux I__5281 (
            .O(N__22946),
            .I(N__22914));
    InMux I__5280 (
            .O(N__22945),
            .I(N__22907));
    InMux I__5279 (
            .O(N__22944),
            .I(N__22907));
    InMux I__5278 (
            .O(N__22943),
            .I(N__22907));
    LocalMux I__5277 (
            .O(N__22940),
            .I(N__22904));
    LocalMux I__5276 (
            .O(N__22937),
            .I(N__22899));
    LocalMux I__5275 (
            .O(N__22934),
            .I(N__22899));
    Span4Mux_s3_v I__5274 (
            .O(N__22931),
            .I(N__22894));
    Span4Mux_h I__5273 (
            .O(N__22928),
            .I(N__22894));
    Span4Mux_h I__5272 (
            .O(N__22921),
            .I(N__22889));
    LocalMux I__5271 (
            .O(N__22914),
            .I(N__22889));
    LocalMux I__5270 (
            .O(N__22907),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv4 I__5269 (
            .O(N__22904),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv12 I__5268 (
            .O(N__22899),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv4 I__5267 (
            .O(N__22894),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv4 I__5266 (
            .O(N__22889),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    InMux I__5265 (
            .O(N__22878),
            .I(N__22875));
    LocalMux I__5264 (
            .O(N__22875),
            .I(N__22872));
    Span4Mux_h I__5263 (
            .O(N__22872),
            .I(N__22869));
    Odrv4 I__5262 (
            .O(N__22869),
            .I(\Lab_UT.dictrl.N_79_0 ));
    InMux I__5261 (
            .O(N__22866),
            .I(N__22863));
    LocalMux I__5260 (
            .O(N__22863),
            .I(N__22860));
    Span4Mux_v I__5259 (
            .O(N__22860),
            .I(N__22857));
    Odrv4 I__5258 (
            .O(N__22857),
            .I(\Lab_UT.dictrl.N_40_5 ));
    InMux I__5257 (
            .O(N__22854),
            .I(N__22851));
    LocalMux I__5256 (
            .O(N__22851),
            .I(N__22848));
    Odrv4 I__5255 (
            .O(N__22848),
            .I(\Lab_UT.dictrl.g1_2 ));
    InMux I__5254 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__5253 (
            .O(N__22842),
            .I(N__22839));
    Span4Mux_s2_h I__5252 (
            .O(N__22839),
            .I(N__22836));
    Odrv4 I__5251 (
            .O(N__22836),
            .I(\Lab_UT.dictrl.N_40_2 ));
    InMux I__5250 (
            .O(N__22833),
            .I(N__22830));
    LocalMux I__5249 (
            .O(N__22830),
            .I(N__22827));
    Odrv4 I__5248 (
            .O(N__22827),
            .I(\Lab_UT.dictrl.g1_0 ));
    InMux I__5247 (
            .O(N__22824),
            .I(N__22809));
    InMux I__5246 (
            .O(N__22823),
            .I(N__22802));
    InMux I__5245 (
            .O(N__22822),
            .I(N__22802));
    InMux I__5244 (
            .O(N__22821),
            .I(N__22802));
    CascadeMux I__5243 (
            .O(N__22820),
            .I(N__22798));
    InMux I__5242 (
            .O(N__22819),
            .I(N__22795));
    InMux I__5241 (
            .O(N__22818),
            .I(N__22792));
    InMux I__5240 (
            .O(N__22817),
            .I(N__22781));
    InMux I__5239 (
            .O(N__22816),
            .I(N__22781));
    InMux I__5238 (
            .O(N__22815),
            .I(N__22781));
    InMux I__5237 (
            .O(N__22814),
            .I(N__22781));
    InMux I__5236 (
            .O(N__22813),
            .I(N__22781));
    InMux I__5235 (
            .O(N__22812),
            .I(N__22778));
    LocalMux I__5234 (
            .O(N__22809),
            .I(N__22770));
    LocalMux I__5233 (
            .O(N__22802),
            .I(N__22770));
    InMux I__5232 (
            .O(N__22801),
            .I(N__22767));
    InMux I__5231 (
            .O(N__22798),
            .I(N__22762));
    LocalMux I__5230 (
            .O(N__22795),
            .I(N__22759));
    LocalMux I__5229 (
            .O(N__22792),
            .I(N__22756));
    LocalMux I__5228 (
            .O(N__22781),
            .I(N__22751));
    LocalMux I__5227 (
            .O(N__22778),
            .I(N__22751));
    InMux I__5226 (
            .O(N__22777),
            .I(N__22745));
    InMux I__5225 (
            .O(N__22776),
            .I(N__22745));
    InMux I__5224 (
            .O(N__22775),
            .I(N__22742));
    Sp12to4 I__5223 (
            .O(N__22770),
            .I(N__22737));
    LocalMux I__5222 (
            .O(N__22767),
            .I(N__22737));
    InMux I__5221 (
            .O(N__22766),
            .I(N__22734));
    InMux I__5220 (
            .O(N__22765),
            .I(N__22731));
    LocalMux I__5219 (
            .O(N__22762),
            .I(N__22726));
    Span4Mux_s3_v I__5218 (
            .O(N__22759),
            .I(N__22726));
    Span4Mux_v I__5217 (
            .O(N__22756),
            .I(N__22721));
    Span4Mux_s2_h I__5216 (
            .O(N__22751),
            .I(N__22721));
    InMux I__5215 (
            .O(N__22750),
            .I(N__22718));
    LocalMux I__5214 (
            .O(N__22745),
            .I(N__22713));
    LocalMux I__5213 (
            .O(N__22742),
            .I(N__22713));
    Span12Mux_s7_v I__5212 (
            .O(N__22737),
            .I(N__22706));
    LocalMux I__5211 (
            .O(N__22734),
            .I(N__22706));
    LocalMux I__5210 (
            .O(N__22731),
            .I(N__22706));
    Span4Mux_v I__5209 (
            .O(N__22726),
            .I(N__22703));
    Span4Mux_h I__5208 (
            .O(N__22721),
            .I(N__22700));
    LocalMux I__5207 (
            .O(N__22718),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv12 I__5206 (
            .O(N__22713),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv12 I__5205 (
            .O(N__22706),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5204 (
            .O(N__22703),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__5203 (
            .O(N__22700),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    InMux I__5202 (
            .O(N__22689),
            .I(N__22686));
    LocalMux I__5201 (
            .O(N__22686),
            .I(N__22683));
    Span4Mux_s2_h I__5200 (
            .O(N__22683),
            .I(N__22680));
    Span4Mux_v I__5199 (
            .O(N__22680),
            .I(N__22677));
    Odrv4 I__5198 (
            .O(N__22677),
            .I(\Lab_UT.dictrl.N_1460_4 ));
    CascadeMux I__5197 (
            .O(N__22674),
            .I(N__22671));
    InMux I__5196 (
            .O(N__22671),
            .I(N__22668));
    LocalMux I__5195 (
            .O(N__22668),
            .I(N__22665));
    Odrv4 I__5194 (
            .O(N__22665),
            .I(\Lab_UT.dictrl.g2_4 ));
    CascadeMux I__5193 (
            .O(N__22662),
            .I(\Lab_UT.dictrl.next_state_4_1_cascade_ ));
    InMux I__5192 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__5191 (
            .O(N__22656),
            .I(N__22653));
    Odrv4 I__5190 (
            .O(N__22653),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__5189 (
            .O(N__22650),
            .I(N__22647));
    LocalMux I__5188 (
            .O(N__22647),
            .I(\Lab_UT.LdSones_i_4 ));
    InMux I__5187 (
            .O(N__22644),
            .I(N__22638));
    InMux I__5186 (
            .O(N__22643),
            .I(N__22635));
    InMux I__5185 (
            .O(N__22642),
            .I(N__22630));
    InMux I__5184 (
            .O(N__22641),
            .I(N__22630));
    LocalMux I__5183 (
            .O(N__22638),
            .I(N__22627));
    LocalMux I__5182 (
            .O(N__22635),
            .I(N__22624));
    LocalMux I__5181 (
            .O(N__22630),
            .I(N__22621));
    Span4Mux_v I__5180 (
            .O(N__22627),
            .I(N__22618));
    Span4Mux_h I__5179 (
            .O(N__22624),
            .I(N__22615));
    Span4Mux_h I__5178 (
            .O(N__22621),
            .I(N__22612));
    Odrv4 I__5177 (
            .O(N__22618),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    Odrv4 I__5176 (
            .O(N__22615),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    Odrv4 I__5175 (
            .O(N__22612),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    InMux I__5174 (
            .O(N__22605),
            .I(N__22600));
    InMux I__5173 (
            .O(N__22604),
            .I(N__22595));
    InMux I__5172 (
            .O(N__22603),
            .I(N__22595));
    LocalMux I__5171 (
            .O(N__22600),
            .I(N__22590));
    LocalMux I__5170 (
            .O(N__22595),
            .I(N__22590));
    Span4Mux_h I__5169 (
            .O(N__22590),
            .I(N__22584));
    InMux I__5168 (
            .O(N__22589),
            .I(N__22579));
    InMux I__5167 (
            .O(N__22588),
            .I(N__22579));
    InMux I__5166 (
            .O(N__22587),
            .I(N__22576));
    Odrv4 I__5165 (
            .O(N__22584),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    LocalMux I__5164 (
            .O(N__22579),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    LocalMux I__5163 (
            .O(N__22576),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    CascadeMux I__5162 (
            .O(N__22569),
            .I(N__22564));
    CascadeMux I__5161 (
            .O(N__22568),
            .I(N__22561));
    InMux I__5160 (
            .O(N__22567),
            .I(N__22553));
    InMux I__5159 (
            .O(N__22564),
            .I(N__22553));
    InMux I__5158 (
            .O(N__22561),
            .I(N__22553));
    CascadeMux I__5157 (
            .O(N__22560),
            .I(N__22547));
    LocalMux I__5156 (
            .O(N__22553),
            .I(N__22544));
    InMux I__5155 (
            .O(N__22552),
            .I(N__22541));
    InMux I__5154 (
            .O(N__22551),
            .I(N__22538));
    InMux I__5153 (
            .O(N__22550),
            .I(N__22533));
    InMux I__5152 (
            .O(N__22547),
            .I(N__22533));
    Odrv12 I__5151 (
            .O(N__22544),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    LocalMux I__5150 (
            .O(N__22541),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    LocalMux I__5149 (
            .O(N__22538),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    LocalMux I__5148 (
            .O(N__22533),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    CascadeMux I__5147 (
            .O(N__22524),
            .I(N__22518));
    InMux I__5146 (
            .O(N__22523),
            .I(N__22513));
    InMux I__5145 (
            .O(N__22522),
            .I(N__22513));
    InMux I__5144 (
            .O(N__22521),
            .I(N__22508));
    InMux I__5143 (
            .O(N__22518),
            .I(N__22508));
    LocalMux I__5142 (
            .O(N__22513),
            .I(N__22505));
    LocalMux I__5141 (
            .O(N__22508),
            .I(N__22502));
    Span4Mux_h I__5140 (
            .O(N__22505),
            .I(N__22499));
    Span4Mux_h I__5139 (
            .O(N__22502),
            .I(N__22496));
    Odrv4 I__5138 (
            .O(N__22499),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__5137 (
            .O(N__22496),
            .I(\Lab_UT.LdSones ));
    CEMux I__5136 (
            .O(N__22491),
            .I(N__22473));
    CEMux I__5135 (
            .O(N__22490),
            .I(N__22473));
    CEMux I__5134 (
            .O(N__22489),
            .I(N__22473));
    CEMux I__5133 (
            .O(N__22488),
            .I(N__22473));
    CEMux I__5132 (
            .O(N__22487),
            .I(N__22473));
    CEMux I__5131 (
            .O(N__22486),
            .I(N__22473));
    GlobalMux I__5130 (
            .O(N__22473),
            .I(N__22470));
    gio2CtrlBuf I__5129 (
            .O(N__22470),
            .I(bu_rx_data_rdy_0_g));
    CascadeMux I__5128 (
            .O(N__22467),
            .I(N__22464));
    InMux I__5127 (
            .O(N__22464),
            .I(N__22459));
    CascadeMux I__5126 (
            .O(N__22463),
            .I(N__22455));
    CascadeMux I__5125 (
            .O(N__22462),
            .I(N__22452));
    LocalMux I__5124 (
            .O(N__22459),
            .I(N__22449));
    InMux I__5123 (
            .O(N__22458),
            .I(N__22442));
    InMux I__5122 (
            .O(N__22455),
            .I(N__22442));
    InMux I__5121 (
            .O(N__22452),
            .I(N__22442));
    Span4Mux_v I__5120 (
            .O(N__22449),
            .I(N__22439));
    LocalMux I__5119 (
            .O(N__22442),
            .I(N__22436));
    Span4Mux_h I__5118 (
            .O(N__22439),
            .I(N__22433));
    Span4Mux_h I__5117 (
            .O(N__22436),
            .I(N__22430));
    Odrv4 I__5116 (
            .O(N__22433),
            .I(\Lab_UT.dictrl.g2_5 ));
    Odrv4 I__5115 (
            .O(N__22430),
            .I(\Lab_UT.dictrl.g2_5 ));
    InMux I__5114 (
            .O(N__22425),
            .I(N__22422));
    LocalMux I__5113 (
            .O(N__22422),
            .I(N__22415));
    InMux I__5112 (
            .O(N__22421),
            .I(N__22408));
    InMux I__5111 (
            .O(N__22420),
            .I(N__22408));
    InMux I__5110 (
            .O(N__22419),
            .I(N__22408));
    InMux I__5109 (
            .O(N__22418),
            .I(N__22405));
    Span4Mux_v I__5108 (
            .O(N__22415),
            .I(N__22402));
    LocalMux I__5107 (
            .O(N__22408),
            .I(N__22399));
    LocalMux I__5106 (
            .O(N__22405),
            .I(N__22396));
    Span4Mux_v I__5105 (
            .O(N__22402),
            .I(N__22393));
    Span4Mux_h I__5104 (
            .O(N__22399),
            .I(N__22388));
    Span4Mux_s2_h I__5103 (
            .O(N__22396),
            .I(N__22388));
    Odrv4 I__5102 (
            .O(N__22393),
            .I(\Lab_UT.dictrl.g1_3 ));
    Odrv4 I__5101 (
            .O(N__22388),
            .I(\Lab_UT.dictrl.g1_3 ));
    CascadeMux I__5100 (
            .O(N__22383),
            .I(\Lab_UT.dictrl.g2_5_cascade_ ));
    InMux I__5099 (
            .O(N__22380),
            .I(N__22376));
    CascadeMux I__5098 (
            .O(N__22379),
            .I(N__22373));
    LocalMux I__5097 (
            .O(N__22376),
            .I(N__22367));
    InMux I__5096 (
            .O(N__22373),
            .I(N__22360));
    InMux I__5095 (
            .O(N__22372),
            .I(N__22360));
    InMux I__5094 (
            .O(N__22371),
            .I(N__22360));
    InMux I__5093 (
            .O(N__22370),
            .I(N__22357));
    Span4Mux_h I__5092 (
            .O(N__22367),
            .I(N__22354));
    LocalMux I__5091 (
            .O(N__22360),
            .I(N__22351));
    LocalMux I__5090 (
            .O(N__22357),
            .I(N__22348));
    Span4Mux_v I__5089 (
            .O(N__22354),
            .I(N__22345));
    Span4Mux_h I__5088 (
            .O(N__22351),
            .I(N__22340));
    Span4Mux_s2_h I__5087 (
            .O(N__22348),
            .I(N__22340));
    Odrv4 I__5086 (
            .O(N__22345),
            .I(\Lab_UT.dictrl.N_1460_5 ));
    Odrv4 I__5085 (
            .O(N__22340),
            .I(\Lab_UT.dictrl.N_1460_5 ));
    InMux I__5084 (
            .O(N__22335),
            .I(N__22329));
    InMux I__5083 (
            .O(N__22334),
            .I(N__22329));
    LocalMux I__5082 (
            .O(N__22329),
            .I(N__22326));
    Span4Mux_h I__5081 (
            .O(N__22326),
            .I(N__22323));
    Odrv4 I__5080 (
            .O(N__22323),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    InMux I__5079 (
            .O(N__22320),
            .I(N__22316));
    InMux I__5078 (
            .O(N__22319),
            .I(N__22313));
    LocalMux I__5077 (
            .O(N__22316),
            .I(N__22308));
    LocalMux I__5076 (
            .O(N__22313),
            .I(N__22308));
    Odrv4 I__5075 (
            .O(N__22308),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    CascadeMux I__5074 (
            .O(N__22305),
            .I(N__22299));
    InMux I__5073 (
            .O(N__22304),
            .I(N__22287));
    InMux I__5072 (
            .O(N__22303),
            .I(N__22287));
    InMux I__5071 (
            .O(N__22302),
            .I(N__22287));
    InMux I__5070 (
            .O(N__22299),
            .I(N__22287));
    InMux I__5069 (
            .O(N__22298),
            .I(N__22287));
    LocalMux I__5068 (
            .O(N__22287),
            .I(N__22284));
    Odrv12 I__5067 (
            .O(N__22284),
            .I(\Lab_UT.didp.un24_ce_2 ));
    InMux I__5066 (
            .O(N__22281),
            .I(N__22276));
    InMux I__5065 (
            .O(N__22280),
            .I(N__22273));
    InMux I__5064 (
            .O(N__22279),
            .I(N__22270));
    LocalMux I__5063 (
            .O(N__22276),
            .I(N__22263));
    LocalMux I__5062 (
            .O(N__22273),
            .I(N__22260));
    LocalMux I__5061 (
            .O(N__22270),
            .I(N__22257));
    InMux I__5060 (
            .O(N__22269),
            .I(N__22254));
    InMux I__5059 (
            .O(N__22268),
            .I(N__22251));
    InMux I__5058 (
            .O(N__22267),
            .I(N__22248));
    InMux I__5057 (
            .O(N__22266),
            .I(N__22245));
    Span4Mux_h I__5056 (
            .O(N__22263),
            .I(N__22242));
    Span4Mux_s3_h I__5055 (
            .O(N__22260),
            .I(N__22237));
    Span4Mux_h I__5054 (
            .O(N__22257),
            .I(N__22237));
    LocalMux I__5053 (
            .O(N__22254),
            .I(N__22234));
    LocalMux I__5052 (
            .O(N__22251),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__5051 (
            .O(N__22248),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__5050 (
            .O(N__22245),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__5049 (
            .O(N__22242),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__5048 (
            .O(N__22237),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__5047 (
            .O(N__22234),
            .I(\Lab_UT.di_Mtens_1 ));
    CascadeMux I__5046 (
            .O(N__22221),
            .I(\Lab_UT.didp.ce_12_3_cascade_ ));
    InMux I__5045 (
            .O(N__22218),
            .I(N__22215));
    LocalMux I__5044 (
            .O(N__22215),
            .I(N__22210));
    CascadeMux I__5043 (
            .O(N__22214),
            .I(N__22205));
    InMux I__5042 (
            .O(N__22213),
            .I(N__22202));
    Span4Mux_h I__5041 (
            .O(N__22210),
            .I(N__22199));
    InMux I__5040 (
            .O(N__22209),
            .I(N__22192));
    InMux I__5039 (
            .O(N__22208),
            .I(N__22192));
    InMux I__5038 (
            .O(N__22205),
            .I(N__22192));
    LocalMux I__5037 (
            .O(N__22202),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__5036 (
            .O(N__22199),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__5035 (
            .O(N__22192),
            .I(\Lab_UT.di_Mtens_3 ));
    InMux I__5034 (
            .O(N__22185),
            .I(N__22179));
    InMux I__5033 (
            .O(N__22184),
            .I(N__22179));
    LocalMux I__5032 (
            .O(N__22179),
            .I(N__22174));
    InMux I__5031 (
            .O(N__22178),
            .I(N__22171));
    InMux I__5030 (
            .O(N__22177),
            .I(N__22168));
    Span4Mux_v I__5029 (
            .O(N__22174),
            .I(N__22165));
    LocalMux I__5028 (
            .O(N__22171),
            .I(N__22160));
    LocalMux I__5027 (
            .O(N__22168),
            .I(N__22160));
    Span4Mux_h I__5026 (
            .O(N__22165),
            .I(N__22157));
    Span4Mux_h I__5025 (
            .O(N__22160),
            .I(N__22154));
    Odrv4 I__5024 (
            .O(N__22157),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    Odrv4 I__5023 (
            .O(N__22154),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    InMux I__5022 (
            .O(N__22149),
            .I(N__22130));
    InMux I__5021 (
            .O(N__22148),
            .I(N__22130));
    InMux I__5020 (
            .O(N__22147),
            .I(N__22130));
    InMux I__5019 (
            .O(N__22146),
            .I(N__22130));
    InMux I__5018 (
            .O(N__22145),
            .I(N__22130));
    InMux I__5017 (
            .O(N__22144),
            .I(N__22130));
    InMux I__5016 (
            .O(N__22143),
            .I(N__22127));
    LocalMux I__5015 (
            .O(N__22130),
            .I(N__22124));
    LocalMux I__5014 (
            .O(N__22127),
            .I(N__22121));
    Span4Mux_s2_h I__5013 (
            .O(N__22124),
            .I(N__22118));
    Odrv12 I__5012 (
            .O(N__22121),
            .I(\Lab_UT.didp.un18_ce ));
    Odrv4 I__5011 (
            .O(N__22118),
            .I(\Lab_UT.didp.un18_ce ));
    CascadeMux I__5010 (
            .O(N__22113),
            .I(N__22105));
    CascadeMux I__5009 (
            .O(N__22112),
            .I(N__22102));
    CascadeMux I__5008 (
            .O(N__22111),
            .I(N__22099));
    CascadeMux I__5007 (
            .O(N__22110),
            .I(N__22096));
    CascadeMux I__5006 (
            .O(N__22109),
            .I(N__22091));
    InMux I__5005 (
            .O(N__22108),
            .I(N__22084));
    InMux I__5004 (
            .O(N__22105),
            .I(N__22084));
    InMux I__5003 (
            .O(N__22102),
            .I(N__22071));
    InMux I__5002 (
            .O(N__22099),
            .I(N__22071));
    InMux I__5001 (
            .O(N__22096),
            .I(N__22071));
    InMux I__5000 (
            .O(N__22095),
            .I(N__22071));
    InMux I__4999 (
            .O(N__22094),
            .I(N__22071));
    InMux I__4998 (
            .O(N__22091),
            .I(N__22071));
    CascadeMux I__4997 (
            .O(N__22090),
            .I(N__22066));
    InMux I__4996 (
            .O(N__22089),
            .I(N__22062));
    LocalMux I__4995 (
            .O(N__22084),
            .I(N__22059));
    LocalMux I__4994 (
            .O(N__22071),
            .I(N__22056));
    CascadeMux I__4993 (
            .O(N__22070),
            .I(N__22053));
    InMux I__4992 (
            .O(N__22069),
            .I(N__22047));
    InMux I__4991 (
            .O(N__22066),
            .I(N__22047));
    CascadeMux I__4990 (
            .O(N__22065),
            .I(N__22044));
    LocalMux I__4989 (
            .O(N__22062),
            .I(N__22041));
    Span4Mux_v I__4988 (
            .O(N__22059),
            .I(N__22036));
    Span4Mux_s2_h I__4987 (
            .O(N__22056),
            .I(N__22036));
    InMux I__4986 (
            .O(N__22053),
            .I(N__22031));
    InMux I__4985 (
            .O(N__22052),
            .I(N__22028));
    LocalMux I__4984 (
            .O(N__22047),
            .I(N__22025));
    InMux I__4983 (
            .O(N__22044),
            .I(N__22022));
    Span4Mux_h I__4982 (
            .O(N__22041),
            .I(N__22017));
    Span4Mux_h I__4981 (
            .O(N__22036),
            .I(N__22017));
    InMux I__4980 (
            .O(N__22035),
            .I(N__22012));
    InMux I__4979 (
            .O(N__22034),
            .I(N__22012));
    LocalMux I__4978 (
            .O(N__22031),
            .I(oneSecStrb));
    LocalMux I__4977 (
            .O(N__22028),
            .I(oneSecStrb));
    Odrv4 I__4976 (
            .O(N__22025),
            .I(oneSecStrb));
    LocalMux I__4975 (
            .O(N__22022),
            .I(oneSecStrb));
    Odrv4 I__4974 (
            .O(N__22017),
            .I(oneSecStrb));
    LocalMux I__4973 (
            .O(N__22012),
            .I(oneSecStrb));
    CascadeMux I__4972 (
            .O(N__21999),
            .I(N__21994));
    InMux I__4971 (
            .O(N__21998),
            .I(N__21987));
    InMux I__4970 (
            .O(N__21997),
            .I(N__21987));
    InMux I__4969 (
            .O(N__21994),
            .I(N__21987));
    LocalMux I__4968 (
            .O(N__21987),
            .I(N__21983));
    InMux I__4967 (
            .O(N__21986),
            .I(N__21980));
    Span12Mux_s7_v I__4966 (
            .O(N__21983),
            .I(N__21975));
    LocalMux I__4965 (
            .O(N__21980),
            .I(N__21975));
    Odrv12 I__4964 (
            .O(N__21975),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    InMux I__4963 (
            .O(N__21972),
            .I(N__21967));
    InMux I__4962 (
            .O(N__21971),
            .I(N__21964));
    InMux I__4961 (
            .O(N__21970),
            .I(N__21961));
    LocalMux I__4960 (
            .O(N__21967),
            .I(N__21956));
    LocalMux I__4959 (
            .O(N__21964),
            .I(N__21953));
    LocalMux I__4958 (
            .O(N__21961),
            .I(N__21949));
    InMux I__4957 (
            .O(N__21960),
            .I(N__21943));
    InMux I__4956 (
            .O(N__21959),
            .I(N__21943));
    Span4Mux_v I__4955 (
            .O(N__21956),
            .I(N__21938));
    Span4Mux_v I__4954 (
            .O(N__21953),
            .I(N__21938));
    InMux I__4953 (
            .O(N__21952),
            .I(N__21935));
    Span4Mux_h I__4952 (
            .O(N__21949),
            .I(N__21932));
    InMux I__4951 (
            .O(N__21948),
            .I(N__21929));
    LocalMux I__4950 (
            .O(N__21943),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__4949 (
            .O(N__21938),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4948 (
            .O(N__21935),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__4947 (
            .O(N__21932),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4946 (
            .O(N__21929),
            .I(\Lab_UT.di_Mtens_0 ));
    InMux I__4945 (
            .O(N__21918),
            .I(N__21915));
    LocalMux I__4944 (
            .O(N__21915),
            .I(N__21911));
    InMux I__4943 (
            .O(N__21914),
            .I(N__21908));
    Span4Mux_v I__4942 (
            .O(N__21911),
            .I(N__21899));
    LocalMux I__4941 (
            .O(N__21908),
            .I(N__21899));
    InMux I__4940 (
            .O(N__21907),
            .I(N__21896));
    InMux I__4939 (
            .O(N__21906),
            .I(N__21889));
    InMux I__4938 (
            .O(N__21905),
            .I(N__21889));
    InMux I__4937 (
            .O(N__21904),
            .I(N__21889));
    Odrv4 I__4936 (
            .O(N__21899),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__4935 (
            .O(N__21896),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__4934 (
            .O(N__21889),
            .I(\Lab_UT.di_Mtens_2 ));
    InMux I__4933 (
            .O(N__21882),
            .I(N__21879));
    LocalMux I__4932 (
            .O(N__21879),
            .I(\Lab_UT.didp.reset_12_1_3 ));
    InMux I__4931 (
            .O(N__21876),
            .I(N__21873));
    LocalMux I__4930 (
            .O(N__21873),
            .I(N__21870));
    Span4Mux_s2_h I__4929 (
            .O(N__21870),
            .I(N__21867));
    Odrv4 I__4928 (
            .O(N__21867),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__4927 (
            .O(N__21864),
            .I(N__21861));
    LocalMux I__4926 (
            .O(N__21861),
            .I(N__21858));
    Span4Mux_s3_h I__4925 (
            .O(N__21858),
            .I(N__21855));
    Odrv4 I__4924 (
            .O(N__21855),
            .I(\Lab_UT.LdStens_i_4 ));
    InMux I__4923 (
            .O(N__21852),
            .I(N__21849));
    LocalMux I__4922 (
            .O(N__21849),
            .I(N__21844));
    InMux I__4921 (
            .O(N__21848),
            .I(N__21839));
    InMux I__4920 (
            .O(N__21847),
            .I(N__21839));
    Span4Mux_v I__4919 (
            .O(N__21844),
            .I(N__21834));
    LocalMux I__4918 (
            .O(N__21839),
            .I(N__21834));
    Span4Mux_h I__4917 (
            .O(N__21834),
            .I(N__21831));
    Odrv4 I__4916 (
            .O(N__21831),
            .I(\Lab_UT.di_AMones_3 ));
    CEMux I__4915 (
            .O(N__21828),
            .I(N__21825));
    LocalMux I__4914 (
            .O(N__21825),
            .I(N__21822));
    Span4Mux_v I__4913 (
            .O(N__21822),
            .I(N__21818));
    CEMux I__4912 (
            .O(N__21821),
            .I(N__21815));
    Span4Mux_s1_h I__4911 (
            .O(N__21818),
            .I(N__21810));
    LocalMux I__4910 (
            .O(N__21815),
            .I(N__21810));
    Odrv4 I__4909 (
            .O(N__21810),
            .I(\Lab_UT.didp.regrce3.LdAMones_0 ));
    InMux I__4908 (
            .O(N__21807),
            .I(N__21799));
    InMux I__4907 (
            .O(N__21806),
            .I(N__21796));
    InMux I__4906 (
            .O(N__21805),
            .I(N__21793));
    InMux I__4905 (
            .O(N__21804),
            .I(N__21790));
    InMux I__4904 (
            .O(N__21803),
            .I(N__21787));
    InMux I__4903 (
            .O(N__21802),
            .I(N__21783));
    LocalMux I__4902 (
            .O(N__21799),
            .I(N__21780));
    LocalMux I__4901 (
            .O(N__21796),
            .I(N__21776));
    LocalMux I__4900 (
            .O(N__21793),
            .I(N__21771));
    LocalMux I__4899 (
            .O(N__21790),
            .I(N__21767));
    LocalMux I__4898 (
            .O(N__21787),
            .I(N__21764));
    InMux I__4897 (
            .O(N__21786),
            .I(N__21761));
    LocalMux I__4896 (
            .O(N__21783),
            .I(N__21756));
    Span4Mux_s2_h I__4895 (
            .O(N__21780),
            .I(N__21756));
    InMux I__4894 (
            .O(N__21779),
            .I(N__21753));
    Span4Mux_s2_h I__4893 (
            .O(N__21776),
            .I(N__21750));
    InMux I__4892 (
            .O(N__21775),
            .I(N__21746));
    InMux I__4891 (
            .O(N__21774),
            .I(N__21743));
    Span4Mux_h I__4890 (
            .O(N__21771),
            .I(N__21740));
    InMux I__4889 (
            .O(N__21770),
            .I(N__21737));
    Span4Mux_v I__4888 (
            .O(N__21767),
            .I(N__21730));
    Span4Mux_v I__4887 (
            .O(N__21764),
            .I(N__21730));
    LocalMux I__4886 (
            .O(N__21761),
            .I(N__21730));
    Span4Mux_h I__4885 (
            .O(N__21756),
            .I(N__21725));
    LocalMux I__4884 (
            .O(N__21753),
            .I(N__21725));
    Span4Mux_h I__4883 (
            .O(N__21750),
            .I(N__21722));
    InMux I__4882 (
            .O(N__21749),
            .I(N__21719));
    LocalMux I__4881 (
            .O(N__21746),
            .I(N__21714));
    LocalMux I__4880 (
            .O(N__21743),
            .I(N__21714));
    Span4Mux_v I__4879 (
            .O(N__21740),
            .I(N__21711));
    LocalMux I__4878 (
            .O(N__21737),
            .I(N__21704));
    Span4Mux_h I__4877 (
            .O(N__21730),
            .I(N__21704));
    Span4Mux_h I__4876 (
            .O(N__21725),
            .I(N__21701));
    Span4Mux_v I__4875 (
            .O(N__21722),
            .I(N__21696));
    LocalMux I__4874 (
            .O(N__21719),
            .I(N__21696));
    Span12Mux_s10_h I__4873 (
            .O(N__21714),
            .I(N__21693));
    Span4Mux_h I__4872 (
            .O(N__21711),
            .I(N__21690));
    InMux I__4871 (
            .O(N__21710),
            .I(N__21685));
    InMux I__4870 (
            .O(N__21709),
            .I(N__21685));
    Span4Mux_h I__4869 (
            .O(N__21704),
            .I(N__21680));
    Span4Mux_v I__4868 (
            .O(N__21701),
            .I(N__21680));
    Span4Mux_h I__4867 (
            .O(N__21696),
            .I(N__21677));
    Odrv12 I__4866 (
            .O(N__21693),
            .I(bu_rx_data_0));
    Odrv4 I__4865 (
            .O(N__21690),
            .I(bu_rx_data_0));
    LocalMux I__4864 (
            .O(N__21685),
            .I(bu_rx_data_0));
    Odrv4 I__4863 (
            .O(N__21680),
            .I(bu_rx_data_0));
    Odrv4 I__4862 (
            .O(N__21677),
            .I(bu_rx_data_0));
    InMux I__4861 (
            .O(N__21666),
            .I(N__21663));
    LocalMux I__4860 (
            .O(N__21663),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    CascadeMux I__4859 (
            .O(N__21660),
            .I(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ));
    InMux I__4858 (
            .O(N__21657),
            .I(N__21654));
    LocalMux I__4857 (
            .O(N__21654),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    InMux I__4856 (
            .O(N__21651),
            .I(N__21647));
    InMux I__4855 (
            .O(N__21650),
            .I(N__21644));
    LocalMux I__4854 (
            .O(N__21647),
            .I(N__21641));
    LocalMux I__4853 (
            .O(N__21644),
            .I(N__21637));
    Span4Mux_v I__4852 (
            .O(N__21641),
            .I(N__21634));
    InMux I__4851 (
            .O(N__21640),
            .I(N__21631));
    Odrv12 I__4850 (
            .O(N__21637),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__4849 (
            .O(N__21634),
            .I(\Lab_UT.di_AMones_2 ));
    LocalMux I__4848 (
            .O(N__21631),
            .I(\Lab_UT.di_AMones_2 ));
    InMux I__4847 (
            .O(N__21624),
            .I(N__21621));
    LocalMux I__4846 (
            .O(N__21621),
            .I(N__21617));
    InMux I__4845 (
            .O(N__21620),
            .I(N__21614));
    Span4Mux_v I__4844 (
            .O(N__21617),
            .I(N__21610));
    LocalMux I__4843 (
            .O(N__21614),
            .I(N__21607));
    CascadeMux I__4842 (
            .O(N__21613),
            .I(N__21604));
    Span4Mux_h I__4841 (
            .O(N__21610),
            .I(N__21601));
    Span4Mux_v I__4840 (
            .O(N__21607),
            .I(N__21598));
    InMux I__4839 (
            .O(N__21604),
            .I(N__21595));
    Odrv4 I__4838 (
            .O(N__21601),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__4837 (
            .O(N__21598),
            .I(\Lab_UT.di_AMones_1 ));
    LocalMux I__4836 (
            .O(N__21595),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__4835 (
            .O(N__21588),
            .I(N__21585));
    LocalMux I__4834 (
            .O(N__21585),
            .I(N__21582));
    Odrv4 I__4833 (
            .O(N__21582),
            .I(\Lab_UT.dispString.m49Z0Z_2 ));
    CascadeMux I__4832 (
            .O(N__21579),
            .I(N__21575));
    CascadeMux I__4831 (
            .O(N__21578),
            .I(N__21572));
    InMux I__4830 (
            .O(N__21575),
            .I(N__21562));
    InMux I__4829 (
            .O(N__21572),
            .I(N__21562));
    InMux I__4828 (
            .O(N__21571),
            .I(N__21562));
    InMux I__4827 (
            .O(N__21570),
            .I(N__21557));
    InMux I__4826 (
            .O(N__21569),
            .I(N__21557));
    LocalMux I__4825 (
            .O(N__21562),
            .I(N__21554));
    LocalMux I__4824 (
            .O(N__21557),
            .I(N__21551));
    Span4Mux_s3_h I__4823 (
            .O(N__21554),
            .I(N__21546));
    Span4Mux_s3_h I__4822 (
            .O(N__21551),
            .I(N__21543));
    InMux I__4821 (
            .O(N__21550),
            .I(N__21538));
    InMux I__4820 (
            .O(N__21549),
            .I(N__21538));
    Odrv4 I__4819 (
            .O(N__21546),
            .I(\Lab_UT.sec2_1 ));
    Odrv4 I__4818 (
            .O(N__21543),
            .I(\Lab_UT.sec2_1 ));
    LocalMux I__4817 (
            .O(N__21538),
            .I(\Lab_UT.sec2_1 ));
    CascadeMux I__4816 (
            .O(N__21531),
            .I(N__21526));
    InMux I__4815 (
            .O(N__21530),
            .I(N__21518));
    InMux I__4814 (
            .O(N__21529),
            .I(N__21518));
    InMux I__4813 (
            .O(N__21526),
            .I(N__21518));
    CascadeMux I__4812 (
            .O(N__21525),
            .I(N__21514));
    LocalMux I__4811 (
            .O(N__21518),
            .I(N__21510));
    InMux I__4810 (
            .O(N__21517),
            .I(N__21505));
    InMux I__4809 (
            .O(N__21514),
            .I(N__21505));
    CascadeMux I__4808 (
            .O(N__21513),
            .I(N__21501));
    Span4Mux_v I__4807 (
            .O(N__21510),
            .I(N__21498));
    LocalMux I__4806 (
            .O(N__21505),
            .I(N__21495));
    InMux I__4805 (
            .O(N__21504),
            .I(N__21490));
    InMux I__4804 (
            .O(N__21501),
            .I(N__21490));
    Span4Mux_s1_h I__4803 (
            .O(N__21498),
            .I(N__21485));
    Span4Mux_v I__4802 (
            .O(N__21495),
            .I(N__21485));
    LocalMux I__4801 (
            .O(N__21490),
            .I(N__21482));
    Odrv4 I__4800 (
            .O(N__21485),
            .I(\Lab_UT.sec2_3 ));
    Odrv4 I__4799 (
            .O(N__21482),
            .I(\Lab_UT.sec2_3 ));
    CascadeMux I__4798 (
            .O(N__21477),
            .I(N__21471));
    InMux I__4797 (
            .O(N__21476),
            .I(N__21463));
    InMux I__4796 (
            .O(N__21475),
            .I(N__21463));
    InMux I__4795 (
            .O(N__21474),
            .I(N__21463));
    InMux I__4794 (
            .O(N__21471),
            .I(N__21458));
    InMux I__4793 (
            .O(N__21470),
            .I(N__21458));
    LocalMux I__4792 (
            .O(N__21463),
            .I(N__21454));
    LocalMux I__4791 (
            .O(N__21458),
            .I(N__21451));
    CascadeMux I__4790 (
            .O(N__21457),
            .I(N__21448));
    Span4Mux_s2_h I__4789 (
            .O(N__21454),
            .I(N__21444));
    Span4Mux_s2_h I__4788 (
            .O(N__21451),
            .I(N__21441));
    InMux I__4787 (
            .O(N__21448),
            .I(N__21436));
    InMux I__4786 (
            .O(N__21447),
            .I(N__21436));
    Odrv4 I__4785 (
            .O(N__21444),
            .I(\Lab_UT.sec2_2 ));
    Odrv4 I__4784 (
            .O(N__21441),
            .I(\Lab_UT.sec2_2 ));
    LocalMux I__4783 (
            .O(N__21436),
            .I(\Lab_UT.sec2_2 ));
    InMux I__4782 (
            .O(N__21429),
            .I(N__21423));
    InMux I__4781 (
            .O(N__21428),
            .I(N__21423));
    LocalMux I__4780 (
            .O(N__21423),
            .I(N__21417));
    InMux I__4779 (
            .O(N__21422),
            .I(N__21410));
    InMux I__4778 (
            .O(N__21421),
            .I(N__21410));
    InMux I__4777 (
            .O(N__21420),
            .I(N__21410));
    Span4Mux_v I__4776 (
            .O(N__21417),
            .I(N__21405));
    LocalMux I__4775 (
            .O(N__21410),
            .I(N__21402));
    InMux I__4774 (
            .O(N__21409),
            .I(N__21397));
    InMux I__4773 (
            .O(N__21408),
            .I(N__21397));
    Sp12to4 I__4772 (
            .O(N__21405),
            .I(N__21394));
    Span4Mux_s3_h I__4771 (
            .O(N__21402),
            .I(N__21389));
    LocalMux I__4770 (
            .O(N__21397),
            .I(N__21389));
    Odrv12 I__4769 (
            .O(N__21394),
            .I(\Lab_UT.sec2_0 ));
    Odrv4 I__4768 (
            .O(N__21389),
            .I(\Lab_UT.sec2_0 ));
    InMux I__4767 (
            .O(N__21384),
            .I(N__21381));
    LocalMux I__4766 (
            .O(N__21381),
            .I(\uu2.bitmapZ0Z_58 ));
    CascadeMux I__4765 (
            .O(N__21378),
            .I(\Lab_UT.didp.countrce2.q_5_0_cascade_ ));
    InMux I__4764 (
            .O(N__21375),
            .I(N__21371));
    InMux I__4763 (
            .O(N__21374),
            .I(N__21368));
    LocalMux I__4762 (
            .O(N__21371),
            .I(N__21365));
    LocalMux I__4761 (
            .O(N__21368),
            .I(N__21362));
    Span4Mux_h I__4760 (
            .O(N__21365),
            .I(N__21356));
    Span4Mux_v I__4759 (
            .O(N__21362),
            .I(N__21356));
    InMux I__4758 (
            .O(N__21361),
            .I(N__21353));
    Odrv4 I__4757 (
            .O(N__21356),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__4756 (
            .O(N__21353),
            .I(\Lab_UT.di_AStens_0 ));
    CascadeMux I__4755 (
            .O(N__21348),
            .I(N__21337));
    InMux I__4754 (
            .O(N__21347),
            .I(N__21333));
    InMux I__4753 (
            .O(N__21346),
            .I(N__21328));
    InMux I__4752 (
            .O(N__21345),
            .I(N__21328));
    InMux I__4751 (
            .O(N__21344),
            .I(N__21321));
    InMux I__4750 (
            .O(N__21343),
            .I(N__21321));
    InMux I__4749 (
            .O(N__21342),
            .I(N__21318));
    InMux I__4748 (
            .O(N__21341),
            .I(N__21309));
    InMux I__4747 (
            .O(N__21340),
            .I(N__21309));
    InMux I__4746 (
            .O(N__21337),
            .I(N__21309));
    InMux I__4745 (
            .O(N__21336),
            .I(N__21309));
    LocalMux I__4744 (
            .O(N__21333),
            .I(N__21304));
    LocalMux I__4743 (
            .O(N__21328),
            .I(N__21304));
    InMux I__4742 (
            .O(N__21327),
            .I(N__21298));
    InMux I__4741 (
            .O(N__21326),
            .I(N__21295));
    LocalMux I__4740 (
            .O(N__21321),
            .I(N__21288));
    LocalMux I__4739 (
            .O(N__21318),
            .I(N__21288));
    LocalMux I__4738 (
            .O(N__21309),
            .I(N__21288));
    Span4Mux_s3_h I__4737 (
            .O(N__21304),
            .I(N__21285));
    InMux I__4736 (
            .O(N__21303),
            .I(N__21282));
    InMux I__4735 (
            .O(N__21302),
            .I(N__21277));
    InMux I__4734 (
            .O(N__21301),
            .I(N__21277));
    LocalMux I__4733 (
            .O(N__21298),
            .I(\Lab_UT.loadalarm_0 ));
    LocalMux I__4732 (
            .O(N__21295),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv4 I__4731 (
            .O(N__21288),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv4 I__4730 (
            .O(N__21285),
            .I(\Lab_UT.loadalarm_0 ));
    LocalMux I__4729 (
            .O(N__21282),
            .I(\Lab_UT.loadalarm_0 ));
    LocalMux I__4728 (
            .O(N__21277),
            .I(\Lab_UT.loadalarm_0 ));
    InMux I__4727 (
            .O(N__21264),
            .I(N__21260));
    InMux I__4726 (
            .O(N__21263),
            .I(N__21252));
    LocalMux I__4725 (
            .O(N__21260),
            .I(N__21249));
    InMux I__4724 (
            .O(N__21259),
            .I(N__21240));
    InMux I__4723 (
            .O(N__21258),
            .I(N__21240));
    InMux I__4722 (
            .O(N__21257),
            .I(N__21240));
    InMux I__4721 (
            .O(N__21256),
            .I(N__21240));
    InMux I__4720 (
            .O(N__21255),
            .I(N__21237));
    LocalMux I__4719 (
            .O(N__21252),
            .I(N__21232));
    Span4Mux_s2_h I__4718 (
            .O(N__21249),
            .I(N__21232));
    LocalMux I__4717 (
            .O(N__21240),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__4716 (
            .O(N__21237),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__4715 (
            .O(N__21232),
            .I(\Lab_UT.di_Sones_1 ));
    InMux I__4714 (
            .O(N__21225),
            .I(N__21222));
    LocalMux I__4713 (
            .O(N__21222),
            .I(N__21217));
    InMux I__4712 (
            .O(N__21221),
            .I(N__21212));
    InMux I__4711 (
            .O(N__21220),
            .I(N__21212));
    Span4Mux_v I__4710 (
            .O(N__21217),
            .I(N__21209));
    LocalMux I__4709 (
            .O(N__21212),
            .I(N__21206));
    Span4Mux_h I__4708 (
            .O(N__21209),
            .I(N__21203));
    Span4Mux_v I__4707 (
            .O(N__21206),
            .I(N__21200));
    Odrv4 I__4706 (
            .O(N__21203),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__4705 (
            .O(N__21200),
            .I(\Lab_UT.di_AStens_1 ));
    InMux I__4704 (
            .O(N__21195),
            .I(N__21191));
    InMux I__4703 (
            .O(N__21194),
            .I(N__21187));
    LocalMux I__4702 (
            .O(N__21191),
            .I(N__21184));
    InMux I__4701 (
            .O(N__21190),
            .I(N__21181));
    LocalMux I__4700 (
            .O(N__21187),
            .I(N__21178));
    Odrv4 I__4699 (
            .O(N__21184),
            .I(\Lab_UT.di_ASones_1 ));
    LocalMux I__4698 (
            .O(N__21181),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__4697 (
            .O(N__21178),
            .I(\Lab_UT.di_ASones_1 ));
    InMux I__4696 (
            .O(N__21171),
            .I(N__21168));
    LocalMux I__4695 (
            .O(N__21168),
            .I(N__21165));
    Span4Mux_h I__4694 (
            .O(N__21165),
            .I(N__21162));
    Odrv4 I__4693 (
            .O(N__21162),
            .I(\Lab_UT.dispString.m49Z0Z_5 ));
    InMux I__4692 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__4691 (
            .O(N__21156),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__4690 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__4689 (
            .O(N__21150),
            .I(\uu2.bitmapZ0Z_90 ));
    InMux I__4688 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__4687 (
            .O(N__21144),
            .I(N__21141));
    Span4Mux_h I__4686 (
            .O(N__21141),
            .I(N__21138));
    Odrv4 I__4685 (
            .O(N__21138),
            .I(\uu2.N_20 ));
    InMux I__4684 (
            .O(N__21135),
            .I(N__21128));
    InMux I__4683 (
            .O(N__21134),
            .I(N__21121));
    InMux I__4682 (
            .O(N__21133),
            .I(N__21121));
    InMux I__4681 (
            .O(N__21132),
            .I(N__21118));
    InMux I__4680 (
            .O(N__21131),
            .I(N__21115));
    LocalMux I__4679 (
            .O(N__21128),
            .I(N__21112));
    InMux I__4678 (
            .O(N__21127),
            .I(N__21109));
    InMux I__4677 (
            .O(N__21126),
            .I(N__21106));
    LocalMux I__4676 (
            .O(N__21121),
            .I(N__21103));
    LocalMux I__4675 (
            .O(N__21118),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__4674 (
            .O(N__21115),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__4673 (
            .O(N__21112),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__4672 (
            .O(N__21109),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__4671 (
            .O(N__21106),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__4670 (
            .O(N__21103),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    CascadeMux I__4669 (
            .O(N__21090),
            .I(\uu2.bitmap_RNIE7RKZ0Z_58_cascade_ ));
    InMux I__4668 (
            .O(N__21087),
            .I(N__21084));
    LocalMux I__4667 (
            .O(N__21084),
            .I(\uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7 ));
    InMux I__4666 (
            .O(N__21081),
            .I(N__21076));
    InMux I__4665 (
            .O(N__21080),
            .I(N__21073));
    InMux I__4664 (
            .O(N__21079),
            .I(N__21070));
    LocalMux I__4663 (
            .O(N__21076),
            .I(\uu2.bitmapZ0Z_314 ));
    LocalMux I__4662 (
            .O(N__21073),
            .I(\uu2.bitmapZ0Z_314 ));
    LocalMux I__4661 (
            .O(N__21070),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__4660 (
            .O(N__21063),
            .I(N__21060));
    LocalMux I__4659 (
            .O(N__21060),
            .I(\uu2.bitmap_RNI020QZ0Z_186 ));
    InMux I__4658 (
            .O(N__21057),
            .I(N__21054));
    LocalMux I__4657 (
            .O(N__21054),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__4656 (
            .O(N__21051),
            .I(N__21044));
    InMux I__4655 (
            .O(N__21050),
            .I(N__21044));
    CascadeMux I__4654 (
            .O(N__21049),
            .I(N__21041));
    LocalMux I__4653 (
            .O(N__21044),
            .I(N__21038));
    InMux I__4652 (
            .O(N__21041),
            .I(N__21034));
    Span4Mux_h I__4651 (
            .O(N__21038),
            .I(N__21031));
    InMux I__4650 (
            .O(N__21037),
            .I(N__21028));
    LocalMux I__4649 (
            .O(N__21034),
            .I(N__21025));
    Span4Mux_h I__4648 (
            .O(N__21031),
            .I(N__21022));
    LocalMux I__4647 (
            .O(N__21028),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv12 I__4646 (
            .O(N__21025),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__4645 (
            .O(N__21022),
            .I(\uu2.w_addr_userZ0Z_5 ));
    InMux I__4644 (
            .O(N__21015),
            .I(N__21009));
    InMux I__4643 (
            .O(N__21014),
            .I(N__21006));
    InMux I__4642 (
            .O(N__21013),
            .I(N__21003));
    CascadeMux I__4641 (
            .O(N__21012),
            .I(N__21000));
    LocalMux I__4640 (
            .O(N__21009),
            .I(N__20996));
    LocalMux I__4639 (
            .O(N__21006),
            .I(N__20991));
    LocalMux I__4638 (
            .O(N__21003),
            .I(N__20991));
    InMux I__4637 (
            .O(N__21000),
            .I(N__20986));
    InMux I__4636 (
            .O(N__20999),
            .I(N__20986));
    Span4Mux_s0_v I__4635 (
            .O(N__20996),
            .I(N__20983));
    Span12Mux_s10_h I__4634 (
            .O(N__20991),
            .I(N__20980));
    LocalMux I__4633 (
            .O(N__20986),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__4632 (
            .O(N__20983),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv12 I__4631 (
            .O(N__20980),
            .I(\uu2.w_addr_userZ0Z_4 ));
    InMux I__4630 (
            .O(N__20973),
            .I(N__20964));
    InMux I__4629 (
            .O(N__20972),
            .I(N__20964));
    InMux I__4628 (
            .O(N__20971),
            .I(N__20964));
    LocalMux I__4627 (
            .O(N__20964),
            .I(N__20961));
    Span4Mux_s1_h I__4626 (
            .O(N__20961),
            .I(N__20955));
    InMux I__4625 (
            .O(N__20960),
            .I(N__20948));
    InMux I__4624 (
            .O(N__20959),
            .I(N__20948));
    InMux I__4623 (
            .O(N__20958),
            .I(N__20948));
    Span4Mux_h I__4622 (
            .O(N__20955),
            .I(N__20944));
    LocalMux I__4621 (
            .O(N__20948),
            .I(N__20941));
    InMux I__4620 (
            .O(N__20947),
            .I(N__20938));
    Odrv4 I__4619 (
            .O(N__20944),
            .I(\uu2.un28_w_addr_user_i ));
    Odrv4 I__4618 (
            .O(N__20941),
            .I(\uu2.un28_w_addr_user_i ));
    LocalMux I__4617 (
            .O(N__20938),
            .I(\uu2.un28_w_addr_user_i ));
    InMux I__4616 (
            .O(N__20931),
            .I(N__20922));
    InMux I__4615 (
            .O(N__20930),
            .I(N__20922));
    InMux I__4614 (
            .O(N__20929),
            .I(N__20922));
    LocalMux I__4613 (
            .O(N__20922),
            .I(N__20917));
    InMux I__4612 (
            .O(N__20921),
            .I(N__20912));
    InMux I__4611 (
            .O(N__20920),
            .I(N__20912));
    Odrv12 I__4610 (
            .O(N__20917),
            .I(\uu2.un404_ci ));
    LocalMux I__4609 (
            .O(N__20912),
            .I(\uu2.un404_ci ));
    CascadeMux I__4608 (
            .O(N__20907),
            .I(N__20904));
    InMux I__4607 (
            .O(N__20904),
            .I(N__20901));
    LocalMux I__4606 (
            .O(N__20901),
            .I(N__20898));
    Span4Mux_s1_v I__4605 (
            .O(N__20898),
            .I(N__20895));
    Span4Mux_h I__4604 (
            .O(N__20895),
            .I(N__20891));
    InMux I__4603 (
            .O(N__20894),
            .I(N__20888));
    Odrv4 I__4602 (
            .O(N__20891),
            .I(\uu2.un426_ci_3 ));
    LocalMux I__4601 (
            .O(N__20888),
            .I(\uu2.un426_ci_3 ));
    InMux I__4600 (
            .O(N__20883),
            .I(N__20876));
    InMux I__4599 (
            .O(N__20882),
            .I(N__20876));
    CascadeMux I__4598 (
            .O(N__20881),
            .I(N__20873));
    LocalMux I__4597 (
            .O(N__20876),
            .I(N__20868));
    InMux I__4596 (
            .O(N__20873),
            .I(N__20865));
    InMux I__4595 (
            .O(N__20872),
            .I(N__20862));
    InMux I__4594 (
            .O(N__20871),
            .I(N__20859));
    Span12Mux_v I__4593 (
            .O(N__20868),
            .I(N__20854));
    LocalMux I__4592 (
            .O(N__20865),
            .I(N__20854));
    LocalMux I__4591 (
            .O(N__20862),
            .I(N__20851));
    LocalMux I__4590 (
            .O(N__20859),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv12 I__4589 (
            .O(N__20854),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__4588 (
            .O(N__20851),
            .I(\uu2.w_addr_userZ0Z_6 ));
    SRMux I__4587 (
            .O(N__20844),
            .I(N__20839));
    SRMux I__4586 (
            .O(N__20843),
            .I(N__20836));
    SRMux I__4585 (
            .O(N__20842),
            .I(N__20833));
    LocalMux I__4584 (
            .O(N__20839),
            .I(N__20830));
    LocalMux I__4583 (
            .O(N__20836),
            .I(N__20827));
    LocalMux I__4582 (
            .O(N__20833),
            .I(N__20824));
    Span12Mux_s2_v I__4581 (
            .O(N__20830),
            .I(N__20820));
    Span4Mux_s2_v I__4580 (
            .O(N__20827),
            .I(N__20817));
    Span4Mux_h I__4579 (
            .O(N__20824),
            .I(N__20814));
    InMux I__4578 (
            .O(N__20823),
            .I(N__20811));
    Odrv12 I__4577 (
            .O(N__20820),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    Odrv4 I__4576 (
            .O(N__20817),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    Odrv4 I__4575 (
            .O(N__20814),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    LocalMux I__4574 (
            .O(N__20811),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_2 ));
    CascadeMux I__4573 (
            .O(N__20802),
            .I(\uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_ ));
    InMux I__4572 (
            .O(N__20799),
            .I(N__20796));
    LocalMux I__4571 (
            .O(N__20796),
            .I(N__20793));
    Odrv12 I__4570 (
            .O(N__20793),
            .I(\uu2.N_397 ));
    InMux I__4569 (
            .O(N__20790),
            .I(N__20785));
    InMux I__4568 (
            .O(N__20789),
            .I(N__20778));
    InMux I__4567 (
            .O(N__20788),
            .I(N__20778));
    LocalMux I__4566 (
            .O(N__20785),
            .I(N__20775));
    InMux I__4565 (
            .O(N__20784),
            .I(N__20770));
    InMux I__4564 (
            .O(N__20783),
            .I(N__20770));
    LocalMux I__4563 (
            .O(N__20778),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    Odrv4 I__4562 (
            .O(N__20775),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    LocalMux I__4561 (
            .O(N__20770),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    InMux I__4560 (
            .O(N__20763),
            .I(N__20745));
    InMux I__4559 (
            .O(N__20762),
            .I(N__20745));
    InMux I__4558 (
            .O(N__20761),
            .I(N__20745));
    InMux I__4557 (
            .O(N__20760),
            .I(N__20745));
    InMux I__4556 (
            .O(N__20759),
            .I(N__20737));
    InMux I__4555 (
            .O(N__20758),
            .I(N__20737));
    InMux I__4554 (
            .O(N__20757),
            .I(N__20734));
    InMux I__4553 (
            .O(N__20756),
            .I(N__20731));
    InMux I__4552 (
            .O(N__20755),
            .I(N__20728));
    InMux I__4551 (
            .O(N__20754),
            .I(N__20725));
    LocalMux I__4550 (
            .O(N__20745),
            .I(N__20722));
    InMux I__4549 (
            .O(N__20744),
            .I(N__20717));
    InMux I__4548 (
            .O(N__20743),
            .I(N__20717));
    InMux I__4547 (
            .O(N__20742),
            .I(N__20714));
    LocalMux I__4546 (
            .O(N__20737),
            .I(N__20711));
    LocalMux I__4545 (
            .O(N__20734),
            .I(N__20706));
    LocalMux I__4544 (
            .O(N__20731),
            .I(N__20706));
    LocalMux I__4543 (
            .O(N__20728),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    LocalMux I__4542 (
            .O(N__20725),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    Odrv4 I__4541 (
            .O(N__20722),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    LocalMux I__4540 (
            .O(N__20717),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    LocalMux I__4539 (
            .O(N__20714),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    Odrv4 I__4538 (
            .O(N__20711),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    Odrv4 I__4537 (
            .O(N__20706),
            .I(\uu2.w_addr_displayingZ1Z_3 ));
    InMux I__4536 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__4535 (
            .O(N__20688),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    CascadeMux I__4534 (
            .O(N__20685),
            .I(N__20682));
    InMux I__4533 (
            .O(N__20682),
            .I(N__20679));
    LocalMux I__4532 (
            .O(N__20679),
            .I(\uu2.N_32 ));
    InMux I__4531 (
            .O(N__20676),
            .I(N__20669));
    InMux I__4530 (
            .O(N__20675),
            .I(N__20664));
    InMux I__4529 (
            .O(N__20674),
            .I(N__20664));
    InMux I__4528 (
            .O(N__20673),
            .I(N__20656));
    InMux I__4527 (
            .O(N__20672),
            .I(N__20656));
    LocalMux I__4526 (
            .O(N__20669),
            .I(N__20653));
    LocalMux I__4525 (
            .O(N__20664),
            .I(N__20650));
    InMux I__4524 (
            .O(N__20663),
            .I(N__20643));
    InMux I__4523 (
            .O(N__20662),
            .I(N__20643));
    InMux I__4522 (
            .O(N__20661),
            .I(N__20643));
    LocalMux I__4521 (
            .O(N__20656),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__4520 (
            .O(N__20653),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv12 I__4519 (
            .O(N__20650),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__4518 (
            .O(N__20643),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__4517 (
            .O(N__20634),
            .I(N__20630));
    InMux I__4516 (
            .O(N__20633),
            .I(N__20625));
    LocalMux I__4515 (
            .O(N__20630),
            .I(N__20622));
    InMux I__4514 (
            .O(N__20629),
            .I(N__20617));
    InMux I__4513 (
            .O(N__20628),
            .I(N__20617));
    LocalMux I__4512 (
            .O(N__20625),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__4511 (
            .O(N__20622),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__4510 (
            .O(N__20617),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__4509 (
            .O(N__20610),
            .I(N__20607));
    LocalMux I__4508 (
            .O(N__20607),
            .I(N__20604));
    Odrv4 I__4507 (
            .O(N__20604),
            .I(\uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2 ));
    CascadeMux I__4506 (
            .O(N__20601),
            .I(N__20598));
    InMux I__4505 (
            .O(N__20598),
            .I(N__20586));
    InMux I__4504 (
            .O(N__20597),
            .I(N__20586));
    InMux I__4503 (
            .O(N__20596),
            .I(N__20581));
    InMux I__4502 (
            .O(N__20595),
            .I(N__20581));
    InMux I__4501 (
            .O(N__20594),
            .I(N__20567));
    InMux I__4500 (
            .O(N__20593),
            .I(N__20567));
    InMux I__4499 (
            .O(N__20592),
            .I(N__20567));
    InMux I__4498 (
            .O(N__20591),
            .I(N__20567));
    LocalMux I__4497 (
            .O(N__20586),
            .I(N__20562));
    LocalMux I__4496 (
            .O(N__20581),
            .I(N__20562));
    InMux I__4495 (
            .O(N__20580),
            .I(N__20555));
    InMux I__4494 (
            .O(N__20579),
            .I(N__20555));
    InMux I__4493 (
            .O(N__20578),
            .I(N__20555));
    InMux I__4492 (
            .O(N__20577),
            .I(N__20552));
    InMux I__4491 (
            .O(N__20576),
            .I(N__20549));
    LocalMux I__4490 (
            .O(N__20567),
            .I(N__20546));
    Span4Mux_v I__4489 (
            .O(N__20562),
            .I(N__20541));
    LocalMux I__4488 (
            .O(N__20555),
            .I(N__20541));
    LocalMux I__4487 (
            .O(N__20552),
            .I(\Lab_UT.dictrl.m23_aZ0Z0 ));
    LocalMux I__4486 (
            .O(N__20549),
            .I(\Lab_UT.dictrl.m23_aZ0Z0 ));
    Odrv12 I__4485 (
            .O(N__20546),
            .I(\Lab_UT.dictrl.m23_aZ0Z0 ));
    Odrv4 I__4484 (
            .O(N__20541),
            .I(\Lab_UT.dictrl.m23_aZ0Z0 ));
    InMux I__4483 (
            .O(N__20532),
            .I(N__20529));
    LocalMux I__4482 (
            .O(N__20529),
            .I(\Lab_UT.dictrl.N_40_7 ));
    CascadeMux I__4481 (
            .O(N__20526),
            .I(\Lab_UT.dictrl.N_40_7_cascade_ ));
    InMux I__4480 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__4479 (
            .O(N__20520),
            .I(\Lab_UT.dictrl.g2_1_5 ));
    CascadeMux I__4478 (
            .O(N__20517),
            .I(\Lab_UT.dictrl.N_1462_5_cascade_ ));
    InMux I__4477 (
            .O(N__20514),
            .I(N__20511));
    LocalMux I__4476 (
            .O(N__20511),
            .I(\Lab_UT.dictrl.N_1102_5 ));
    InMux I__4475 (
            .O(N__20508),
            .I(N__20505));
    LocalMux I__4474 (
            .O(N__20505),
            .I(N__20499));
    InMux I__4473 (
            .O(N__20504),
            .I(N__20494));
    CascadeMux I__4472 (
            .O(N__20503),
            .I(N__20490));
    InMux I__4471 (
            .O(N__20502),
            .I(N__20484));
    Span4Mux_v I__4470 (
            .O(N__20499),
            .I(N__20481));
    InMux I__4469 (
            .O(N__20498),
            .I(N__20476));
    InMux I__4468 (
            .O(N__20497),
            .I(N__20476));
    LocalMux I__4467 (
            .O(N__20494),
            .I(N__20473));
    InMux I__4466 (
            .O(N__20493),
            .I(N__20470));
    InMux I__4465 (
            .O(N__20490),
            .I(N__20465));
    InMux I__4464 (
            .O(N__20489),
            .I(N__20465));
    CascadeMux I__4463 (
            .O(N__20488),
            .I(N__20462));
    InMux I__4462 (
            .O(N__20487),
            .I(N__20459));
    LocalMux I__4461 (
            .O(N__20484),
            .I(N__20456));
    Sp12to4 I__4460 (
            .O(N__20481),
            .I(N__20453));
    LocalMux I__4459 (
            .O(N__20476),
            .I(N__20450));
    Span4Mux_h I__4458 (
            .O(N__20473),
            .I(N__20445));
    LocalMux I__4457 (
            .O(N__20470),
            .I(N__20445));
    LocalMux I__4456 (
            .O(N__20465),
            .I(N__20442));
    InMux I__4455 (
            .O(N__20462),
            .I(N__20439));
    LocalMux I__4454 (
            .O(N__20459),
            .I(N__20436));
    Span4Mux_v I__4453 (
            .O(N__20456),
            .I(N__20433));
    Span12Mux_s8_h I__4452 (
            .O(N__20453),
            .I(N__20430));
    Span4Mux_h I__4451 (
            .O(N__20450),
            .I(N__20423));
    Span4Mux_h I__4450 (
            .O(N__20445),
            .I(N__20423));
    Span4Mux_s3_h I__4449 (
            .O(N__20442),
            .I(N__20423));
    LocalMux I__4448 (
            .O(N__20439),
            .I(N__20418));
    Span4Mux_h I__4447 (
            .O(N__20436),
            .I(N__20418));
    Odrv4 I__4446 (
            .O(N__20433),
            .I(bu_rx_data_0_rep1));
    Odrv12 I__4445 (
            .O(N__20430),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__4444 (
            .O(N__20423),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__4443 (
            .O(N__20418),
            .I(bu_rx_data_0_rep1));
    CascadeMux I__4442 (
            .O(N__20409),
            .I(N__20403));
    InMux I__4441 (
            .O(N__20408),
            .I(N__20399));
    CascadeMux I__4440 (
            .O(N__20407),
            .I(N__20396));
    InMux I__4439 (
            .O(N__20406),
            .I(N__20387));
    InMux I__4438 (
            .O(N__20403),
            .I(N__20387));
    InMux I__4437 (
            .O(N__20402),
            .I(N__20387));
    LocalMux I__4436 (
            .O(N__20399),
            .I(N__20384));
    InMux I__4435 (
            .O(N__20396),
            .I(N__20379));
    InMux I__4434 (
            .O(N__20395),
            .I(N__20379));
    InMux I__4433 (
            .O(N__20394),
            .I(N__20376));
    LocalMux I__4432 (
            .O(N__20387),
            .I(N__20372));
    Span4Mux_s2_v I__4431 (
            .O(N__20384),
            .I(N__20367));
    LocalMux I__4430 (
            .O(N__20379),
            .I(N__20367));
    LocalMux I__4429 (
            .O(N__20376),
            .I(N__20364));
    CascadeMux I__4428 (
            .O(N__20375),
            .I(N__20361));
    Span4Mux_s2_v I__4427 (
            .O(N__20372),
            .I(N__20357));
    Span4Mux_v I__4426 (
            .O(N__20367),
            .I(N__20354));
    Span4Mux_s2_v I__4425 (
            .O(N__20364),
            .I(N__20351));
    InMux I__4424 (
            .O(N__20361),
            .I(N__20348));
    InMux I__4423 (
            .O(N__20360),
            .I(N__20345));
    Span4Mux_v I__4422 (
            .O(N__20357),
            .I(N__20342));
    Span4Mux_h I__4421 (
            .O(N__20354),
            .I(N__20337));
    Span4Mux_v I__4420 (
            .O(N__20351),
            .I(N__20337));
    LocalMux I__4419 (
            .O(N__20348),
            .I(N__20332));
    LocalMux I__4418 (
            .O(N__20345),
            .I(N__20332));
    Odrv4 I__4417 (
            .O(N__20342),
            .I(bu_rx_data_5_rep1));
    Odrv4 I__4416 (
            .O(N__20337),
            .I(bu_rx_data_5_rep1));
    Odrv12 I__4415 (
            .O(N__20332),
            .I(bu_rx_data_5_rep1));
    InMux I__4414 (
            .O(N__20325),
            .I(N__20311));
    InMux I__4413 (
            .O(N__20324),
            .I(N__20311));
    InMux I__4412 (
            .O(N__20323),
            .I(N__20311));
    InMux I__4411 (
            .O(N__20322),
            .I(N__20301));
    InMux I__4410 (
            .O(N__20321),
            .I(N__20301));
    InMux I__4409 (
            .O(N__20320),
            .I(N__20301));
    InMux I__4408 (
            .O(N__20319),
            .I(N__20301));
    InMux I__4407 (
            .O(N__20318),
            .I(N__20298));
    LocalMux I__4406 (
            .O(N__20311),
            .I(N__20292));
    InMux I__4405 (
            .O(N__20310),
            .I(N__20289));
    LocalMux I__4404 (
            .O(N__20301),
            .I(N__20284));
    LocalMux I__4403 (
            .O(N__20298),
            .I(N__20284));
    InMux I__4402 (
            .O(N__20297),
            .I(N__20279));
    InMux I__4401 (
            .O(N__20296),
            .I(N__20274));
    InMux I__4400 (
            .O(N__20295),
            .I(N__20274));
    Span4Mux_v I__4399 (
            .O(N__20292),
            .I(N__20269));
    LocalMux I__4398 (
            .O(N__20289),
            .I(N__20269));
    Span4Mux_s3_v I__4397 (
            .O(N__20284),
            .I(N__20264));
    InMux I__4396 (
            .O(N__20283),
            .I(N__20259));
    InMux I__4395 (
            .O(N__20282),
            .I(N__20259));
    LocalMux I__4394 (
            .O(N__20279),
            .I(N__20256));
    LocalMux I__4393 (
            .O(N__20274),
            .I(N__20251));
    Span4Mux_h I__4392 (
            .O(N__20269),
            .I(N__20251));
    InMux I__4391 (
            .O(N__20268),
            .I(N__20246));
    InMux I__4390 (
            .O(N__20267),
            .I(N__20246));
    Span4Mux_h I__4389 (
            .O(N__20264),
            .I(N__20241));
    LocalMux I__4388 (
            .O(N__20259),
            .I(N__20241));
    Odrv4 I__4387 (
            .O(N__20256),
            .I(bu_rx_data_4_rep2));
    Odrv4 I__4386 (
            .O(N__20251),
            .I(bu_rx_data_4_rep2));
    LocalMux I__4385 (
            .O(N__20246),
            .I(bu_rx_data_4_rep2));
    Odrv4 I__4384 (
            .O(N__20241),
            .I(bu_rx_data_4_rep2));
    InMux I__4383 (
            .O(N__20232),
            .I(N__20229));
    LocalMux I__4382 (
            .O(N__20229),
            .I(N__20226));
    Odrv4 I__4381 (
            .O(N__20226),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_4_8 ));
    CascadeMux I__4380 (
            .O(N__20223),
            .I(N__20211));
    CascadeMux I__4379 (
            .O(N__20222),
            .I(N__20208));
    CascadeMux I__4378 (
            .O(N__20221),
            .I(N__20202));
    CascadeMux I__4377 (
            .O(N__20220),
            .I(N__20199));
    InMux I__4376 (
            .O(N__20219),
            .I(N__20193));
    InMux I__4375 (
            .O(N__20218),
            .I(N__20186));
    InMux I__4374 (
            .O(N__20217),
            .I(N__20186));
    InMux I__4373 (
            .O(N__20216),
            .I(N__20183));
    InMux I__4372 (
            .O(N__20215),
            .I(N__20178));
    InMux I__4371 (
            .O(N__20214),
            .I(N__20178));
    InMux I__4370 (
            .O(N__20211),
            .I(N__20169));
    InMux I__4369 (
            .O(N__20208),
            .I(N__20169));
    InMux I__4368 (
            .O(N__20207),
            .I(N__20169));
    InMux I__4367 (
            .O(N__20206),
            .I(N__20169));
    InMux I__4366 (
            .O(N__20205),
            .I(N__20160));
    InMux I__4365 (
            .O(N__20202),
            .I(N__20160));
    InMux I__4364 (
            .O(N__20199),
            .I(N__20160));
    InMux I__4363 (
            .O(N__20198),
            .I(N__20160));
    InMux I__4362 (
            .O(N__20197),
            .I(N__20152));
    InMux I__4361 (
            .O(N__20196),
            .I(N__20152));
    LocalMux I__4360 (
            .O(N__20193),
            .I(N__20149));
    InMux I__4359 (
            .O(N__20192),
            .I(N__20144));
    InMux I__4358 (
            .O(N__20191),
            .I(N__20144));
    LocalMux I__4357 (
            .O(N__20186),
            .I(N__20140));
    LocalMux I__4356 (
            .O(N__20183),
            .I(N__20135));
    LocalMux I__4355 (
            .O(N__20178),
            .I(N__20135));
    LocalMux I__4354 (
            .O(N__20169),
            .I(N__20130));
    LocalMux I__4353 (
            .O(N__20160),
            .I(N__20130));
    InMux I__4352 (
            .O(N__20159),
            .I(N__20123));
    InMux I__4351 (
            .O(N__20158),
            .I(N__20123));
    InMux I__4350 (
            .O(N__20157),
            .I(N__20123));
    LocalMux I__4349 (
            .O(N__20152),
            .I(N__20116));
    Span4Mux_v I__4348 (
            .O(N__20149),
            .I(N__20116));
    LocalMux I__4347 (
            .O(N__20144),
            .I(N__20116));
    InMux I__4346 (
            .O(N__20143),
            .I(N__20113));
    Span4Mux_v I__4345 (
            .O(N__20140),
            .I(N__20104));
    Span4Mux_s2_v I__4344 (
            .O(N__20135),
            .I(N__20104));
    Span4Mux_h I__4343 (
            .O(N__20130),
            .I(N__20104));
    LocalMux I__4342 (
            .O(N__20123),
            .I(N__20104));
    Span4Mux_h I__4341 (
            .O(N__20116),
            .I(N__20099));
    LocalMux I__4340 (
            .O(N__20113),
            .I(N__20099));
    Odrv4 I__4339 (
            .O(N__20104),
            .I(\Lab_UT.dictrl.N_19_0 ));
    Odrv4 I__4338 (
            .O(N__20099),
            .I(\Lab_UT.dictrl.N_19_0 ));
    CascadeMux I__4337 (
            .O(N__20094),
            .I(N__20087));
    CascadeMux I__4336 (
            .O(N__20093),
            .I(N__20083));
    CascadeMux I__4335 (
            .O(N__20092),
            .I(N__20079));
    CascadeMux I__4334 (
            .O(N__20091),
            .I(N__20072));
    InMux I__4333 (
            .O(N__20090),
            .I(N__20067));
    InMux I__4332 (
            .O(N__20087),
            .I(N__20064));
    InMux I__4331 (
            .O(N__20086),
            .I(N__20055));
    InMux I__4330 (
            .O(N__20083),
            .I(N__20055));
    InMux I__4329 (
            .O(N__20082),
            .I(N__20055));
    InMux I__4328 (
            .O(N__20079),
            .I(N__20055));
    InMux I__4327 (
            .O(N__20078),
            .I(N__20050));
    InMux I__4326 (
            .O(N__20077),
            .I(N__20050));
    CascadeMux I__4325 (
            .O(N__20076),
            .I(N__20046));
    InMux I__4324 (
            .O(N__20075),
            .I(N__20040));
    InMux I__4323 (
            .O(N__20072),
            .I(N__20040));
    InMux I__4322 (
            .O(N__20071),
            .I(N__20035));
    InMux I__4321 (
            .O(N__20070),
            .I(N__20035));
    LocalMux I__4320 (
            .O(N__20067),
            .I(N__20032));
    LocalMux I__4319 (
            .O(N__20064),
            .I(N__20028));
    LocalMux I__4318 (
            .O(N__20055),
            .I(N__20023));
    LocalMux I__4317 (
            .O(N__20050),
            .I(N__20023));
    InMux I__4316 (
            .O(N__20049),
            .I(N__20018));
    InMux I__4315 (
            .O(N__20046),
            .I(N__20018));
    CascadeMux I__4314 (
            .O(N__20045),
            .I(N__20015));
    LocalMux I__4313 (
            .O(N__20040),
            .I(N__20012));
    LocalMux I__4312 (
            .O(N__20035),
            .I(N__20009));
    Span4Mux_s1_v I__4311 (
            .O(N__20032),
            .I(N__20006));
    InMux I__4310 (
            .O(N__20031),
            .I(N__20003));
    Span4Mux_h I__4309 (
            .O(N__20028),
            .I(N__19998));
    Span4Mux_h I__4308 (
            .O(N__20023),
            .I(N__19998));
    LocalMux I__4307 (
            .O(N__20018),
            .I(N__19995));
    InMux I__4306 (
            .O(N__20015),
            .I(N__19992));
    Span4Mux_v I__4305 (
            .O(N__20012),
            .I(N__19987));
    Span4Mux_h I__4304 (
            .O(N__20009),
            .I(N__19987));
    Sp12to4 I__4303 (
            .O(N__20006),
            .I(N__19982));
    LocalMux I__4302 (
            .O(N__20003),
            .I(N__19982));
    Span4Mux_h I__4301 (
            .O(N__19998),
            .I(N__19979));
    Span4Mux_h I__4300 (
            .O(N__19995),
            .I(N__19974));
    LocalMux I__4299 (
            .O(N__19992),
            .I(N__19974));
    Span4Mux_h I__4298 (
            .O(N__19987),
            .I(N__19971));
    Odrv12 I__4297 (
            .O(N__19982),
            .I(bu_rx_data_6_rep2));
    Odrv4 I__4296 (
            .O(N__19979),
            .I(bu_rx_data_6_rep2));
    Odrv4 I__4295 (
            .O(N__19974),
            .I(bu_rx_data_6_rep2));
    Odrv4 I__4294 (
            .O(N__19971),
            .I(bu_rx_data_6_rep2));
    InMux I__4293 (
            .O(N__19962),
            .I(N__19948));
    InMux I__4292 (
            .O(N__19961),
            .I(N__19945));
    InMux I__4291 (
            .O(N__19960),
            .I(N__19942));
    InMux I__4290 (
            .O(N__19959),
            .I(N__19939));
    InMux I__4289 (
            .O(N__19958),
            .I(N__19936));
    InMux I__4288 (
            .O(N__19957),
            .I(N__19933));
    InMux I__4287 (
            .O(N__19956),
            .I(N__19926));
    InMux I__4286 (
            .O(N__19955),
            .I(N__19926));
    InMux I__4285 (
            .O(N__19954),
            .I(N__19926));
    InMux I__4284 (
            .O(N__19953),
            .I(N__19921));
    InMux I__4283 (
            .O(N__19952),
            .I(N__19921));
    InMux I__4282 (
            .O(N__19951),
            .I(N__19918));
    LocalMux I__4281 (
            .O(N__19948),
            .I(N__19914));
    LocalMux I__4280 (
            .O(N__19945),
            .I(N__19909));
    LocalMux I__4279 (
            .O(N__19942),
            .I(N__19909));
    LocalMux I__4278 (
            .O(N__19939),
            .I(N__19904));
    LocalMux I__4277 (
            .O(N__19936),
            .I(N__19904));
    LocalMux I__4276 (
            .O(N__19933),
            .I(N__19901));
    LocalMux I__4275 (
            .O(N__19926),
            .I(N__19898));
    LocalMux I__4274 (
            .O(N__19921),
            .I(N__19893));
    LocalMux I__4273 (
            .O(N__19918),
            .I(N__19893));
    InMux I__4272 (
            .O(N__19917),
            .I(N__19890));
    Span12Mux_s2_v I__4271 (
            .O(N__19914),
            .I(N__19885));
    Span12Mux_v I__4270 (
            .O(N__19909),
            .I(N__19885));
    Span4Mux_v I__4269 (
            .O(N__19904),
            .I(N__19880));
    Span4Mux_s2_v I__4268 (
            .O(N__19901),
            .I(N__19880));
    Span4Mux_h I__4267 (
            .O(N__19898),
            .I(N__19875));
    Span4Mux_s2_v I__4266 (
            .O(N__19893),
            .I(N__19875));
    LocalMux I__4265 (
            .O(N__19890),
            .I(N__19872));
    Odrv12 I__4264 (
            .O(N__19885),
            .I(\Lab_UT.dictrl.m40Z0Z_1 ));
    Odrv4 I__4263 (
            .O(N__19880),
            .I(\Lab_UT.dictrl.m40Z0Z_1 ));
    Odrv4 I__4262 (
            .O(N__19875),
            .I(\Lab_UT.dictrl.m40Z0Z_1 ));
    Odrv12 I__4261 (
            .O(N__19872),
            .I(\Lab_UT.dictrl.m40Z0Z_1 ));
    InMux I__4260 (
            .O(N__19863),
            .I(N__19860));
    LocalMux I__4259 (
            .O(N__19860),
            .I(N__19857));
    Span4Mux_h I__4258 (
            .O(N__19857),
            .I(N__19854));
    Odrv4 I__4257 (
            .O(N__19854),
            .I(\Lab_UT.dictrl.m53_d_1_4 ));
    InMux I__4256 (
            .O(N__19851),
            .I(N__19845));
    InMux I__4255 (
            .O(N__19850),
            .I(N__19845));
    LocalMux I__4254 (
            .O(N__19845),
            .I(N__19840));
    InMux I__4253 (
            .O(N__19844),
            .I(N__19837));
    InMux I__4252 (
            .O(N__19843),
            .I(N__19834));
    Span4Mux_v I__4251 (
            .O(N__19840),
            .I(N__19825));
    LocalMux I__4250 (
            .O(N__19837),
            .I(N__19825));
    LocalMux I__4249 (
            .O(N__19834),
            .I(N__19816));
    InMux I__4248 (
            .O(N__19833),
            .I(N__19813));
    InMux I__4247 (
            .O(N__19832),
            .I(N__19810));
    InMux I__4246 (
            .O(N__19831),
            .I(N__19805));
    InMux I__4245 (
            .O(N__19830),
            .I(N__19805));
    Span4Mux_v I__4244 (
            .O(N__19825),
            .I(N__19802));
    InMux I__4243 (
            .O(N__19824),
            .I(N__19799));
    InMux I__4242 (
            .O(N__19823),
            .I(N__19788));
    InMux I__4241 (
            .O(N__19822),
            .I(N__19788));
    InMux I__4240 (
            .O(N__19821),
            .I(N__19788));
    InMux I__4239 (
            .O(N__19820),
            .I(N__19788));
    InMux I__4238 (
            .O(N__19819),
            .I(N__19788));
    Span4Mux_s3_v I__4237 (
            .O(N__19816),
            .I(N__19783));
    LocalMux I__4236 (
            .O(N__19813),
            .I(N__19783));
    LocalMux I__4235 (
            .O(N__19810),
            .I(N__19780));
    LocalMux I__4234 (
            .O(N__19805),
            .I(N__19775));
    Span4Mux_s0_v I__4233 (
            .O(N__19802),
            .I(N__19768));
    LocalMux I__4232 (
            .O(N__19799),
            .I(N__19768));
    LocalMux I__4231 (
            .O(N__19788),
            .I(N__19768));
    Span4Mux_v I__4230 (
            .O(N__19783),
            .I(N__19762));
    Span4Mux_v I__4229 (
            .O(N__19780),
            .I(N__19762));
    InMux I__4228 (
            .O(N__19779),
            .I(N__19757));
    InMux I__4227 (
            .O(N__19778),
            .I(N__19757));
    Span4Mux_v I__4226 (
            .O(N__19775),
            .I(N__19752));
    Span4Mux_v I__4225 (
            .O(N__19768),
            .I(N__19752));
    InMux I__4224 (
            .O(N__19767),
            .I(N__19749));
    Odrv4 I__4223 (
            .O(N__19762),
            .I(\Lab_UT.dictrl.state_2_rep2 ));
    LocalMux I__4222 (
            .O(N__19757),
            .I(\Lab_UT.dictrl.state_2_rep2 ));
    Odrv4 I__4221 (
            .O(N__19752),
            .I(\Lab_UT.dictrl.state_2_rep2 ));
    LocalMux I__4220 (
            .O(N__19749),
            .I(\Lab_UT.dictrl.state_2_rep2 ));
    CascadeMux I__4219 (
            .O(N__19740),
            .I(\Lab_UT.dictrl.N_97_mux_6_cascade_ ));
    CascadeMux I__4218 (
            .O(N__19737),
            .I(N__19731));
    CascadeMux I__4217 (
            .O(N__19736),
            .I(N__19726));
    InMux I__4216 (
            .O(N__19735),
            .I(N__19721));
    InMux I__4215 (
            .O(N__19734),
            .I(N__19717));
    InMux I__4214 (
            .O(N__19731),
            .I(N__19707));
    InMux I__4213 (
            .O(N__19730),
            .I(N__19704));
    InMux I__4212 (
            .O(N__19729),
            .I(N__19701));
    InMux I__4211 (
            .O(N__19726),
            .I(N__19697));
    InMux I__4210 (
            .O(N__19725),
            .I(N__19694));
    InMux I__4209 (
            .O(N__19724),
            .I(N__19691));
    LocalMux I__4208 (
            .O(N__19721),
            .I(N__19688));
    InMux I__4207 (
            .O(N__19720),
            .I(N__19685));
    LocalMux I__4206 (
            .O(N__19717),
            .I(N__19682));
    InMux I__4205 (
            .O(N__19716),
            .I(N__19679));
    InMux I__4204 (
            .O(N__19715),
            .I(N__19672));
    InMux I__4203 (
            .O(N__19714),
            .I(N__19672));
    InMux I__4202 (
            .O(N__19713),
            .I(N__19672));
    InMux I__4201 (
            .O(N__19712),
            .I(N__19667));
    InMux I__4200 (
            .O(N__19711),
            .I(N__19667));
    InMux I__4199 (
            .O(N__19710),
            .I(N__19662));
    LocalMux I__4198 (
            .O(N__19707),
            .I(N__19655));
    LocalMux I__4197 (
            .O(N__19704),
            .I(N__19655));
    LocalMux I__4196 (
            .O(N__19701),
            .I(N__19655));
    InMux I__4195 (
            .O(N__19700),
            .I(N__19652));
    LocalMux I__4194 (
            .O(N__19697),
            .I(N__19645));
    LocalMux I__4193 (
            .O(N__19694),
            .I(N__19645));
    LocalMux I__4192 (
            .O(N__19691),
            .I(N__19645));
    Span4Mux_s2_v I__4191 (
            .O(N__19688),
            .I(N__19642));
    LocalMux I__4190 (
            .O(N__19685),
            .I(N__19639));
    Span4Mux_s2_v I__4189 (
            .O(N__19682),
            .I(N__19632));
    LocalMux I__4188 (
            .O(N__19679),
            .I(N__19632));
    LocalMux I__4187 (
            .O(N__19672),
            .I(N__19632));
    LocalMux I__4186 (
            .O(N__19667),
            .I(N__19629));
    InMux I__4185 (
            .O(N__19666),
            .I(N__19624));
    InMux I__4184 (
            .O(N__19665),
            .I(N__19624));
    LocalMux I__4183 (
            .O(N__19662),
            .I(N__19619));
    Span4Mux_v I__4182 (
            .O(N__19655),
            .I(N__19619));
    LocalMux I__4181 (
            .O(N__19652),
            .I(N__19610));
    Span4Mux_s3_v I__4180 (
            .O(N__19645),
            .I(N__19610));
    Span4Mux_v I__4179 (
            .O(N__19642),
            .I(N__19607));
    Span4Mux_v I__4178 (
            .O(N__19639),
            .I(N__19596));
    Span4Mux_v I__4177 (
            .O(N__19632),
            .I(N__19596));
    Span4Mux_v I__4176 (
            .O(N__19629),
            .I(N__19596));
    LocalMux I__4175 (
            .O(N__19624),
            .I(N__19596));
    Span4Mux_h I__4174 (
            .O(N__19619),
            .I(N__19596));
    InMux I__4173 (
            .O(N__19618),
            .I(N__19593));
    InMux I__4172 (
            .O(N__19617),
            .I(N__19590));
    InMux I__4171 (
            .O(N__19616),
            .I(N__19585));
    InMux I__4170 (
            .O(N__19615),
            .I(N__19585));
    Odrv4 I__4169 (
            .O(N__19610),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv4 I__4168 (
            .O(N__19607),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv4 I__4167 (
            .O(N__19596),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    LocalMux I__4166 (
            .O(N__19593),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    LocalMux I__4165 (
            .O(N__19590),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    LocalMux I__4164 (
            .O(N__19585),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    InMux I__4163 (
            .O(N__19572),
            .I(N__19569));
    LocalMux I__4162 (
            .O(N__19569),
            .I(N__19566));
    Span4Mux_h I__4161 (
            .O(N__19566),
            .I(N__19563));
    Span4Mux_v I__4160 (
            .O(N__19563),
            .I(N__19560));
    Odrv4 I__4159 (
            .O(N__19560),
            .I(\Lab_UT.dictrl.g2_1_4 ));
    InMux I__4158 (
            .O(N__19557),
            .I(N__19554));
    LocalMux I__4157 (
            .O(N__19554),
            .I(\Lab_UT.dictrl.N_1462_4 ));
    CascadeMux I__4156 (
            .O(N__19551),
            .I(\Lab_UT.dictrl.N_1102_4_cascade_ ));
    InMux I__4155 (
            .O(N__19548),
            .I(N__19545));
    LocalMux I__4154 (
            .O(N__19545),
            .I(\Lab_UT.dictrl.N_6_0 ));
    CascadeMux I__4153 (
            .O(N__19542),
            .I(N__19539));
    InMux I__4152 (
            .O(N__19539),
            .I(N__19535));
    InMux I__4151 (
            .O(N__19538),
            .I(N__19529));
    LocalMux I__4150 (
            .O(N__19535),
            .I(N__19524));
    InMux I__4149 (
            .O(N__19534),
            .I(N__19519));
    InMux I__4148 (
            .O(N__19533),
            .I(N__19519));
    InMux I__4147 (
            .O(N__19532),
            .I(N__19516));
    LocalMux I__4146 (
            .O(N__19529),
            .I(N__19513));
    InMux I__4145 (
            .O(N__19528),
            .I(N__19510));
    CascadeMux I__4144 (
            .O(N__19527),
            .I(N__19507));
    Span4Mux_s2_v I__4143 (
            .O(N__19524),
            .I(N__19502));
    LocalMux I__4142 (
            .O(N__19519),
            .I(N__19502));
    LocalMux I__4141 (
            .O(N__19516),
            .I(N__19497));
    Span4Mux_s2_v I__4140 (
            .O(N__19513),
            .I(N__19497));
    LocalMux I__4139 (
            .O(N__19510),
            .I(N__19494));
    InMux I__4138 (
            .O(N__19507),
            .I(N__19491));
    Span4Mux_v I__4137 (
            .O(N__19502),
            .I(N__19488));
    Span4Mux_v I__4136 (
            .O(N__19497),
            .I(N__19485));
    Span4Mux_v I__4135 (
            .O(N__19494),
            .I(N__19478));
    LocalMux I__4134 (
            .O(N__19491),
            .I(N__19478));
    Span4Mux_s2_h I__4133 (
            .O(N__19488),
            .I(N__19478));
    Odrv4 I__4132 (
            .O(N__19485),
            .I(\Lab_UT.dictrl.next_state_2_1 ));
    Odrv4 I__4131 (
            .O(N__19478),
            .I(\Lab_UT.dictrl.next_state_2_1 ));
    InMux I__4130 (
            .O(N__19473),
            .I(N__19470));
    LocalMux I__4129 (
            .O(N__19470),
            .I(N__19467));
    Span4Mux_h I__4128 (
            .O(N__19467),
            .I(N__19464));
    Span4Mux_h I__4127 (
            .O(N__19464),
            .I(N__19461));
    Odrv4 I__4126 (
            .O(N__19461),
            .I(\Lab_UT.dictrl.g0_i_0 ));
    CascadeMux I__4125 (
            .O(N__19458),
            .I(N__19455));
    InMux I__4124 (
            .O(N__19455),
            .I(N__19452));
    LocalMux I__4123 (
            .O(N__19452),
            .I(\Lab_UT.dictrl.g1_1_1_0 ));
    InMux I__4122 (
            .O(N__19449),
            .I(N__19440));
    InMux I__4121 (
            .O(N__19448),
            .I(N__19440));
    InMux I__4120 (
            .O(N__19447),
            .I(N__19434));
    InMux I__4119 (
            .O(N__19446),
            .I(N__19434));
    InMux I__4118 (
            .O(N__19445),
            .I(N__19431));
    LocalMux I__4117 (
            .O(N__19440),
            .I(N__19428));
    InMux I__4116 (
            .O(N__19439),
            .I(N__19425));
    LocalMux I__4115 (
            .O(N__19434),
            .I(N__19418));
    LocalMux I__4114 (
            .O(N__19431),
            .I(N__19415));
    Span4Mux_v I__4113 (
            .O(N__19428),
            .I(N__19412));
    LocalMux I__4112 (
            .O(N__19425),
            .I(N__19409));
    InMux I__4111 (
            .O(N__19424),
            .I(N__19404));
    InMux I__4110 (
            .O(N__19423),
            .I(N__19404));
    InMux I__4109 (
            .O(N__19422),
            .I(N__19399));
    InMux I__4108 (
            .O(N__19421),
            .I(N__19399));
    Span12Mux_s10_h I__4107 (
            .O(N__19418),
            .I(N__19396));
    Span4Mux_v I__4106 (
            .O(N__19415),
            .I(N__19385));
    Span4Mux_h I__4105 (
            .O(N__19412),
            .I(N__19385));
    Span4Mux_v I__4104 (
            .O(N__19409),
            .I(N__19385));
    LocalMux I__4103 (
            .O(N__19404),
            .I(N__19385));
    LocalMux I__4102 (
            .O(N__19399),
            .I(N__19385));
    Odrv12 I__4101 (
            .O(N__19396),
            .I(bu_rx_data_7_rep1));
    Odrv4 I__4100 (
            .O(N__19385),
            .I(bu_rx_data_7_rep1));
    InMux I__4099 (
            .O(N__19380),
            .I(N__19377));
    LocalMux I__4098 (
            .O(N__19377),
            .I(N__19374));
    Span4Mux_h I__4097 (
            .O(N__19374),
            .I(N__19371));
    Odrv4 I__4096 (
            .O(N__19371),
            .I(\Lab_UT.dictrl.N_59 ));
    InMux I__4095 (
            .O(N__19368),
            .I(N__19363));
    InMux I__4094 (
            .O(N__19367),
            .I(N__19358));
    InMux I__4093 (
            .O(N__19366),
            .I(N__19358));
    LocalMux I__4092 (
            .O(N__19363),
            .I(N__19352));
    LocalMux I__4091 (
            .O(N__19358),
            .I(N__19352));
    InMux I__4090 (
            .O(N__19357),
            .I(N__19348));
    Span4Mux_v I__4089 (
            .O(N__19352),
            .I(N__19345));
    InMux I__4088 (
            .O(N__19351),
            .I(N__19342));
    LocalMux I__4087 (
            .O(N__19348),
            .I(\Lab_UT.dictrl.N_97_mux ));
    Odrv4 I__4086 (
            .O(N__19345),
            .I(\Lab_UT.dictrl.N_97_mux ));
    LocalMux I__4085 (
            .O(N__19342),
            .I(\Lab_UT.dictrl.N_97_mux ));
    CascadeMux I__4084 (
            .O(N__19335),
            .I(\Lab_UT.dictrl.N_59_cascade_ ));
    InMux I__4083 (
            .O(N__19332),
            .I(N__19321));
    InMux I__4082 (
            .O(N__19331),
            .I(N__19321));
    CascadeMux I__4081 (
            .O(N__19330),
            .I(N__19318));
    CascadeMux I__4080 (
            .O(N__19329),
            .I(N__19307));
    InMux I__4079 (
            .O(N__19328),
            .I(N__19298));
    InMux I__4078 (
            .O(N__19327),
            .I(N__19298));
    InMux I__4077 (
            .O(N__19326),
            .I(N__19298));
    LocalMux I__4076 (
            .O(N__19321),
            .I(N__19295));
    InMux I__4075 (
            .O(N__19318),
            .I(N__19290));
    InMux I__4074 (
            .O(N__19317),
            .I(N__19290));
    InMux I__4073 (
            .O(N__19316),
            .I(N__19285));
    InMux I__4072 (
            .O(N__19315),
            .I(N__19285));
    InMux I__4071 (
            .O(N__19314),
            .I(N__19280));
    InMux I__4070 (
            .O(N__19313),
            .I(N__19280));
    InMux I__4069 (
            .O(N__19312),
            .I(N__19275));
    InMux I__4068 (
            .O(N__19311),
            .I(N__19275));
    CascadeMux I__4067 (
            .O(N__19310),
            .I(N__19272));
    InMux I__4066 (
            .O(N__19307),
            .I(N__19264));
    InMux I__4065 (
            .O(N__19306),
            .I(N__19264));
    InMux I__4064 (
            .O(N__19305),
            .I(N__19264));
    LocalMux I__4063 (
            .O(N__19298),
            .I(N__19261));
    Span4Mux_h I__4062 (
            .O(N__19295),
            .I(N__19256));
    LocalMux I__4061 (
            .O(N__19290),
            .I(N__19256));
    LocalMux I__4060 (
            .O(N__19285),
            .I(N__19249));
    LocalMux I__4059 (
            .O(N__19280),
            .I(N__19249));
    LocalMux I__4058 (
            .O(N__19275),
            .I(N__19249));
    InMux I__4057 (
            .O(N__19272),
            .I(N__19246));
    InMux I__4056 (
            .O(N__19271),
            .I(N__19243));
    LocalMux I__4055 (
            .O(N__19264),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    Odrv4 I__4054 (
            .O(N__19261),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    Odrv4 I__4053 (
            .O(N__19256),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    Odrv12 I__4052 (
            .O(N__19249),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    LocalMux I__4051 (
            .O(N__19246),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    LocalMux I__4050 (
            .O(N__19243),
            .I(\Lab_UT.dictrl.state_0_rep2 ));
    CascadeMux I__4049 (
            .O(N__19230),
            .I(\Lab_UT.dictrl.N_40_5_cascade_ ));
    InMux I__4048 (
            .O(N__19227),
            .I(N__19223));
    InMux I__4047 (
            .O(N__19226),
            .I(N__19220));
    LocalMux I__4046 (
            .O(N__19223),
            .I(\Lab_UT.dictrl.N_40_4 ));
    LocalMux I__4045 (
            .O(N__19220),
            .I(\Lab_UT.dictrl.N_40_4 ));
    CascadeMux I__4044 (
            .O(N__19215),
            .I(\Lab_UT.dictrl.N_40_2_cascade_ ));
    InMux I__4043 (
            .O(N__19212),
            .I(N__19205));
    CascadeMux I__4042 (
            .O(N__19211),
            .I(N__19200));
    CascadeMux I__4041 (
            .O(N__19210),
            .I(N__19194));
    InMux I__4040 (
            .O(N__19209),
            .I(N__19185));
    InMux I__4039 (
            .O(N__19208),
            .I(N__19185));
    LocalMux I__4038 (
            .O(N__19205),
            .I(N__19182));
    InMux I__4037 (
            .O(N__19204),
            .I(N__19177));
    InMux I__4036 (
            .O(N__19203),
            .I(N__19177));
    InMux I__4035 (
            .O(N__19200),
            .I(N__19172));
    InMux I__4034 (
            .O(N__19199),
            .I(N__19172));
    InMux I__4033 (
            .O(N__19198),
            .I(N__19165));
    InMux I__4032 (
            .O(N__19197),
            .I(N__19165));
    InMux I__4031 (
            .O(N__19194),
            .I(N__19165));
    CascadeMux I__4030 (
            .O(N__19193),
            .I(N__19161));
    CascadeMux I__4029 (
            .O(N__19192),
            .I(N__19158));
    InMux I__4028 (
            .O(N__19191),
            .I(N__19154));
    CascadeMux I__4027 (
            .O(N__19190),
            .I(N__19151));
    LocalMux I__4026 (
            .O(N__19185),
            .I(N__19146));
    Span4Mux_s3_h I__4025 (
            .O(N__19182),
            .I(N__19143));
    LocalMux I__4024 (
            .O(N__19177),
            .I(N__19140));
    LocalMux I__4023 (
            .O(N__19172),
            .I(N__19137));
    LocalMux I__4022 (
            .O(N__19165),
            .I(N__19134));
    InMux I__4021 (
            .O(N__19164),
            .I(N__19129));
    InMux I__4020 (
            .O(N__19161),
            .I(N__19129));
    InMux I__4019 (
            .O(N__19158),
            .I(N__19124));
    InMux I__4018 (
            .O(N__19157),
            .I(N__19124));
    LocalMux I__4017 (
            .O(N__19154),
            .I(N__19121));
    InMux I__4016 (
            .O(N__19151),
            .I(N__19118));
    CascadeMux I__4015 (
            .O(N__19150),
            .I(N__19112));
    InMux I__4014 (
            .O(N__19149),
            .I(N__19109));
    Span4Mux_s3_h I__4013 (
            .O(N__19146),
            .I(N__19106));
    Sp12to4 I__4012 (
            .O(N__19143),
            .I(N__19101));
    Span12Mux_s8_h I__4011 (
            .O(N__19140),
            .I(N__19101));
    Span4Mux_v I__4010 (
            .O(N__19137),
            .I(N__19094));
    Span4Mux_v I__4009 (
            .O(N__19134),
            .I(N__19094));
    LocalMux I__4008 (
            .O(N__19129),
            .I(N__19094));
    LocalMux I__4007 (
            .O(N__19124),
            .I(N__19091));
    Span4Mux_s3_h I__4006 (
            .O(N__19121),
            .I(N__19088));
    LocalMux I__4005 (
            .O(N__19118),
            .I(N__19085));
    InMux I__4004 (
            .O(N__19117),
            .I(N__19076));
    InMux I__4003 (
            .O(N__19116),
            .I(N__19076));
    InMux I__4002 (
            .O(N__19115),
            .I(N__19076));
    InMux I__4001 (
            .O(N__19112),
            .I(N__19076));
    LocalMux I__4000 (
            .O(N__19109),
            .I(bu_rx_data_6));
    Odrv4 I__3999 (
            .O(N__19106),
            .I(bu_rx_data_6));
    Odrv12 I__3998 (
            .O(N__19101),
            .I(bu_rx_data_6));
    Odrv4 I__3997 (
            .O(N__19094),
            .I(bu_rx_data_6));
    Odrv4 I__3996 (
            .O(N__19091),
            .I(bu_rx_data_6));
    Odrv4 I__3995 (
            .O(N__19088),
            .I(bu_rx_data_6));
    Odrv12 I__3994 (
            .O(N__19085),
            .I(bu_rx_data_6));
    LocalMux I__3993 (
            .O(N__19076),
            .I(bu_rx_data_6));
    InMux I__3992 (
            .O(N__19059),
            .I(N__19056));
    LocalMux I__3991 (
            .O(N__19056),
            .I(\Lab_UT.dictrl.g0_i_a4_1_5 ));
    CascadeMux I__3990 (
            .O(N__19053),
            .I(\Lab_UT.dictrl.g0_i_a4_1_4_cascade_ ));
    InMux I__3989 (
            .O(N__19050),
            .I(N__19042));
    InMux I__3988 (
            .O(N__19049),
            .I(N__19042));
    CascadeMux I__3987 (
            .O(N__19048),
            .I(N__19037));
    InMux I__3986 (
            .O(N__19047),
            .I(N__19033));
    LocalMux I__3985 (
            .O(N__19042),
            .I(N__19030));
    InMux I__3984 (
            .O(N__19041),
            .I(N__19023));
    InMux I__3983 (
            .O(N__19040),
            .I(N__19023));
    InMux I__3982 (
            .O(N__19037),
            .I(N__19023));
    InMux I__3981 (
            .O(N__19036),
            .I(N__19020));
    LocalMux I__3980 (
            .O(N__19033),
            .I(N__19014));
    Span4Mux_v I__3979 (
            .O(N__19030),
            .I(N__19009));
    LocalMux I__3978 (
            .O(N__19023),
            .I(N__19009));
    LocalMux I__3977 (
            .O(N__19020),
            .I(N__19006));
    InMux I__3976 (
            .O(N__19019),
            .I(N__18999));
    InMux I__3975 (
            .O(N__19018),
            .I(N__18999));
    InMux I__3974 (
            .O(N__19017),
            .I(N__18999));
    Span12Mux_s3_h I__3973 (
            .O(N__19014),
            .I(N__18991));
    Span4Mux_h I__3972 (
            .O(N__19009),
            .I(N__18988));
    Span4Mux_s3_h I__3971 (
            .O(N__19006),
            .I(N__18985));
    LocalMux I__3970 (
            .O(N__18999),
            .I(N__18982));
    InMux I__3969 (
            .O(N__18998),
            .I(N__18971));
    InMux I__3968 (
            .O(N__18997),
            .I(N__18971));
    InMux I__3967 (
            .O(N__18996),
            .I(N__18971));
    InMux I__3966 (
            .O(N__18995),
            .I(N__18971));
    InMux I__3965 (
            .O(N__18994),
            .I(N__18971));
    Odrv12 I__3964 (
            .O(N__18991),
            .I(bu_rx_data_5));
    Odrv4 I__3963 (
            .O(N__18988),
            .I(bu_rx_data_5));
    Odrv4 I__3962 (
            .O(N__18985),
            .I(bu_rx_data_5));
    Odrv12 I__3961 (
            .O(N__18982),
            .I(bu_rx_data_5));
    LocalMux I__3960 (
            .O(N__18971),
            .I(bu_rx_data_5));
    InMux I__3959 (
            .O(N__18960),
            .I(N__18957));
    LocalMux I__3958 (
            .O(N__18957),
            .I(N__18954));
    Span4Mux_h I__3957 (
            .O(N__18954),
            .I(N__18951));
    Odrv4 I__3956 (
            .O(N__18951),
            .I(\Lab_UT.dictrl.N_12 ));
    InMux I__3955 (
            .O(N__18948),
            .I(N__18945));
    LocalMux I__3954 (
            .O(N__18945),
            .I(N__18942));
    Odrv12 I__3953 (
            .O(N__18942),
            .I(\Lab_UT.dictrl.N_4 ));
    CascadeMux I__3952 (
            .O(N__18939),
            .I(N__18928));
    CascadeMux I__3951 (
            .O(N__18938),
            .I(N__18924));
    CascadeMux I__3950 (
            .O(N__18937),
            .I(N__18921));
    InMux I__3949 (
            .O(N__18936),
            .I(N__18914));
    InMux I__3948 (
            .O(N__18935),
            .I(N__18914));
    CascadeMux I__3947 (
            .O(N__18934),
            .I(N__18911));
    InMux I__3946 (
            .O(N__18933),
            .I(N__18906));
    InMux I__3945 (
            .O(N__18932),
            .I(N__18901));
    InMux I__3944 (
            .O(N__18931),
            .I(N__18901));
    InMux I__3943 (
            .O(N__18928),
            .I(N__18898));
    InMux I__3942 (
            .O(N__18927),
            .I(N__18893));
    InMux I__3941 (
            .O(N__18924),
            .I(N__18893));
    InMux I__3940 (
            .O(N__18921),
            .I(N__18886));
    InMux I__3939 (
            .O(N__18920),
            .I(N__18886));
    CascadeMux I__3938 (
            .O(N__18919),
            .I(N__18883));
    LocalMux I__3937 (
            .O(N__18914),
            .I(N__18880));
    InMux I__3936 (
            .O(N__18911),
            .I(N__18877));
    InMux I__3935 (
            .O(N__18910),
            .I(N__18872));
    InMux I__3934 (
            .O(N__18909),
            .I(N__18869));
    LocalMux I__3933 (
            .O(N__18906),
            .I(N__18864));
    LocalMux I__3932 (
            .O(N__18901),
            .I(N__18864));
    LocalMux I__3931 (
            .O(N__18898),
            .I(N__18861));
    LocalMux I__3930 (
            .O(N__18893),
            .I(N__18858));
    CascadeMux I__3929 (
            .O(N__18892),
            .I(N__18855));
    InMux I__3928 (
            .O(N__18891),
            .I(N__18850));
    LocalMux I__3927 (
            .O(N__18886),
            .I(N__18847));
    InMux I__3926 (
            .O(N__18883),
            .I(N__18844));
    Span4Mux_v I__3925 (
            .O(N__18880),
            .I(N__18839));
    LocalMux I__3924 (
            .O(N__18877),
            .I(N__18839));
    InMux I__3923 (
            .O(N__18876),
            .I(N__18834));
    InMux I__3922 (
            .O(N__18875),
            .I(N__18834));
    LocalMux I__3921 (
            .O(N__18872),
            .I(N__18831));
    LocalMux I__3920 (
            .O(N__18869),
            .I(N__18822));
    Span4Mux_v I__3919 (
            .O(N__18864),
            .I(N__18822));
    Span4Mux_v I__3918 (
            .O(N__18861),
            .I(N__18822));
    Span4Mux_v I__3917 (
            .O(N__18858),
            .I(N__18822));
    InMux I__3916 (
            .O(N__18855),
            .I(N__18817));
    InMux I__3915 (
            .O(N__18854),
            .I(N__18817));
    InMux I__3914 (
            .O(N__18853),
            .I(N__18814));
    LocalMux I__3913 (
            .O(N__18850),
            .I(N__18811));
    Span4Mux_v I__3912 (
            .O(N__18847),
            .I(N__18804));
    LocalMux I__3911 (
            .O(N__18844),
            .I(N__18804));
    Span4Mux_h I__3910 (
            .O(N__18839),
            .I(N__18804));
    LocalMux I__3909 (
            .O(N__18834),
            .I(N__18797));
    Span4Mux_v I__3908 (
            .O(N__18831),
            .I(N__18797));
    Span4Mux_h I__3907 (
            .O(N__18822),
            .I(N__18797));
    LocalMux I__3906 (
            .O(N__18817),
            .I(N__18792));
    LocalMux I__3905 (
            .O(N__18814),
            .I(N__18792));
    Span4Mux_h I__3904 (
            .O(N__18811),
            .I(N__18787));
    Span4Mux_h I__3903 (
            .O(N__18804),
            .I(N__18787));
    Odrv4 I__3902 (
            .O(N__18797),
            .I(bu_rx_data_4));
    Odrv12 I__3901 (
            .O(N__18792),
            .I(bu_rx_data_4));
    Odrv4 I__3900 (
            .O(N__18787),
            .I(bu_rx_data_4));
    InMux I__3899 (
            .O(N__18780),
            .I(N__18777));
    LocalMux I__3898 (
            .O(N__18777),
            .I(N__18774));
    Odrv4 I__3897 (
            .O(N__18774),
            .I(\Lab_UT.dictrl.N_7 ));
    CascadeMux I__3896 (
            .O(N__18771),
            .I(N__18768));
    InMux I__3895 (
            .O(N__18768),
            .I(N__18765));
    LocalMux I__3894 (
            .O(N__18765),
            .I(N__18760));
    InMux I__3893 (
            .O(N__18764),
            .I(N__18756));
    CascadeMux I__3892 (
            .O(N__18763),
            .I(N__18753));
    Span4Mux_v I__3891 (
            .O(N__18760),
            .I(N__18747));
    InMux I__3890 (
            .O(N__18759),
            .I(N__18744));
    LocalMux I__3889 (
            .O(N__18756),
            .I(N__18741));
    InMux I__3888 (
            .O(N__18753),
            .I(N__18737));
    CascadeMux I__3887 (
            .O(N__18752),
            .I(N__18734));
    CascadeMux I__3886 (
            .O(N__18751),
            .I(N__18731));
    InMux I__3885 (
            .O(N__18750),
            .I(N__18726));
    Span4Mux_h I__3884 (
            .O(N__18747),
            .I(N__18719));
    LocalMux I__3883 (
            .O(N__18744),
            .I(N__18719));
    Span4Mux_h I__3882 (
            .O(N__18741),
            .I(N__18716));
    InMux I__3881 (
            .O(N__18740),
            .I(N__18713));
    LocalMux I__3880 (
            .O(N__18737),
            .I(N__18710));
    InMux I__3879 (
            .O(N__18734),
            .I(N__18701));
    InMux I__3878 (
            .O(N__18731),
            .I(N__18701));
    InMux I__3877 (
            .O(N__18730),
            .I(N__18701));
    InMux I__3876 (
            .O(N__18729),
            .I(N__18701));
    LocalMux I__3875 (
            .O(N__18726),
            .I(N__18698));
    CascadeMux I__3874 (
            .O(N__18725),
            .I(N__18695));
    CascadeMux I__3873 (
            .O(N__18724),
            .I(N__18692));
    Span4Mux_h I__3872 (
            .O(N__18719),
            .I(N__18689));
    Span4Mux_v I__3871 (
            .O(N__18716),
            .I(N__18686));
    LocalMux I__3870 (
            .O(N__18713),
            .I(N__18679));
    Span4Mux_v I__3869 (
            .O(N__18710),
            .I(N__18679));
    LocalMux I__3868 (
            .O(N__18701),
            .I(N__18679));
    Span4Mux_v I__3867 (
            .O(N__18698),
            .I(N__18676));
    InMux I__3866 (
            .O(N__18695),
            .I(N__18673));
    InMux I__3865 (
            .O(N__18692),
            .I(N__18670));
    Span4Mux_v I__3864 (
            .O(N__18689),
            .I(N__18665));
    Span4Mux_h I__3863 (
            .O(N__18686),
            .I(N__18665));
    Span4Mux_h I__3862 (
            .O(N__18679),
            .I(N__18662));
    Odrv4 I__3861 (
            .O(N__18676),
            .I(bu_rx_data_3_rep2));
    LocalMux I__3860 (
            .O(N__18673),
            .I(bu_rx_data_3_rep2));
    LocalMux I__3859 (
            .O(N__18670),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__3858 (
            .O(N__18665),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__3857 (
            .O(N__18662),
            .I(bu_rx_data_3_rep2));
    InMux I__3856 (
            .O(N__18651),
            .I(N__18646));
    InMux I__3855 (
            .O(N__18650),
            .I(N__18641));
    InMux I__3854 (
            .O(N__18649),
            .I(N__18641));
    LocalMux I__3853 (
            .O(N__18646),
            .I(N__18638));
    LocalMux I__3852 (
            .O(N__18641),
            .I(N__18635));
    Odrv12 I__3851 (
            .O(N__18638),
            .I(\Lab_UT.N_115 ));
    Odrv4 I__3850 (
            .O(N__18635),
            .I(\Lab_UT.N_115 ));
    InMux I__3849 (
            .O(N__18630),
            .I(N__18627));
    LocalMux I__3848 (
            .O(N__18627),
            .I(N__18622));
    InMux I__3847 (
            .O(N__18626),
            .I(N__18617));
    InMux I__3846 (
            .O(N__18625),
            .I(N__18617));
    Span4Mux_h I__3845 (
            .O(N__18622),
            .I(N__18614));
    LocalMux I__3844 (
            .O(N__18617),
            .I(N__18611));
    Odrv4 I__3843 (
            .O(N__18614),
            .I(\Lab_UT.dictrl.N_39 ));
    Odrv12 I__3842 (
            .O(N__18611),
            .I(\Lab_UT.dictrl.N_39 ));
    CascadeMux I__3841 (
            .O(N__18606),
            .I(N__18599));
    CascadeMux I__3840 (
            .O(N__18605),
            .I(N__18596));
    CascadeMux I__3839 (
            .O(N__18604),
            .I(N__18591));
    CascadeMux I__3838 (
            .O(N__18603),
            .I(N__18588));
    InMux I__3837 (
            .O(N__18602),
            .I(N__18580));
    InMux I__3836 (
            .O(N__18599),
            .I(N__18580));
    InMux I__3835 (
            .O(N__18596),
            .I(N__18577));
    InMux I__3834 (
            .O(N__18595),
            .I(N__18574));
    InMux I__3833 (
            .O(N__18594),
            .I(N__18571));
    InMux I__3832 (
            .O(N__18591),
            .I(N__18566));
    InMux I__3831 (
            .O(N__18588),
            .I(N__18563));
    InMux I__3830 (
            .O(N__18587),
            .I(N__18560));
    InMux I__3829 (
            .O(N__18586),
            .I(N__18556));
    CascadeMux I__3828 (
            .O(N__18585),
            .I(N__18553));
    LocalMux I__3827 (
            .O(N__18580),
            .I(N__18548));
    LocalMux I__3826 (
            .O(N__18577),
            .I(N__18548));
    LocalMux I__3825 (
            .O(N__18574),
            .I(N__18545));
    LocalMux I__3824 (
            .O(N__18571),
            .I(N__18542));
    InMux I__3823 (
            .O(N__18570),
            .I(N__18537));
    InMux I__3822 (
            .O(N__18569),
            .I(N__18537));
    LocalMux I__3821 (
            .O(N__18566),
            .I(N__18532));
    LocalMux I__3820 (
            .O(N__18563),
            .I(N__18532));
    LocalMux I__3819 (
            .O(N__18560),
            .I(N__18529));
    InMux I__3818 (
            .O(N__18559),
            .I(N__18526));
    LocalMux I__3817 (
            .O(N__18556),
            .I(N__18523));
    InMux I__3816 (
            .O(N__18553),
            .I(N__18520));
    Span4Mux_v I__3815 (
            .O(N__18548),
            .I(N__18517));
    Span4Mux_v I__3814 (
            .O(N__18545),
            .I(N__18512));
    Span4Mux_v I__3813 (
            .O(N__18542),
            .I(N__18512));
    LocalMux I__3812 (
            .O(N__18537),
            .I(N__18509));
    Span4Mux_s3_v I__3811 (
            .O(N__18532),
            .I(N__18506));
    Span4Mux_h I__3810 (
            .O(N__18529),
            .I(N__18503));
    LocalMux I__3809 (
            .O(N__18526),
            .I(N__18496));
    Span4Mux_v I__3808 (
            .O(N__18523),
            .I(N__18496));
    LocalMux I__3807 (
            .O(N__18520),
            .I(N__18496));
    Span4Mux_v I__3806 (
            .O(N__18517),
            .I(N__18491));
    Span4Mux_v I__3805 (
            .O(N__18512),
            .I(N__18491));
    Span4Mux_v I__3804 (
            .O(N__18509),
            .I(N__18488));
    Span4Mux_v I__3803 (
            .O(N__18506),
            .I(N__18485));
    Span4Mux_v I__3802 (
            .O(N__18503),
            .I(N__18480));
    Span4Mux_h I__3801 (
            .O(N__18496),
            .I(N__18480));
    Odrv4 I__3800 (
            .O(N__18491),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__3799 (
            .O(N__18488),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__3798 (
            .O(N__18485),
            .I(bu_rx_data_6_rep1));
    Odrv4 I__3797 (
            .O(N__18480),
            .I(bu_rx_data_6_rep1));
    InMux I__3796 (
            .O(N__18471),
            .I(N__18468));
    LocalMux I__3795 (
            .O(N__18468),
            .I(N__18465));
    Span4Mux_h I__3794 (
            .O(N__18465),
            .I(N__18462));
    Odrv4 I__3793 (
            .O(N__18462),
            .I(\Lab_UT.dictrl.m53_d_1_0 ));
    CascadeMux I__3792 (
            .O(N__18459),
            .I(\Lab_UT.dictrl.N_97_mux_2_cascade_ ));
    InMux I__3791 (
            .O(N__18456),
            .I(N__18453));
    LocalMux I__3790 (
            .O(N__18453),
            .I(N__18450));
    Span4Mux_v I__3789 (
            .O(N__18450),
            .I(N__18447));
    Odrv4 I__3788 (
            .O(N__18447),
            .I(\Lab_UT.dictrl.g2_1 ));
    InMux I__3787 (
            .O(N__18444),
            .I(N__18441));
    LocalMux I__3786 (
            .O(N__18441),
            .I(N__18438));
    Odrv4 I__3785 (
            .O(N__18438),
            .I(\Lab_UT.dictrl.N_1462_0 ));
    CascadeMux I__3784 (
            .O(N__18435),
            .I(\Lab_UT.dictrl.N_1102_0_cascade_ ));
    CascadeMux I__3783 (
            .O(N__18432),
            .I(N__18428));
    InMux I__3782 (
            .O(N__18431),
            .I(N__18425));
    InMux I__3781 (
            .O(N__18428),
            .I(N__18422));
    LocalMux I__3780 (
            .O(N__18425),
            .I(\Lab_UT.dictrl.N_97_mux_7 ));
    LocalMux I__3779 (
            .O(N__18422),
            .I(\Lab_UT.dictrl.N_97_mux_7 ));
    CascadeMux I__3778 (
            .O(N__18417),
            .I(\Lab_UT.dictrl.N_1106_1_cascade_ ));
    CascadeMux I__3777 (
            .O(N__18414),
            .I(\Lab_UT.didp.countrce4.q_5_0_cascade_ ));
    InMux I__3776 (
            .O(N__18411),
            .I(N__18408));
    LocalMux I__3775 (
            .O(N__18408),
            .I(N__18403));
    InMux I__3774 (
            .O(N__18407),
            .I(N__18400));
    CascadeMux I__3773 (
            .O(N__18406),
            .I(N__18396));
    Span4Mux_h I__3772 (
            .O(N__18403),
            .I(N__18392));
    LocalMux I__3771 (
            .O(N__18400),
            .I(N__18389));
    InMux I__3770 (
            .O(N__18399),
            .I(N__18382));
    InMux I__3769 (
            .O(N__18396),
            .I(N__18382));
    InMux I__3768 (
            .O(N__18395),
            .I(N__18382));
    Odrv4 I__3767 (
            .O(N__18392),
            .I(\Lab_UT.LdMtens ));
    Odrv4 I__3766 (
            .O(N__18389),
            .I(\Lab_UT.LdMtens ));
    LocalMux I__3765 (
            .O(N__18382),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__3764 (
            .O(N__18375),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__3763 (
            .O(N__18372),
            .I(N__18368));
    InMux I__3762 (
            .O(N__18371),
            .I(N__18365));
    LocalMux I__3761 (
            .O(N__18368),
            .I(N__18360));
    LocalMux I__3760 (
            .O(N__18365),
            .I(N__18360));
    Span4Mux_h I__3759 (
            .O(N__18360),
            .I(N__18356));
    InMux I__3758 (
            .O(N__18359),
            .I(N__18353));
    Odrv4 I__3757 (
            .O(N__18356),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    LocalMux I__3756 (
            .O(N__18353),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    CascadeMux I__3755 (
            .O(N__18348),
            .I(N__18342));
    InMux I__3754 (
            .O(N__18347),
            .I(N__18328));
    InMux I__3753 (
            .O(N__18346),
            .I(N__18328));
    InMux I__3752 (
            .O(N__18345),
            .I(N__18328));
    InMux I__3751 (
            .O(N__18342),
            .I(N__18328));
    InMux I__3750 (
            .O(N__18341),
            .I(N__18325));
    InMux I__3749 (
            .O(N__18340),
            .I(N__18316));
    InMux I__3748 (
            .O(N__18339),
            .I(N__18316));
    InMux I__3747 (
            .O(N__18338),
            .I(N__18313));
    InMux I__3746 (
            .O(N__18337),
            .I(N__18310));
    LocalMux I__3745 (
            .O(N__18328),
            .I(N__18307));
    LocalMux I__3744 (
            .O(N__18325),
            .I(N__18304));
    InMux I__3743 (
            .O(N__18324),
            .I(N__18297));
    InMux I__3742 (
            .O(N__18323),
            .I(N__18297));
    InMux I__3741 (
            .O(N__18322),
            .I(N__18297));
    InMux I__3740 (
            .O(N__18321),
            .I(N__18294));
    LocalMux I__3739 (
            .O(N__18316),
            .I(N__18291));
    LocalMux I__3738 (
            .O(N__18313),
            .I(N__18288));
    LocalMux I__3737 (
            .O(N__18310),
            .I(N__18284));
    Span4Mux_v I__3736 (
            .O(N__18307),
            .I(N__18275));
    Span4Mux_s3_v I__3735 (
            .O(N__18304),
            .I(N__18275));
    LocalMux I__3734 (
            .O(N__18297),
            .I(N__18275));
    LocalMux I__3733 (
            .O(N__18294),
            .I(N__18275));
    Span4Mux_s3_h I__3732 (
            .O(N__18291),
            .I(N__18272));
    Span4Mux_v I__3731 (
            .O(N__18288),
            .I(N__18268));
    InMux I__3730 (
            .O(N__18287),
            .I(N__18265));
    Span4Mux_h I__3729 (
            .O(N__18284),
            .I(N__18260));
    Span4Mux_h I__3728 (
            .O(N__18275),
            .I(N__18260));
    Span4Mux_h I__3727 (
            .O(N__18272),
            .I(N__18257));
    InMux I__3726 (
            .O(N__18271),
            .I(N__18254));
    Odrv4 I__3725 (
            .O(N__18268),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    LocalMux I__3724 (
            .O(N__18265),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv4 I__3723 (
            .O(N__18260),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv4 I__3722 (
            .O(N__18257),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    LocalMux I__3721 (
            .O(N__18254),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    InMux I__3720 (
            .O(N__18243),
            .I(N__18240));
    LocalMux I__3719 (
            .O(N__18240),
            .I(N__18237));
    Odrv4 I__3718 (
            .O(N__18237),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0 ));
    InMux I__3717 (
            .O(N__18234),
            .I(N__18229));
    InMux I__3716 (
            .O(N__18233),
            .I(N__18226));
    InMux I__3715 (
            .O(N__18232),
            .I(N__18221));
    LocalMux I__3714 (
            .O(N__18229),
            .I(N__18218));
    LocalMux I__3713 (
            .O(N__18226),
            .I(N__18214));
    InMux I__3712 (
            .O(N__18225),
            .I(N__18211));
    CascadeMux I__3711 (
            .O(N__18224),
            .I(N__18208));
    LocalMux I__3710 (
            .O(N__18221),
            .I(N__18203));
    Span4Mux_v I__3709 (
            .O(N__18218),
            .I(N__18203));
    CascadeMux I__3708 (
            .O(N__18217),
            .I(N__18200));
    Span4Mux_v I__3707 (
            .O(N__18214),
            .I(N__18194));
    LocalMux I__3706 (
            .O(N__18211),
            .I(N__18194));
    InMux I__3705 (
            .O(N__18208),
            .I(N__18191));
    Span4Mux_h I__3704 (
            .O(N__18203),
            .I(N__18188));
    InMux I__3703 (
            .O(N__18200),
            .I(N__18185));
    InMux I__3702 (
            .O(N__18199),
            .I(N__18182));
    Odrv4 I__3701 (
            .O(N__18194),
            .I(\Lab_UT.state_i_4_0 ));
    LocalMux I__3700 (
            .O(N__18191),
            .I(\Lab_UT.state_i_4_0 ));
    Odrv4 I__3699 (
            .O(N__18188),
            .I(\Lab_UT.state_i_4_0 ));
    LocalMux I__3698 (
            .O(N__18185),
            .I(\Lab_UT.state_i_4_0 ));
    LocalMux I__3697 (
            .O(N__18182),
            .I(\Lab_UT.state_i_4_0 ));
    InMux I__3696 (
            .O(N__18171),
            .I(N__18167));
    InMux I__3695 (
            .O(N__18170),
            .I(N__18164));
    LocalMux I__3694 (
            .O(N__18167),
            .I(\Lab_UT.dicRun_2 ));
    LocalMux I__3693 (
            .O(N__18164),
            .I(\Lab_UT.dicRun_2 ));
    InMux I__3692 (
            .O(N__18159),
            .I(N__18145));
    InMux I__3691 (
            .O(N__18158),
            .I(N__18145));
    CascadeMux I__3690 (
            .O(N__18157),
            .I(N__18142));
    InMux I__3689 (
            .O(N__18156),
            .I(N__18138));
    InMux I__3688 (
            .O(N__18155),
            .I(N__18130));
    InMux I__3687 (
            .O(N__18154),
            .I(N__18130));
    InMux I__3686 (
            .O(N__18153),
            .I(N__18130));
    CascadeMux I__3685 (
            .O(N__18152),
            .I(N__18126));
    InMux I__3684 (
            .O(N__18151),
            .I(N__18123));
    InMux I__3683 (
            .O(N__18150),
            .I(N__18120));
    LocalMux I__3682 (
            .O(N__18145),
            .I(N__18117));
    InMux I__3681 (
            .O(N__18142),
            .I(N__18114));
    CascadeMux I__3680 (
            .O(N__18141),
            .I(N__18111));
    LocalMux I__3679 (
            .O(N__18138),
            .I(N__18108));
    InMux I__3678 (
            .O(N__18137),
            .I(N__18105));
    LocalMux I__3677 (
            .O(N__18130),
            .I(N__18102));
    InMux I__3676 (
            .O(N__18129),
            .I(N__18099));
    InMux I__3675 (
            .O(N__18126),
            .I(N__18096));
    LocalMux I__3674 (
            .O(N__18123),
            .I(N__18087));
    LocalMux I__3673 (
            .O(N__18120),
            .I(N__18087));
    Span4Mux_h I__3672 (
            .O(N__18117),
            .I(N__18087));
    LocalMux I__3671 (
            .O(N__18114),
            .I(N__18087));
    InMux I__3670 (
            .O(N__18111),
            .I(N__18084));
    Span4Mux_v I__3669 (
            .O(N__18108),
            .I(N__18079));
    LocalMux I__3668 (
            .O(N__18105),
            .I(N__18079));
    Span4Mux_h I__3667 (
            .O(N__18102),
            .I(N__18076));
    LocalMux I__3666 (
            .O(N__18099),
            .I(N__18071));
    LocalMux I__3665 (
            .O(N__18096),
            .I(N__18071));
    Span4Mux_v I__3664 (
            .O(N__18087),
            .I(N__18066));
    LocalMux I__3663 (
            .O(N__18084),
            .I(N__18066));
    Span4Mux_h I__3662 (
            .O(N__18079),
            .I(N__18063));
    Span4Mux_h I__3661 (
            .O(N__18076),
            .I(N__18060));
    Span4Mux_v I__3660 (
            .O(N__18071),
            .I(N__18055));
    Span4Mux_h I__3659 (
            .O(N__18066),
            .I(N__18055));
    Odrv4 I__3658 (
            .O(N__18063),
            .I(bu_rx_data_7));
    Odrv4 I__3657 (
            .O(N__18060),
            .I(bu_rx_data_7));
    Odrv4 I__3656 (
            .O(N__18055),
            .I(bu_rx_data_7));
    InMux I__3655 (
            .O(N__18048),
            .I(N__18045));
    LocalMux I__3654 (
            .O(N__18045),
            .I(N__18042));
    Odrv4 I__3653 (
            .O(N__18042),
            .I(\Lab_UT.didp.countrce1.q_5_1 ));
    InMux I__3652 (
            .O(N__18039),
            .I(N__18036));
    LocalMux I__3651 (
            .O(N__18036),
            .I(N__18033));
    Span4Mux_h I__3650 (
            .O(N__18033),
            .I(N__18029));
    InMux I__3649 (
            .O(N__18032),
            .I(N__18026));
    Odrv4 I__3648 (
            .O(N__18029),
            .I(\Lab_UT.LdASones ));
    LocalMux I__3647 (
            .O(N__18026),
            .I(\Lab_UT.LdASones ));
    CEMux I__3646 (
            .O(N__18021),
            .I(N__18018));
    LocalMux I__3645 (
            .O(N__18018),
            .I(N__18015));
    Span4Mux_h I__3644 (
            .O(N__18015),
            .I(N__18011));
    CEMux I__3643 (
            .O(N__18014),
            .I(N__18008));
    Odrv4 I__3642 (
            .O(N__18011),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    LocalMux I__3641 (
            .O(N__18008),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    InMux I__3640 (
            .O(N__18003),
            .I(N__18000));
    LocalMux I__3639 (
            .O(N__18000),
            .I(N__17995));
    InMux I__3638 (
            .O(N__17999),
            .I(N__17992));
    InMux I__3637 (
            .O(N__17998),
            .I(N__17989));
    Odrv4 I__3636 (
            .O(N__17995),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__3635 (
            .O(N__17992),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__3634 (
            .O(N__17989),
            .I(\Lab_UT.di_ASones_0 ));
    CascadeMux I__3633 (
            .O(N__17982),
            .I(N__17979));
    InMux I__3632 (
            .O(N__17979),
            .I(N__17976));
    LocalMux I__3631 (
            .O(N__17976),
            .I(N__17973));
    Odrv12 I__3630 (
            .O(N__17973),
            .I(\Lab_UT.dispString.N_180 ));
    InMux I__3629 (
            .O(N__17970),
            .I(N__17967));
    LocalMux I__3628 (
            .O(N__17967),
            .I(\Lab_UT.dispString.m49Z0Z_7 ));
    InMux I__3627 (
            .O(N__17964),
            .I(N__17961));
    LocalMux I__3626 (
            .O(N__17961),
            .I(\Lab_UT.dispString.m49Z0Z_11 ));
    CascadeMux I__3625 (
            .O(N__17958),
            .I(\Lab_UT.didp.countrce1.q_5_0_cascade_ ));
    CascadeMux I__3624 (
            .O(N__17955),
            .I(N__17950));
    CascadeMux I__3623 (
            .O(N__17954),
            .I(N__17947));
    InMux I__3622 (
            .O(N__17953),
            .I(N__17940));
    InMux I__3621 (
            .O(N__17950),
            .I(N__17940));
    InMux I__3620 (
            .O(N__17947),
            .I(N__17940));
    LocalMux I__3619 (
            .O(N__17940),
            .I(N__17932));
    InMux I__3618 (
            .O(N__17939),
            .I(N__17929));
    InMux I__3617 (
            .O(N__17938),
            .I(N__17920));
    InMux I__3616 (
            .O(N__17937),
            .I(N__17920));
    InMux I__3615 (
            .O(N__17936),
            .I(N__17920));
    InMux I__3614 (
            .O(N__17935),
            .I(N__17920));
    Odrv4 I__3613 (
            .O(N__17932),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3612 (
            .O(N__17929),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3611 (
            .O(N__17920),
            .I(\Lab_UT.di_Sones_0 ));
    CascadeMux I__3610 (
            .O(N__17913),
            .I(\Lab_UT.LdMtens_cascade_ ));
    CascadeMux I__3609 (
            .O(N__17910),
            .I(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ));
    CascadeMux I__3608 (
            .O(N__17907),
            .I(\Lab_UT.didp.countrce1.q_5_2_cascade_ ));
    InMux I__3607 (
            .O(N__17904),
            .I(N__17896));
    InMux I__3606 (
            .O(N__17903),
            .I(N__17889));
    InMux I__3605 (
            .O(N__17902),
            .I(N__17889));
    InMux I__3604 (
            .O(N__17901),
            .I(N__17889));
    InMux I__3603 (
            .O(N__17900),
            .I(N__17886));
    InMux I__3602 (
            .O(N__17899),
            .I(N__17883));
    LocalMux I__3601 (
            .O(N__17896),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3600 (
            .O(N__17889),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3599 (
            .O(N__17886),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3598 (
            .O(N__17883),
            .I(\Lab_UT.di_Sones_2 ));
    InMux I__3597 (
            .O(N__17874),
            .I(N__17871));
    LocalMux I__3596 (
            .O(N__17871),
            .I(\Lab_UT.dispString.m49Z0Z_12 ));
    CascadeMux I__3595 (
            .O(N__17868),
            .I(\Lab_UT.dispString.m49Z0Z_4_cascade_ ));
    InMux I__3594 (
            .O(N__17865),
            .I(N__17861));
    InMux I__3593 (
            .O(N__17864),
            .I(N__17858));
    LocalMux I__3592 (
            .O(N__17861),
            .I(N__17853));
    LocalMux I__3591 (
            .O(N__17858),
            .I(N__17853));
    Odrv12 I__3590 (
            .O(N__17853),
            .I(\Lab_UT.dispString.N_128_mux ));
    InMux I__3589 (
            .O(N__17850),
            .I(N__17847));
    LocalMux I__3588 (
            .O(N__17847),
            .I(N__17842));
    InMux I__3587 (
            .O(N__17846),
            .I(N__17837));
    InMux I__3586 (
            .O(N__17845),
            .I(N__17837));
    Odrv4 I__3585 (
            .O(N__17842),
            .I(\Lab_UT.di_AStens_2 ));
    LocalMux I__3584 (
            .O(N__17837),
            .I(\Lab_UT.di_AStens_2 ));
    InMux I__3583 (
            .O(N__17832),
            .I(N__17829));
    LocalMux I__3582 (
            .O(N__17829),
            .I(N__17825));
    InMux I__3581 (
            .O(N__17828),
            .I(N__17822));
    Span4Mux_v I__3580 (
            .O(N__17825),
            .I(N__17818));
    LocalMux I__3579 (
            .O(N__17822),
            .I(N__17815));
    InMux I__3578 (
            .O(N__17821),
            .I(N__17812));
    Odrv4 I__3577 (
            .O(N__17818),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__3576 (
            .O(N__17815),
            .I(\Lab_UT.di_ASones_2 ));
    LocalMux I__3575 (
            .O(N__17812),
            .I(\Lab_UT.di_ASones_2 ));
    InMux I__3574 (
            .O(N__17805),
            .I(N__17802));
    LocalMux I__3573 (
            .O(N__17802),
            .I(N__17794));
    InMux I__3572 (
            .O(N__17801),
            .I(N__17791));
    InMux I__3571 (
            .O(N__17800),
            .I(N__17782));
    InMux I__3570 (
            .O(N__17799),
            .I(N__17782));
    InMux I__3569 (
            .O(N__17798),
            .I(N__17782));
    InMux I__3568 (
            .O(N__17797),
            .I(N__17782));
    Span4Mux_h I__3567 (
            .O(N__17794),
            .I(N__17777));
    LocalMux I__3566 (
            .O(N__17791),
            .I(N__17777));
    LocalMux I__3565 (
            .O(N__17782),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3564 (
            .O(N__17777),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    CascadeMux I__3563 (
            .O(N__17772),
            .I(N__17769));
    InMux I__3562 (
            .O(N__17769),
            .I(N__17766));
    LocalMux I__3561 (
            .O(N__17766),
            .I(N__17763));
    Odrv4 I__3560 (
            .O(N__17763),
            .I(\uu2.N_15 ));
    InMux I__3559 (
            .O(N__17760),
            .I(N__17757));
    LocalMux I__3558 (
            .O(N__17757),
            .I(\uu2.N_17 ));
    CascadeMux I__3557 (
            .O(N__17754),
            .I(\uu2.bitmap_pmux_25_i_m2_ns_1_cascade_ ));
    CascadeMux I__3556 (
            .O(N__17751),
            .I(N__17748));
    InMux I__3555 (
            .O(N__17748),
            .I(N__17745));
    LocalMux I__3554 (
            .O(N__17745),
            .I(N__17742));
    Odrv4 I__3553 (
            .O(N__17742),
            .I(\uu2.N_49 ));
    InMux I__3552 (
            .O(N__17739),
            .I(N__17736));
    LocalMux I__3551 (
            .O(N__17736),
            .I(\uu2.bitmapZ0Z_221 ));
    InMux I__3550 (
            .O(N__17733),
            .I(N__17730));
    LocalMux I__3549 (
            .O(N__17730),
            .I(\uu2.bitmapZ0Z_93 ));
    InMux I__3548 (
            .O(N__17727),
            .I(N__17724));
    LocalMux I__3547 (
            .O(N__17724),
            .I(\uu2.N_13 ));
    CascadeMux I__3546 (
            .O(N__17721),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    CascadeMux I__3545 (
            .O(N__17718),
            .I(\Lab_UT.didp.countrce1.q_5_3_cascade_ ));
    CascadeMux I__3544 (
            .O(N__17715),
            .I(N__17708));
    InMux I__3543 (
            .O(N__17714),
            .I(N__17705));
    InMux I__3542 (
            .O(N__17713),
            .I(N__17700));
    InMux I__3541 (
            .O(N__17712),
            .I(N__17700));
    InMux I__3540 (
            .O(N__17711),
            .I(N__17695));
    InMux I__3539 (
            .O(N__17708),
            .I(N__17695));
    LocalMux I__3538 (
            .O(N__17705),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3537 (
            .O(N__17700),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3536 (
            .O(N__17695),
            .I(\Lab_UT.di_Sones_3 ));
    InMux I__3535 (
            .O(N__17688),
            .I(N__17682));
    InMux I__3534 (
            .O(N__17687),
            .I(N__17682));
    LocalMux I__3533 (
            .O(N__17682),
            .I(\uu2.w_addr_displaying_0_rep1_RNIDASJZ0 ));
    CascadeMux I__3532 (
            .O(N__17679),
            .I(N__17676));
    InMux I__3531 (
            .O(N__17676),
            .I(N__17673));
    LocalMux I__3530 (
            .O(N__17673),
            .I(\uu2.w_addr_displaying_RNIR2PLZ0Z_8 ));
    InMux I__3529 (
            .O(N__17670),
            .I(N__17667));
    LocalMux I__3528 (
            .O(N__17667),
            .I(\uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1 ));
    InMux I__3527 (
            .O(N__17664),
            .I(N__17661));
    LocalMux I__3526 (
            .O(N__17661),
            .I(N__17658));
    Odrv4 I__3525 (
            .O(N__17658),
            .I(\uu2.bitmap_pmux_29_0 ));
    InMux I__3524 (
            .O(N__17655),
            .I(N__17650));
    InMux I__3523 (
            .O(N__17654),
            .I(N__17647));
    InMux I__3522 (
            .O(N__17653),
            .I(N__17644));
    LocalMux I__3521 (
            .O(N__17650),
            .I(\uu2.N_24_0 ));
    LocalMux I__3520 (
            .O(N__17647),
            .I(\uu2.N_24_0 ));
    LocalMux I__3519 (
            .O(N__17644),
            .I(\uu2.N_24_0 ));
    InMux I__3518 (
            .O(N__17637),
            .I(N__17634));
    LocalMux I__3517 (
            .O(N__17634),
            .I(\uu2.w_addr_displaying_RNIU1AF7Z0Z_0 ));
    InMux I__3516 (
            .O(N__17631),
            .I(N__17625));
    InMux I__3515 (
            .O(N__17630),
            .I(N__17625));
    LocalMux I__3514 (
            .O(N__17625),
            .I(N__17622));
    Span4Mux_h I__3513 (
            .O(N__17622),
            .I(N__17619));
    Span4Mux_v I__3512 (
            .O(N__17619),
            .I(N__17616));
    Odrv4 I__3511 (
            .O(N__17616),
            .I(\Lab_UT.dictrl.m12Z0Z_2 ));
    InMux I__3510 (
            .O(N__17613),
            .I(N__17610));
    LocalMux I__3509 (
            .O(N__17610),
            .I(\uu2.bitmapZ0Z_215 ));
    CascadeMux I__3508 (
            .O(N__17607),
            .I(\uu2.N_198_cascade_ ));
    InMux I__3507 (
            .O(N__17604),
            .I(N__17601));
    LocalMux I__3506 (
            .O(N__17601),
            .I(N__17598));
    Odrv4 I__3505 (
            .O(N__17598),
            .I(\uu2.N_199 ));
    CascadeMux I__3504 (
            .O(N__17595),
            .I(\uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_ ));
    InMux I__3503 (
            .O(N__17592),
            .I(N__17589));
    LocalMux I__3502 (
            .O(N__17589),
            .I(\uu2.N_196 ));
    InMux I__3501 (
            .O(N__17586),
            .I(N__17583));
    LocalMux I__3500 (
            .O(N__17583),
            .I(\uu2.bitmap_pmux_27_i_m2_ns_1 ));
    InMux I__3499 (
            .O(N__17580),
            .I(N__17577));
    LocalMux I__3498 (
            .O(N__17577),
            .I(N__17574));
    Span4Mux_s3_v I__3497 (
            .O(N__17574),
            .I(N__17571));
    Odrv4 I__3496 (
            .O(N__17571),
            .I(\Lab_UT.dictrl.m53_d_1_1 ));
    CascadeMux I__3495 (
            .O(N__17568),
            .I(\Lab_UT.dictrl.N_97_mux_3_cascade_ ));
    InMux I__3494 (
            .O(N__17565),
            .I(N__17562));
    LocalMux I__3493 (
            .O(N__17562),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    CascadeMux I__3492 (
            .O(N__17559),
            .I(N__17552));
    InMux I__3491 (
            .O(N__17558),
            .I(N__17548));
    InMux I__3490 (
            .O(N__17557),
            .I(N__17545));
    InMux I__3489 (
            .O(N__17556),
            .I(N__17540));
    InMux I__3488 (
            .O(N__17555),
            .I(N__17540));
    InMux I__3487 (
            .O(N__17552),
            .I(N__17535));
    InMux I__3486 (
            .O(N__17551),
            .I(N__17535));
    LocalMux I__3485 (
            .O(N__17548),
            .I(N__17532));
    LocalMux I__3484 (
            .O(N__17545),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__3483 (
            .O(N__17540),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__3482 (
            .O(N__17535),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv12 I__3481 (
            .O(N__17532),
            .I(\uu2.w_addr_userZ0Z_1 ));
    InMux I__3480 (
            .O(N__17523),
            .I(N__17519));
    CascadeMux I__3479 (
            .O(N__17522),
            .I(N__17515));
    LocalMux I__3478 (
            .O(N__17519),
            .I(N__17510));
    InMux I__3477 (
            .O(N__17518),
            .I(N__17507));
    InMux I__3476 (
            .O(N__17515),
            .I(N__17502));
    InMux I__3475 (
            .O(N__17514),
            .I(N__17502));
    InMux I__3474 (
            .O(N__17513),
            .I(N__17499));
    Span4Mux_s0_v I__3473 (
            .O(N__17510),
            .I(N__17496));
    LocalMux I__3472 (
            .O(N__17507),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__3471 (
            .O(N__17502),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__3470 (
            .O(N__17499),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__3469 (
            .O(N__17496),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__3468 (
            .O(N__17487),
            .I(\uu2.un3_w_addr_user_4_cascade_ ));
    InMux I__3467 (
            .O(N__17484),
            .I(N__17481));
    LocalMux I__3466 (
            .O(N__17481),
            .I(N__17478));
    Span4Mux_s1_v I__3465 (
            .O(N__17478),
            .I(N__17475));
    Odrv4 I__3464 (
            .O(N__17475),
            .I(\uu2.un3_w_addr_user_5 ));
    CascadeMux I__3463 (
            .O(N__17472),
            .I(N__17469));
    InMux I__3462 (
            .O(N__17469),
            .I(N__17465));
    InMux I__3461 (
            .O(N__17468),
            .I(N__17462));
    LocalMux I__3460 (
            .O(N__17465),
            .I(N__17457));
    LocalMux I__3459 (
            .O(N__17462),
            .I(N__17457));
    IoSpan4Mux I__3458 (
            .O(N__17457),
            .I(N__17454));
    Span4Mux_s0_v I__3457 (
            .O(N__17454),
            .I(N__17451));
    Odrv4 I__3456 (
            .O(N__17451),
            .I(\uu2.un3_w_addr_user ));
    CEMux I__3455 (
            .O(N__17448),
            .I(N__17445));
    LocalMux I__3454 (
            .O(N__17445),
            .I(N__17442));
    Span4Mux_s0_v I__3453 (
            .O(N__17442),
            .I(N__17439));
    Span4Mux_h I__3452 (
            .O(N__17439),
            .I(N__17436));
    Odrv4 I__3451 (
            .O(N__17436),
            .I(\uu2.un21_w_addr_displaying_0_0 ));
    InMux I__3450 (
            .O(N__17433),
            .I(N__17430));
    LocalMux I__3449 (
            .O(N__17430),
            .I(N__17427));
    Span4Mux_s1_v I__3448 (
            .O(N__17427),
            .I(N__17424));
    Odrv4 I__3447 (
            .O(N__17424),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    CascadeMux I__3446 (
            .O(N__17421),
            .I(N__17416));
    CascadeMux I__3445 (
            .O(N__17420),
            .I(N__17410));
    InMux I__3444 (
            .O(N__17419),
            .I(N__17402));
    InMux I__3443 (
            .O(N__17416),
            .I(N__17402));
    InMux I__3442 (
            .O(N__17415),
            .I(N__17402));
    InMux I__3441 (
            .O(N__17414),
            .I(N__17393));
    InMux I__3440 (
            .O(N__17413),
            .I(N__17393));
    InMux I__3439 (
            .O(N__17410),
            .I(N__17393));
    InMux I__3438 (
            .O(N__17409),
            .I(N__17393));
    LocalMux I__3437 (
            .O(N__17402),
            .I(N__17390));
    LocalMux I__3436 (
            .O(N__17393),
            .I(\uu2.w_addr_displayingZ1Z_4 ));
    Odrv4 I__3435 (
            .O(N__17390),
            .I(\uu2.w_addr_displayingZ1Z_4 ));
    CascadeMux I__3434 (
            .O(N__17385),
            .I(\uu2.bitmap_pmux_sn_N_33_cascade_ ));
    CascadeMux I__3433 (
            .O(N__17382),
            .I(N__17378));
    CascadeMux I__3432 (
            .O(N__17381),
            .I(N__17371));
    InMux I__3431 (
            .O(N__17378),
            .I(N__17368));
    CascadeMux I__3430 (
            .O(N__17377),
            .I(N__17363));
    CascadeMux I__3429 (
            .O(N__17376),
            .I(N__17360));
    InMux I__3428 (
            .O(N__17375),
            .I(N__17353));
    InMux I__3427 (
            .O(N__17374),
            .I(N__17353));
    InMux I__3426 (
            .O(N__17371),
            .I(N__17353));
    LocalMux I__3425 (
            .O(N__17368),
            .I(N__17350));
    InMux I__3424 (
            .O(N__17367),
            .I(N__17345));
    InMux I__3423 (
            .O(N__17366),
            .I(N__17345));
    InMux I__3422 (
            .O(N__17363),
            .I(N__17342));
    InMux I__3421 (
            .O(N__17360),
            .I(N__17339));
    LocalMux I__3420 (
            .O(N__17353),
            .I(N__17334));
    Span4Mux_s1_v I__3419 (
            .O(N__17350),
            .I(N__17334));
    LocalMux I__3418 (
            .O(N__17345),
            .I(N__17331));
    LocalMux I__3417 (
            .O(N__17342),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__3416 (
            .O(N__17339),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__3415 (
            .O(N__17334),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__3414 (
            .O(N__17331),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__3413 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__3412 (
            .O(N__17319),
            .I(N__17316));
    Span4Mux_s1_v I__3411 (
            .O(N__17316),
            .I(N__17313));
    Odrv4 I__3410 (
            .O(N__17313),
            .I(\uu2.bitmap_pmux_sn_m15_0_1 ));
    InMux I__3409 (
            .O(N__17310),
            .I(N__17307));
    LocalMux I__3408 (
            .O(N__17307),
            .I(\Lab_UT.dictrl.g1_1 ));
    InMux I__3407 (
            .O(N__17304),
            .I(N__17301));
    LocalMux I__3406 (
            .O(N__17301),
            .I(N__17298));
    Odrv4 I__3405 (
            .O(N__17298),
            .I(\Lab_UT.dictrl.N_5 ));
    CascadeMux I__3404 (
            .O(N__17295),
            .I(\Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_ ));
    InMux I__3403 (
            .O(N__17292),
            .I(N__17289));
    LocalMux I__3402 (
            .O(N__17289),
            .I(N__17286));
    Odrv4 I__3401 (
            .O(N__17286),
            .I(\Lab_UT.dictrl.N_9 ));
    InMux I__3400 (
            .O(N__17283),
            .I(N__17280));
    LocalMux I__3399 (
            .O(N__17280),
            .I(\Lab_UT.dictrl.g2_1_3 ));
    CascadeMux I__3398 (
            .O(N__17277),
            .I(\Lab_UT.dictrl.N_1462_3_cascade_ ));
    InMux I__3397 (
            .O(N__17274),
            .I(N__17271));
    LocalMux I__3396 (
            .O(N__17271),
            .I(\Lab_UT.dictrl.N_1102_3 ));
    InMux I__3395 (
            .O(N__17268),
            .I(N__17265));
    LocalMux I__3394 (
            .O(N__17265),
            .I(\Lab_UT.dictrl.N_1460_3 ));
    InMux I__3393 (
            .O(N__17262),
            .I(N__17259));
    LocalMux I__3392 (
            .O(N__17259),
            .I(N__17256));
    Odrv12 I__3391 (
            .O(N__17256),
            .I(\Lab_UT.dictrl.N_6 ));
    CascadeMux I__3390 (
            .O(N__17253),
            .I(\Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_ ));
    InMux I__3389 (
            .O(N__17250),
            .I(N__17247));
    LocalMux I__3388 (
            .O(N__17247),
            .I(\Lab_UT.dictrl.g0_i_m2_i_1 ));
    InMux I__3387 (
            .O(N__17244),
            .I(N__17241));
    LocalMux I__3386 (
            .O(N__17241),
            .I(\Lab_UT.dictrl.N_97_mux_1 ));
    InMux I__3385 (
            .O(N__17238),
            .I(N__17235));
    LocalMux I__3384 (
            .O(N__17235),
            .I(N__17232));
    Odrv12 I__3383 (
            .O(N__17232),
            .I(\Lab_UT.dictrl.g0_i_a5_0_2 ));
    CascadeMux I__3382 (
            .O(N__17229),
            .I(N__17226));
    InMux I__3381 (
            .O(N__17226),
            .I(N__17223));
    LocalMux I__3380 (
            .O(N__17223),
            .I(N__17220));
    Odrv12 I__3379 (
            .O(N__17220),
            .I(\Lab_UT.dictrl.g2_2 ));
    CascadeMux I__3378 (
            .O(N__17217),
            .I(\Lab_UT.dictrl.g2_3_cascade_ ));
    InMux I__3377 (
            .O(N__17214),
            .I(N__17211));
    LocalMux I__3376 (
            .O(N__17211),
            .I(N__17208));
    Odrv12 I__3375 (
            .O(N__17208),
            .I(\Lab_UT.dictrl.next_state_3_1 ));
    InMux I__3374 (
            .O(N__17205),
            .I(N__17202));
    LocalMux I__3373 (
            .O(N__17202),
            .I(N__17199));
    Span4Mux_h I__3372 (
            .O(N__17199),
            .I(N__17196));
    Odrv4 I__3371 (
            .O(N__17196),
            .I(\Lab_UT.dictrl.g0_12_a6_2_2 ));
    InMux I__3370 (
            .O(N__17193),
            .I(N__17190));
    LocalMux I__3369 (
            .O(N__17190),
            .I(N__17187));
    Span4Mux_h I__3368 (
            .O(N__17187),
            .I(N__17184));
    Odrv4 I__3367 (
            .O(N__17184),
            .I(\Lab_UT.dictrl.N_19 ));
    CascadeMux I__3366 (
            .O(N__17181),
            .I(\Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_ ));
    InMux I__3365 (
            .O(N__17178),
            .I(N__17175));
    LocalMux I__3364 (
            .O(N__17175),
            .I(N__17172));
    Span4Mux_h I__3363 (
            .O(N__17172),
            .I(N__17169));
    Odrv4 I__3362 (
            .O(N__17169),
            .I(\Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3 ));
    InMux I__3361 (
            .O(N__17166),
            .I(N__17160));
    InMux I__3360 (
            .O(N__17165),
            .I(N__17160));
    LocalMux I__3359 (
            .O(N__17160),
            .I(N__17157));
    Span4Mux_h I__3358 (
            .O(N__17157),
            .I(N__17154));
    Odrv4 I__3357 (
            .O(N__17154),
            .I(\Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2 ));
    CascadeMux I__3356 (
            .O(N__17151),
            .I(\Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_ ));
    InMux I__3355 (
            .O(N__17148),
            .I(N__17133));
    InMux I__3354 (
            .O(N__17147),
            .I(N__17133));
    InMux I__3353 (
            .O(N__17146),
            .I(N__17133));
    InMux I__3352 (
            .O(N__17145),
            .I(N__17133));
    InMux I__3351 (
            .O(N__17144),
            .I(N__17133));
    LocalMux I__3350 (
            .O(N__17133),
            .I(N__17130));
    Odrv4 I__3349 (
            .O(N__17130),
            .I(\Lab_UT.dictrl.N_1792_0_0_0 ));
    InMux I__3348 (
            .O(N__17127),
            .I(N__17124));
    LocalMux I__3347 (
            .O(N__17124),
            .I(N__17121));
    Odrv4 I__3346 (
            .O(N__17121),
            .I(\Lab_UT.dictrl.m53_d_1_5 ));
    InMux I__3345 (
            .O(N__17118),
            .I(N__17114));
    InMux I__3344 (
            .O(N__17117),
            .I(N__17108));
    LocalMux I__3343 (
            .O(N__17114),
            .I(N__17104));
    InMux I__3342 (
            .O(N__17113),
            .I(N__17097));
    InMux I__3341 (
            .O(N__17112),
            .I(N__17097));
    InMux I__3340 (
            .O(N__17111),
            .I(N__17097));
    LocalMux I__3339 (
            .O(N__17108),
            .I(N__17090));
    InMux I__3338 (
            .O(N__17107),
            .I(N__17087));
    Span4Mux_v I__3337 (
            .O(N__17104),
            .I(N__17082));
    LocalMux I__3336 (
            .O(N__17097),
            .I(N__17082));
    InMux I__3335 (
            .O(N__17096),
            .I(N__17075));
    InMux I__3334 (
            .O(N__17095),
            .I(N__17075));
    InMux I__3333 (
            .O(N__17094),
            .I(N__17075));
    InMux I__3332 (
            .O(N__17093),
            .I(N__17072));
    Span4Mux_s3_h I__3331 (
            .O(N__17090),
            .I(N__17069));
    LocalMux I__3330 (
            .O(N__17087),
            .I(N__17066));
    Span4Mux_h I__3329 (
            .O(N__17082),
            .I(N__17061));
    LocalMux I__3328 (
            .O(N__17075),
            .I(N__17061));
    LocalMux I__3327 (
            .O(N__17072),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__3326 (
            .O(N__17069),
            .I(bu_rx_data_4_rep1));
    Odrv12 I__3325 (
            .O(N__17066),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__3324 (
            .O(N__17061),
            .I(bu_rx_data_4_rep1));
    InMux I__3323 (
            .O(N__17052),
            .I(N__17049));
    LocalMux I__3322 (
            .O(N__17049),
            .I(\Lab_UT.dictrl.N_40_0 ));
    CascadeMux I__3321 (
            .O(N__17046),
            .I(N__17042));
    CascadeMux I__3320 (
            .O(N__17045),
            .I(N__17038));
    InMux I__3319 (
            .O(N__17042),
            .I(N__17025));
    InMux I__3318 (
            .O(N__17041),
            .I(N__17025));
    InMux I__3317 (
            .O(N__17038),
            .I(N__17025));
    InMux I__3316 (
            .O(N__17037),
            .I(N__17025));
    InMux I__3315 (
            .O(N__17036),
            .I(N__17025));
    LocalMux I__3314 (
            .O(N__17025),
            .I(N__17022));
    Span4Mux_h I__3313 (
            .O(N__17022),
            .I(N__17019));
    Odrv4 I__3312 (
            .O(N__17019),
            .I(\Lab_UT.dictrl.N_23_1 ));
    InMux I__3311 (
            .O(N__17016),
            .I(N__17001));
    InMux I__3310 (
            .O(N__17015),
            .I(N__17001));
    InMux I__3309 (
            .O(N__17014),
            .I(N__17001));
    InMux I__3308 (
            .O(N__17013),
            .I(N__17001));
    InMux I__3307 (
            .O(N__17012),
            .I(N__17001));
    LocalMux I__3306 (
            .O(N__17001),
            .I(N__16998));
    Span4Mux_h I__3305 (
            .O(N__16998),
            .I(N__16995));
    Odrv4 I__3304 (
            .O(N__16995),
            .I(G_17_i_0));
    CascadeMux I__3303 (
            .O(N__16992),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ));
    CascadeMux I__3302 (
            .O(N__16989),
            .I(N__16984));
    CascadeMux I__3301 (
            .O(N__16988),
            .I(N__16980));
    InMux I__3300 (
            .O(N__16987),
            .I(N__16965));
    InMux I__3299 (
            .O(N__16984),
            .I(N__16965));
    InMux I__3298 (
            .O(N__16983),
            .I(N__16965));
    InMux I__3297 (
            .O(N__16980),
            .I(N__16965));
    InMux I__3296 (
            .O(N__16979),
            .I(N__16965));
    InMux I__3295 (
            .O(N__16978),
            .I(N__16965));
    LocalMux I__3294 (
            .O(N__16965),
            .I(N__16962));
    Odrv4 I__3293 (
            .O(N__16962),
            .I(\Lab_UT.dictrl.next_state_latmux_2_1 ));
    CascadeMux I__3292 (
            .O(N__16959),
            .I(N__16956));
    InMux I__3291 (
            .O(N__16956),
            .I(N__16952));
    InMux I__3290 (
            .O(N__16955),
            .I(N__16948));
    LocalMux I__3289 (
            .O(N__16952),
            .I(N__16945));
    IoInMux I__3288 (
            .O(N__16951),
            .I(N__16941));
    LocalMux I__3287 (
            .O(N__16948),
            .I(N__16938));
    Span4Mux_v I__3286 (
            .O(N__16945),
            .I(N__16935));
    SRMux I__3285 (
            .O(N__16944),
            .I(N__16932));
    LocalMux I__3284 (
            .O(N__16941),
            .I(N__16929));
    Span4Mux_v I__3283 (
            .O(N__16938),
            .I(N__16926));
    Span4Mux_v I__3282 (
            .O(N__16935),
            .I(N__16919));
    LocalMux I__3281 (
            .O(N__16932),
            .I(N__16919));
    Span4Mux_s1_v I__3280 (
            .O(N__16929),
            .I(N__16919));
    Span4Mux_v I__3279 (
            .O(N__16926),
            .I(N__16916));
    Span4Mux_h I__3278 (
            .O(N__16919),
            .I(N__16913));
    Odrv4 I__3277 (
            .O(N__16916),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3276 (
            .O(N__16913),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__3275 (
            .O(N__16908),
            .I(N__16905));
    InMux I__3274 (
            .O(N__16905),
            .I(N__16902));
    LocalMux I__3273 (
            .O(N__16902),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    CEMux I__3272 (
            .O(N__16899),
            .I(N__16896));
    LocalMux I__3271 (
            .O(N__16896),
            .I(N__16891));
    CEMux I__3270 (
            .O(N__16895),
            .I(N__16888));
    CEMux I__3269 (
            .O(N__16894),
            .I(N__16885));
    Span4Mux_s3_v I__3268 (
            .O(N__16891),
            .I(N__16881));
    LocalMux I__3267 (
            .O(N__16888),
            .I(N__16878));
    LocalMux I__3266 (
            .O(N__16885),
            .I(N__16875));
    CEMux I__3265 (
            .O(N__16884),
            .I(N__16872));
    Odrv4 I__3264 (
            .O(N__16881),
            .I(\Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ));
    Odrv12 I__3263 (
            .O(N__16878),
            .I(\Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ));
    Odrv4 I__3262 (
            .O(N__16875),
            .I(\Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ));
    LocalMux I__3261 (
            .O(N__16872),
            .I(\Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ));
    CascadeMux I__3260 (
            .O(N__16863),
            .I(N__16857));
    CascadeMux I__3259 (
            .O(N__16862),
            .I(N__16853));
    CascadeMux I__3258 (
            .O(N__16861),
            .I(N__16850));
    InMux I__3257 (
            .O(N__16860),
            .I(N__16839));
    InMux I__3256 (
            .O(N__16857),
            .I(N__16839));
    InMux I__3255 (
            .O(N__16856),
            .I(N__16839));
    InMux I__3254 (
            .O(N__16853),
            .I(N__16839));
    InMux I__3253 (
            .O(N__16850),
            .I(N__16839));
    LocalMux I__3252 (
            .O(N__16839),
            .I(\Lab_UT.dictrl.G_17_i_a5_1_1 ));
    InMux I__3251 (
            .O(N__16836),
            .I(N__16822));
    InMux I__3250 (
            .O(N__16835),
            .I(N__16822));
    InMux I__3249 (
            .O(N__16834),
            .I(N__16822));
    InMux I__3248 (
            .O(N__16833),
            .I(N__16819));
    InMux I__3247 (
            .O(N__16832),
            .I(N__16812));
    InMux I__3246 (
            .O(N__16831),
            .I(N__16812));
    InMux I__3245 (
            .O(N__16830),
            .I(N__16812));
    InMux I__3244 (
            .O(N__16829),
            .I(N__16809));
    LocalMux I__3243 (
            .O(N__16822),
            .I(N__16806));
    LocalMux I__3242 (
            .O(N__16819),
            .I(N__16801));
    LocalMux I__3241 (
            .O(N__16812),
            .I(N__16801));
    LocalMux I__3240 (
            .O(N__16809),
            .I(N__16798));
    Span4Mux_v I__3239 (
            .O(N__16806),
            .I(N__16792));
    Span4Mux_v I__3238 (
            .O(N__16801),
            .I(N__16789));
    Span4Mux_h I__3237 (
            .O(N__16798),
            .I(N__16786));
    InMux I__3236 (
            .O(N__16797),
            .I(N__16779));
    InMux I__3235 (
            .O(N__16796),
            .I(N__16779));
    InMux I__3234 (
            .O(N__16795),
            .I(N__16779));
    Odrv4 I__3233 (
            .O(N__16792),
            .I(\Lab_UT.dictrl.state_1_rep2 ));
    Odrv4 I__3232 (
            .O(N__16789),
            .I(\Lab_UT.dictrl.state_1_rep2 ));
    Odrv4 I__3231 (
            .O(N__16786),
            .I(\Lab_UT.dictrl.state_1_rep2 ));
    LocalMux I__3230 (
            .O(N__16779),
            .I(\Lab_UT.dictrl.state_1_rep2 ));
    InMux I__3229 (
            .O(N__16770),
            .I(N__16767));
    LocalMux I__3228 (
            .O(N__16767),
            .I(N__16764));
    Odrv12 I__3227 (
            .O(N__16764),
            .I(\Lab_UT.dictrl.N_15_0 ));
    InMux I__3226 (
            .O(N__16761),
            .I(N__16758));
    LocalMux I__3225 (
            .O(N__16758),
            .I(N__16755));
    Span4Mux_h I__3224 (
            .O(N__16755),
            .I(N__16752));
    Odrv4 I__3223 (
            .O(N__16752),
            .I(\Lab_UT.dictrl.g0_i_m2_0_1 ));
    CascadeMux I__3222 (
            .O(N__16749),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_ ));
    InMux I__3221 (
            .O(N__16746),
            .I(N__16743));
    LocalMux I__3220 (
            .O(N__16743),
            .I(N__16740));
    Odrv4 I__3219 (
            .O(N__16740),
            .I(\Lab_UT.dictrl.g0_i_m2_0_2 ));
    CascadeMux I__3218 (
            .O(N__16737),
            .I(\Lab_UT.dictrl.next_state_0_0_2_cascade_ ));
    InMux I__3217 (
            .O(N__16734),
            .I(N__16730));
    InMux I__3216 (
            .O(N__16733),
            .I(N__16727));
    LocalMux I__3215 (
            .O(N__16730),
            .I(N__16721));
    LocalMux I__3214 (
            .O(N__16727),
            .I(N__16721));
    InMux I__3213 (
            .O(N__16726),
            .I(N__16716));
    Span4Mux_h I__3212 (
            .O(N__16721),
            .I(N__16713));
    InMux I__3211 (
            .O(N__16720),
            .I(N__16710));
    InMux I__3210 (
            .O(N__16719),
            .I(N__16707));
    LocalMux I__3209 (
            .O(N__16716),
            .I(N__16704));
    Span4Mux_v I__3208 (
            .O(N__16713),
            .I(N__16697));
    LocalMux I__3207 (
            .O(N__16710),
            .I(N__16697));
    LocalMux I__3206 (
            .O(N__16707),
            .I(N__16697));
    Span4Mux_s3_v I__3205 (
            .O(N__16704),
            .I(N__16694));
    Span4Mux_h I__3204 (
            .O(N__16697),
            .I(N__16690));
    Span4Mux_h I__3203 (
            .O(N__16694),
            .I(N__16687));
    IoInMux I__3202 (
            .O(N__16693),
            .I(N__16684));
    Odrv4 I__3201 (
            .O(N__16690),
            .I(rst));
    Odrv4 I__3200 (
            .O(N__16687),
            .I(rst));
    LocalMux I__3199 (
            .O(N__16684),
            .I(rst));
    CascadeMux I__3198 (
            .O(N__16677),
            .I(N__16674));
    InMux I__3197 (
            .O(N__16674),
            .I(N__16671));
    LocalMux I__3196 (
            .O(N__16671),
            .I(N__16668));
    Odrv4 I__3195 (
            .O(N__16668),
            .I(\Lab_UT.didp.countrce4.un13_qPone ));
    InMux I__3194 (
            .O(N__16665),
            .I(N__16662));
    LocalMux I__3193 (
            .O(N__16662),
            .I(N__16659));
    Span4Mux_v I__3192 (
            .O(N__16659),
            .I(N__16656));
    Span4Mux_h I__3191 (
            .O(N__16656),
            .I(N__16652));
    InMux I__3190 (
            .O(N__16655),
            .I(N__16649));
    Odrv4 I__3189 (
            .O(N__16652),
            .I(\Lab_UT.LdAMtens ));
    LocalMux I__3188 (
            .O(N__16649),
            .I(\Lab_UT.LdAMtens ));
    InMux I__3187 (
            .O(N__16644),
            .I(N__16638));
    InMux I__3186 (
            .O(N__16643),
            .I(N__16638));
    LocalMux I__3185 (
            .O(N__16638),
            .I(\Lab_UT.LdAMones ));
    InMux I__3184 (
            .O(N__16635),
            .I(N__16632));
    LocalMux I__3183 (
            .O(N__16632),
            .I(N__16629));
    Span4Mux_s3_h I__3182 (
            .O(N__16629),
            .I(N__16625));
    CascadeMux I__3181 (
            .O(N__16628),
            .I(N__16622));
    Span4Mux_h I__3180 (
            .O(N__16625),
            .I(N__16619));
    InMux I__3179 (
            .O(N__16622),
            .I(N__16616));
    Odrv4 I__3178 (
            .O(N__16619),
            .I(\Lab_UT.LdAStens ));
    LocalMux I__3177 (
            .O(N__16616),
            .I(\Lab_UT.LdAStens ));
    InMux I__3176 (
            .O(N__16611),
            .I(N__16608));
    LocalMux I__3175 (
            .O(N__16608),
            .I(N__16605));
    Odrv4 I__3174 (
            .O(N__16605),
            .I(\Lab_UT.dictrl.N_1460_2 ));
    InMux I__3173 (
            .O(N__16602),
            .I(N__16594));
    InMux I__3172 (
            .O(N__16601),
            .I(N__16594));
    InMux I__3171 (
            .O(N__16600),
            .I(N__16589));
    InMux I__3170 (
            .O(N__16599),
            .I(N__16586));
    LocalMux I__3169 (
            .O(N__16594),
            .I(N__16583));
    InMux I__3168 (
            .O(N__16593),
            .I(N__16578));
    InMux I__3167 (
            .O(N__16592),
            .I(N__16578));
    LocalMux I__3166 (
            .O(N__16589),
            .I(N__16575));
    LocalMux I__3165 (
            .O(N__16586),
            .I(N__16570));
    Span4Mux_s2_v I__3164 (
            .O(N__16583),
            .I(N__16570));
    LocalMux I__3163 (
            .O(N__16578),
            .I(N__16567));
    Span4Mux_v I__3162 (
            .O(N__16575),
            .I(N__16562));
    Span4Mux_v I__3161 (
            .O(N__16570),
            .I(N__16562));
    Odrv12 I__3160 (
            .O(N__16567),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    Odrv4 I__3159 (
            .O(N__16562),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    InMux I__3158 (
            .O(N__16557),
            .I(N__16554));
    LocalMux I__3157 (
            .O(N__16554),
            .I(N__16551));
    Odrv4 I__3156 (
            .O(N__16551),
            .I(\Lab_UT.dispString.m49Z0Z_0 ));
    InMux I__3155 (
            .O(N__16548),
            .I(N__16545));
    LocalMux I__3154 (
            .O(N__16545),
            .I(\Lab_UT.dispString.m49Z0Z_1 ));
    CascadeMux I__3153 (
            .O(N__16542),
            .I(\Lab_UT.dispString.m49Z0Z_3_cascade_ ));
    CascadeMux I__3152 (
            .O(N__16539),
            .I(\Lab_UT.loadalarm_0_cascade_ ));
    InMux I__3151 (
            .O(N__16536),
            .I(N__16517));
    InMux I__3150 (
            .O(N__16535),
            .I(N__16517));
    InMux I__3149 (
            .O(N__16534),
            .I(N__16517));
    InMux I__3148 (
            .O(N__16533),
            .I(N__16517));
    InMux I__3147 (
            .O(N__16532),
            .I(N__16517));
    InMux I__3146 (
            .O(N__16531),
            .I(N__16517));
    InMux I__3145 (
            .O(N__16530),
            .I(N__16514));
    LocalMux I__3144 (
            .O(N__16517),
            .I(N__16511));
    LocalMux I__3143 (
            .O(N__16514),
            .I(N__16508));
    Span4Mux_v I__3142 (
            .O(N__16511),
            .I(N__16505));
    Odrv12 I__3141 (
            .O(N__16508),
            .I(\Lab_UT.min2_0 ));
    Odrv4 I__3140 (
            .O(N__16505),
            .I(\Lab_UT.min2_0 ));
    CascadeMux I__3139 (
            .O(N__16500),
            .I(N__16497));
    InMux I__3138 (
            .O(N__16497),
            .I(N__16494));
    LocalMux I__3137 (
            .O(N__16494),
            .I(N__16491));
    Span4Mux_h I__3136 (
            .O(N__16491),
            .I(N__16486));
    InMux I__3135 (
            .O(N__16490),
            .I(N__16481));
    InMux I__3134 (
            .O(N__16489),
            .I(N__16481));
    Odrv4 I__3133 (
            .O(N__16486),
            .I(\Lab_UT.di_AMones_0 ));
    LocalMux I__3132 (
            .O(N__16481),
            .I(\Lab_UT.di_AMones_0 ));
    CascadeMux I__3131 (
            .O(N__16476),
            .I(N__16472));
    InMux I__3130 (
            .O(N__16475),
            .I(N__16468));
    InMux I__3129 (
            .O(N__16472),
            .I(N__16465));
    InMux I__3128 (
            .O(N__16471),
            .I(N__16462));
    LocalMux I__3127 (
            .O(N__16468),
            .I(N__16457));
    LocalMux I__3126 (
            .O(N__16465),
            .I(N__16457));
    LocalMux I__3125 (
            .O(N__16462),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__3124 (
            .O(N__16457),
            .I(\Lab_UT.di_AMtens_0 ));
    CascadeMux I__3123 (
            .O(N__16452),
            .I(\Lab_UT.dictrl.g0_12_a6_1_3_cascade_ ));
    InMux I__3122 (
            .O(N__16449),
            .I(N__16446));
    LocalMux I__3121 (
            .O(N__16446),
            .I(N__16443));
    Odrv4 I__3120 (
            .O(N__16443),
            .I(\Lab_UT.dictrl.N_18 ));
    CascadeMux I__3119 (
            .O(N__16440),
            .I(N__16437));
    InMux I__3118 (
            .O(N__16437),
            .I(N__16434));
    LocalMux I__3117 (
            .O(N__16434),
            .I(N__16431));
    Span4Mux_v I__3116 (
            .O(N__16431),
            .I(N__16428));
    Odrv4 I__3115 (
            .O(N__16428),
            .I(\Lab_UT.dictrl.m35_0 ));
    InMux I__3114 (
            .O(N__16425),
            .I(N__16419));
    CascadeMux I__3113 (
            .O(N__16424),
            .I(N__16415));
    CascadeMux I__3112 (
            .O(N__16423),
            .I(N__16412));
    CascadeMux I__3111 (
            .O(N__16422),
            .I(N__16409));
    LocalMux I__3110 (
            .O(N__16419),
            .I(N__16404));
    InMux I__3109 (
            .O(N__16418),
            .I(N__16391));
    InMux I__3108 (
            .O(N__16415),
            .I(N__16391));
    InMux I__3107 (
            .O(N__16412),
            .I(N__16391));
    InMux I__3106 (
            .O(N__16409),
            .I(N__16391));
    InMux I__3105 (
            .O(N__16408),
            .I(N__16391));
    InMux I__3104 (
            .O(N__16407),
            .I(N__16391));
    Span4Mux_s1_v I__3103 (
            .O(N__16404),
            .I(N__16386));
    LocalMux I__3102 (
            .O(N__16391),
            .I(N__16386));
    Odrv4 I__3101 (
            .O(N__16386),
            .I(\Lab_UT.min2_1 ));
    InMux I__3100 (
            .O(N__16383),
            .I(N__16380));
    LocalMux I__3099 (
            .O(N__16380),
            .I(N__16371));
    InMux I__3098 (
            .O(N__16379),
            .I(N__16358));
    InMux I__3097 (
            .O(N__16378),
            .I(N__16358));
    InMux I__3096 (
            .O(N__16377),
            .I(N__16358));
    InMux I__3095 (
            .O(N__16376),
            .I(N__16358));
    InMux I__3094 (
            .O(N__16375),
            .I(N__16358));
    InMux I__3093 (
            .O(N__16374),
            .I(N__16358));
    Span4Mux_h I__3092 (
            .O(N__16371),
            .I(N__16353));
    LocalMux I__3091 (
            .O(N__16358),
            .I(N__16353));
    Span4Mux_v I__3090 (
            .O(N__16353),
            .I(N__16350));
    Odrv4 I__3089 (
            .O(N__16350),
            .I(\Lab_UT.min2_2 ));
    CascadeMux I__3088 (
            .O(N__16347),
            .I(N__16344));
    InMux I__3087 (
            .O(N__16344),
            .I(N__16341));
    LocalMux I__3086 (
            .O(N__16341),
            .I(N__16338));
    Span4Mux_h I__3085 (
            .O(N__16338),
            .I(N__16333));
    InMux I__3084 (
            .O(N__16337),
            .I(N__16328));
    InMux I__3083 (
            .O(N__16336),
            .I(N__16328));
    Odrv4 I__3082 (
            .O(N__16333),
            .I(\Lab_UT.di_AStens_3 ));
    LocalMux I__3081 (
            .O(N__16328),
            .I(\Lab_UT.di_AStens_3 ));
    CEMux I__3080 (
            .O(N__16323),
            .I(N__16320));
    LocalMux I__3079 (
            .O(N__16320),
            .I(N__16317));
    Span4Mux_h I__3078 (
            .O(N__16317),
            .I(N__16314));
    Odrv4 I__3077 (
            .O(N__16314),
            .I(\Lab_UT.didp.regrce2.LdAStens_0 ));
    CascadeMux I__3076 (
            .O(N__16311),
            .I(\Lab_UT.didp.countrce4.q_5_2_cascade_ ));
    InMux I__3075 (
            .O(N__16308),
            .I(N__16304));
    InMux I__3074 (
            .O(N__16307),
            .I(N__16300));
    LocalMux I__3073 (
            .O(N__16304),
            .I(N__16297));
    InMux I__3072 (
            .O(N__16303),
            .I(N__16294));
    LocalMux I__3071 (
            .O(N__16300),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__3070 (
            .O(N__16297),
            .I(\Lab_UT.di_AMtens_2 ));
    LocalMux I__3069 (
            .O(N__16294),
            .I(\Lab_UT.di_AMtens_2 ));
    InMux I__3068 (
            .O(N__16287),
            .I(N__16283));
    CascadeMux I__3067 (
            .O(N__16286),
            .I(N__16279));
    LocalMux I__3066 (
            .O(N__16283),
            .I(N__16276));
    InMux I__3065 (
            .O(N__16282),
            .I(N__16273));
    InMux I__3064 (
            .O(N__16279),
            .I(N__16270));
    Span4Mux_v I__3063 (
            .O(N__16276),
            .I(N__16267));
    LocalMux I__3062 (
            .O(N__16273),
            .I(N__16264));
    LocalMux I__3061 (
            .O(N__16270),
            .I(N__16261));
    Odrv4 I__3060 (
            .O(N__16267),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv4 I__3059 (
            .O(N__16264),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv4 I__3058 (
            .O(N__16261),
            .I(\Lab_UT.di_AMtens_1 ));
    InMux I__3057 (
            .O(N__16254),
            .I(N__16246));
    CascadeMux I__3056 (
            .O(N__16253),
            .I(N__16243));
    InMux I__3055 (
            .O(N__16252),
            .I(N__16235));
    InMux I__3054 (
            .O(N__16251),
            .I(N__16232));
    InMux I__3053 (
            .O(N__16250),
            .I(N__16229));
    InMux I__3052 (
            .O(N__16249),
            .I(N__16226));
    LocalMux I__3051 (
            .O(N__16246),
            .I(N__16223));
    InMux I__3050 (
            .O(N__16243),
            .I(N__16214));
    InMux I__3049 (
            .O(N__16242),
            .I(N__16214));
    InMux I__3048 (
            .O(N__16241),
            .I(N__16214));
    InMux I__3047 (
            .O(N__16240),
            .I(N__16214));
    InMux I__3046 (
            .O(N__16239),
            .I(N__16209));
    InMux I__3045 (
            .O(N__16238),
            .I(N__16209));
    LocalMux I__3044 (
            .O(N__16235),
            .I(N__16198));
    LocalMux I__3043 (
            .O(N__16232),
            .I(N__16198));
    LocalMux I__3042 (
            .O(N__16229),
            .I(N__16198));
    LocalMux I__3041 (
            .O(N__16226),
            .I(N__16198));
    Span12Mux_s11_h I__3040 (
            .O(N__16223),
            .I(N__16198));
    LocalMux I__3039 (
            .O(N__16214),
            .I(buart__rx_startbit));
    LocalMux I__3038 (
            .O(N__16209),
            .I(buart__rx_startbit));
    Odrv12 I__3037 (
            .O(N__16198),
            .I(buart__rx_startbit));
    InMux I__3036 (
            .O(N__16191),
            .I(N__16188));
    LocalMux I__3035 (
            .O(N__16188),
            .I(N__16185));
    Span4Mux_h I__3034 (
            .O(N__16185),
            .I(N__16182));
    Span4Mux_v I__3033 (
            .O(N__16182),
            .I(N__16178));
    InMux I__3032 (
            .O(N__16181),
            .I(N__16175));
    Span4Mux_h I__3031 (
            .O(N__16178),
            .I(N__16170));
    LocalMux I__3030 (
            .O(N__16175),
            .I(N__16167));
    InMux I__3029 (
            .O(N__16174),
            .I(N__16164));
    InMux I__3028 (
            .O(N__16173),
            .I(N__16161));
    Odrv4 I__3027 (
            .O(N__16170),
            .I(buart__rx_N_27_0_i));
    Odrv4 I__3026 (
            .O(N__16167),
            .I(buart__rx_N_27_0_i));
    LocalMux I__3025 (
            .O(N__16164),
            .I(buart__rx_N_27_0_i));
    LocalMux I__3024 (
            .O(N__16161),
            .I(buart__rx_N_27_0_i));
    CascadeMux I__3023 (
            .O(N__16152),
            .I(N__16149));
    InMux I__3022 (
            .O(N__16149),
            .I(N__16146));
    LocalMux I__3021 (
            .O(N__16146),
            .I(N__16143));
    Span4Mux_h I__3020 (
            .O(N__16143),
            .I(N__16140));
    Span4Mux_v I__3019 (
            .O(N__16140),
            .I(N__16137));
    Span4Mux_h I__3018 (
            .O(N__16137),
            .I(N__16134));
    Odrv4 I__3017 (
            .O(N__16134),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__3016 (
            .O(N__16131),
            .I(N__16125));
    InMux I__3015 (
            .O(N__16130),
            .I(N__16122));
    InMux I__3014 (
            .O(N__16129),
            .I(N__16117));
    InMux I__3013 (
            .O(N__16128),
            .I(N__16117));
    LocalMux I__3012 (
            .O(N__16125),
            .I(N__16114));
    LocalMux I__3011 (
            .O(N__16122),
            .I(N__16109));
    LocalMux I__3010 (
            .O(N__16117),
            .I(N__16109));
    Span4Mux_v I__3009 (
            .O(N__16114),
            .I(N__16104));
    Span4Mux_v I__3008 (
            .O(N__16109),
            .I(N__16104));
    Span4Mux_h I__3007 (
            .O(N__16104),
            .I(N__16100));
    InMux I__3006 (
            .O(N__16103),
            .I(N__16097));
    Span4Mux_v I__3005 (
            .O(N__16100),
            .I(N__16094));
    LocalMux I__3004 (
            .O(N__16097),
            .I(buart__rx_bitcount_2));
    Odrv4 I__3003 (
            .O(N__16094),
            .I(buart__rx_bitcount_2));
    CEMux I__3002 (
            .O(N__16089),
            .I(N__16086));
    LocalMux I__3001 (
            .O(N__16086),
            .I(N__16082));
    CEMux I__3000 (
            .O(N__16085),
            .I(N__16078));
    Sp12to4 I__2999 (
            .O(N__16082),
            .I(N__16074));
    CEMux I__2998 (
            .O(N__16081),
            .I(N__16071));
    LocalMux I__2997 (
            .O(N__16078),
            .I(N__16068));
    CEMux I__2996 (
            .O(N__16077),
            .I(N__16065));
    Span12Mux_s9_v I__2995 (
            .O(N__16074),
            .I(N__16062));
    LocalMux I__2994 (
            .O(N__16071),
            .I(N__16059));
    Span4Mux_v I__2993 (
            .O(N__16068),
            .I(N__16056));
    LocalMux I__2992 (
            .O(N__16065),
            .I(N__16053));
    Odrv12 I__2991 (
            .O(N__16062),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__2990 (
            .O(N__16059),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__2989 (
            .O(N__16056),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__2988 (
            .O(N__16053),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__2987 (
            .O(N__16044),
            .I(N__16041));
    LocalMux I__2986 (
            .O(N__16041),
            .I(\uu2.bitmapZ0Z_75 ));
    InMux I__2985 (
            .O(N__16038),
            .I(N__16035));
    LocalMux I__2984 (
            .O(N__16035),
            .I(\uu2.bitmapZ0Z_72 ));
    InMux I__2983 (
            .O(N__16032),
            .I(N__16029));
    LocalMux I__2982 (
            .O(N__16029),
            .I(N__16026));
    Odrv4 I__2981 (
            .O(N__16026),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__2980 (
            .O(N__16023),
            .I(N__16019));
    InMux I__2979 (
            .O(N__16022),
            .I(N__16016));
    LocalMux I__2978 (
            .O(N__16019),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    LocalMux I__2977 (
            .O(N__16016),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    CEMux I__2976 (
            .O(N__16011),
            .I(N__16008));
    LocalMux I__2975 (
            .O(N__16008),
            .I(N__16005));
    Span4Mux_s3_h I__2974 (
            .O(N__16005),
            .I(N__16002));
    Span4Mux_h I__2973 (
            .O(N__16002),
            .I(N__15999));
    Odrv4 I__2972 (
            .O(N__15999),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    InMux I__2971 (
            .O(N__15996),
            .I(N__15993));
    LocalMux I__2970 (
            .O(N__15993),
            .I(N__15990));
    Span4Mux_h I__2969 (
            .O(N__15990),
            .I(N__15985));
    InMux I__2968 (
            .O(N__15989),
            .I(N__15980));
    InMux I__2967 (
            .O(N__15988),
            .I(N__15980));
    Odrv4 I__2966 (
            .O(N__15985),
            .I(\Lab_UT.di_ASones_3 ));
    LocalMux I__2965 (
            .O(N__15980),
            .I(\Lab_UT.di_ASones_3 ));
    CascadeMux I__2964 (
            .O(N__15975),
            .I(\uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_ ));
    InMux I__2963 (
            .O(N__15972),
            .I(N__15968));
    CascadeMux I__2962 (
            .O(N__15971),
            .I(N__15965));
    LocalMux I__2961 (
            .O(N__15968),
            .I(N__15957));
    InMux I__2960 (
            .O(N__15965),
            .I(N__15950));
    InMux I__2959 (
            .O(N__15964),
            .I(N__15950));
    InMux I__2958 (
            .O(N__15963),
            .I(N__15950));
    InMux I__2957 (
            .O(N__15962),
            .I(N__15943));
    InMux I__2956 (
            .O(N__15961),
            .I(N__15943));
    InMux I__2955 (
            .O(N__15960),
            .I(N__15943));
    Span4Mux_s3_v I__2954 (
            .O(N__15957),
            .I(N__15940));
    LocalMux I__2953 (
            .O(N__15950),
            .I(N__15935));
    LocalMux I__2952 (
            .O(N__15943),
            .I(N__15935));
    Odrv4 I__2951 (
            .O(N__15940),
            .I(\Lab_UT.min1_2 ));
    Odrv12 I__2950 (
            .O(N__15935),
            .I(\Lab_UT.min1_2 ));
    InMux I__2949 (
            .O(N__15930),
            .I(N__15926));
    CascadeMux I__2948 (
            .O(N__15929),
            .I(N__15919));
    LocalMux I__2947 (
            .O(N__15926),
            .I(N__15915));
    InMux I__2946 (
            .O(N__15925),
            .I(N__15908));
    InMux I__2945 (
            .O(N__15924),
            .I(N__15908));
    InMux I__2944 (
            .O(N__15923),
            .I(N__15908));
    InMux I__2943 (
            .O(N__15922),
            .I(N__15901));
    InMux I__2942 (
            .O(N__15919),
            .I(N__15901));
    InMux I__2941 (
            .O(N__15918),
            .I(N__15901));
    Span4Mux_v I__2940 (
            .O(N__15915),
            .I(N__15898));
    LocalMux I__2939 (
            .O(N__15908),
            .I(N__15895));
    LocalMux I__2938 (
            .O(N__15901),
            .I(N__15892));
    Odrv4 I__2937 (
            .O(N__15898),
            .I(\Lab_UT.min1_1 ));
    Odrv12 I__2936 (
            .O(N__15895),
            .I(\Lab_UT.min1_1 ));
    Odrv4 I__2935 (
            .O(N__15892),
            .I(\Lab_UT.min1_1 ));
    CascadeMux I__2934 (
            .O(N__15885),
            .I(N__15882));
    InMux I__2933 (
            .O(N__15882),
            .I(N__15875));
    CascadeMux I__2932 (
            .O(N__15881),
            .I(N__15871));
    CascadeMux I__2931 (
            .O(N__15880),
            .I(N__15868));
    CascadeMux I__2930 (
            .O(N__15879),
            .I(N__15865));
    CascadeMux I__2929 (
            .O(N__15878),
            .I(N__15861));
    LocalMux I__2928 (
            .O(N__15875),
            .I(N__15858));
    InMux I__2927 (
            .O(N__15874),
            .I(N__15851));
    InMux I__2926 (
            .O(N__15871),
            .I(N__15851));
    InMux I__2925 (
            .O(N__15868),
            .I(N__15851));
    InMux I__2924 (
            .O(N__15865),
            .I(N__15844));
    InMux I__2923 (
            .O(N__15864),
            .I(N__15844));
    InMux I__2922 (
            .O(N__15861),
            .I(N__15844));
    Span4Mux_h I__2921 (
            .O(N__15858),
            .I(N__15839));
    LocalMux I__2920 (
            .O(N__15851),
            .I(N__15839));
    LocalMux I__2919 (
            .O(N__15844),
            .I(N__15836));
    Odrv4 I__2918 (
            .O(N__15839),
            .I(\Lab_UT.min1_3 ));
    Odrv4 I__2917 (
            .O(N__15836),
            .I(\Lab_UT.min1_3 ));
    InMux I__2916 (
            .O(N__15831),
            .I(N__15828));
    LocalMux I__2915 (
            .O(N__15828),
            .I(N__15819));
    InMux I__2914 (
            .O(N__15827),
            .I(N__15812));
    InMux I__2913 (
            .O(N__15826),
            .I(N__15812));
    InMux I__2912 (
            .O(N__15825),
            .I(N__15812));
    InMux I__2911 (
            .O(N__15824),
            .I(N__15805));
    InMux I__2910 (
            .O(N__15823),
            .I(N__15805));
    InMux I__2909 (
            .O(N__15822),
            .I(N__15805));
    Span4Mux_s3_v I__2908 (
            .O(N__15819),
            .I(N__15802));
    LocalMux I__2907 (
            .O(N__15812),
            .I(N__15799));
    LocalMux I__2906 (
            .O(N__15805),
            .I(N__15796));
    Odrv4 I__2905 (
            .O(N__15802),
            .I(\Lab_UT.min1_0 ));
    Odrv12 I__2904 (
            .O(N__15799),
            .I(\Lab_UT.min1_0 ));
    Odrv4 I__2903 (
            .O(N__15796),
            .I(\Lab_UT.min1_0 ));
    InMux I__2902 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__2901 (
            .O(N__15786),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__2900 (
            .O(N__15783),
            .I(N__15780));
    LocalMux I__2899 (
            .O(N__15780),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__2898 (
            .O(N__15777),
            .I(N__15757));
    InMux I__2897 (
            .O(N__15776),
            .I(N__15757));
    InMux I__2896 (
            .O(N__15775),
            .I(N__15757));
    InMux I__2895 (
            .O(N__15774),
            .I(N__15757));
    InMux I__2894 (
            .O(N__15773),
            .I(N__15757));
    InMux I__2893 (
            .O(N__15772),
            .I(N__15750));
    InMux I__2892 (
            .O(N__15771),
            .I(N__15750));
    InMux I__2891 (
            .O(N__15770),
            .I(N__15750));
    InMux I__2890 (
            .O(N__15769),
            .I(N__15745));
    InMux I__2889 (
            .O(N__15768),
            .I(N__15745));
    LocalMux I__2888 (
            .O(N__15757),
            .I(N__15742));
    LocalMux I__2887 (
            .O(N__15750),
            .I(N__15737));
    LocalMux I__2886 (
            .O(N__15745),
            .I(N__15737));
    Odrv4 I__2885 (
            .O(N__15742),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__2884 (
            .O(N__15737),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    InMux I__2883 (
            .O(N__15732),
            .I(N__15729));
    LocalMux I__2882 (
            .O(N__15729),
            .I(\uu2.bitmap_pmux_sn_N_65 ));
    InMux I__2881 (
            .O(N__15726),
            .I(N__15723));
    LocalMux I__2880 (
            .O(N__15723),
            .I(\uu2.N_54 ));
    InMux I__2879 (
            .O(N__15720),
            .I(N__15717));
    LocalMux I__2878 (
            .O(N__15717),
            .I(\uu2.N_53 ));
    InMux I__2877 (
            .O(N__15714),
            .I(N__15711));
    LocalMux I__2876 (
            .O(N__15711),
            .I(N__15708));
    Odrv4 I__2875 (
            .O(N__15708),
            .I(\Lab_UT.dictrl.m53_d_1_3 ));
    CascadeMux I__2874 (
            .O(N__15705),
            .I(\Lab_UT.dictrl.N_97_mux_5_cascade_ ));
    InMux I__2873 (
            .O(N__15702),
            .I(N__15697));
    InMux I__2872 (
            .O(N__15701),
            .I(N__15694));
    CascadeMux I__2871 (
            .O(N__15700),
            .I(N__15689));
    LocalMux I__2870 (
            .O(N__15697),
            .I(N__15684));
    LocalMux I__2869 (
            .O(N__15694),
            .I(N__15684));
    InMux I__2868 (
            .O(N__15693),
            .I(N__15681));
    InMux I__2867 (
            .O(N__15692),
            .I(N__15676));
    InMux I__2866 (
            .O(N__15689),
            .I(N__15676));
    Span4Mux_s1_v I__2865 (
            .O(N__15684),
            .I(N__15673));
    LocalMux I__2864 (
            .O(N__15681),
            .I(\Lab_UT.dictrl.N_40 ));
    LocalMux I__2863 (
            .O(N__15676),
            .I(\Lab_UT.dictrl.N_40 ));
    Odrv4 I__2862 (
            .O(N__15673),
            .I(\Lab_UT.dictrl.N_40 ));
    InMux I__2861 (
            .O(N__15666),
            .I(N__15662));
    InMux I__2860 (
            .O(N__15665),
            .I(N__15659));
    LocalMux I__2859 (
            .O(N__15662),
            .I(N__15656));
    LocalMux I__2858 (
            .O(N__15659),
            .I(\Lab_UT.dictrl.N_62 ));
    Odrv12 I__2857 (
            .O(N__15656),
            .I(\Lab_UT.dictrl.N_62 ));
    CascadeMux I__2856 (
            .O(N__15651),
            .I(\Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_ ));
    InMux I__2855 (
            .O(N__15648),
            .I(N__15645));
    LocalMux I__2854 (
            .O(N__15645),
            .I(\Lab_UT.dictrl.next_state_RNO_1Z0Z_2 ));
    InMux I__2853 (
            .O(N__15642),
            .I(N__15639));
    LocalMux I__2852 (
            .O(N__15639),
            .I(\Lab_UT.dictrl.next_state_RNO_0Z0Z_2 ));
    InMux I__2851 (
            .O(N__15636),
            .I(N__15633));
    LocalMux I__2850 (
            .O(N__15633),
            .I(N__15620));
    InMux I__2849 (
            .O(N__15632),
            .I(N__15615));
    InMux I__2848 (
            .O(N__15631),
            .I(N__15615));
    InMux I__2847 (
            .O(N__15630),
            .I(N__15608));
    InMux I__2846 (
            .O(N__15629),
            .I(N__15608));
    InMux I__2845 (
            .O(N__15628),
            .I(N__15608));
    InMux I__2844 (
            .O(N__15627),
            .I(N__15603));
    InMux I__2843 (
            .O(N__15626),
            .I(N__15598));
    InMux I__2842 (
            .O(N__15625),
            .I(N__15598));
    InMux I__2841 (
            .O(N__15624),
            .I(N__15595));
    InMux I__2840 (
            .O(N__15623),
            .I(N__15592));
    Span4Mux_h I__2839 (
            .O(N__15620),
            .I(N__15587));
    LocalMux I__2838 (
            .O(N__15615),
            .I(N__15587));
    LocalMux I__2837 (
            .O(N__15608),
            .I(N__15584));
    InMux I__2836 (
            .O(N__15607),
            .I(N__15581));
    InMux I__2835 (
            .O(N__15606),
            .I(N__15578));
    LocalMux I__2834 (
            .O(N__15603),
            .I(N__15575));
    LocalMux I__2833 (
            .O(N__15598),
            .I(N__15564));
    LocalMux I__2832 (
            .O(N__15595),
            .I(N__15564));
    LocalMux I__2831 (
            .O(N__15592),
            .I(N__15564));
    Sp12to4 I__2830 (
            .O(N__15587),
            .I(N__15564));
    Sp12to4 I__2829 (
            .O(N__15584),
            .I(N__15564));
    LocalMux I__2828 (
            .O(N__15581),
            .I(N__15561));
    LocalMux I__2827 (
            .O(N__15578),
            .I(N__15558));
    Span12Mux_s5_h I__2826 (
            .O(N__15575),
            .I(N__15553));
    Span12Mux_s6_v I__2825 (
            .O(N__15564),
            .I(N__15553));
    Span4Mux_s3_v I__2824 (
            .O(N__15561),
            .I(N__15548));
    Span4Mux_h I__2823 (
            .O(N__15558),
            .I(N__15548));
    Odrv12 I__2822 (
            .O(N__15553),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    Odrv4 I__2821 (
            .O(N__15548),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    InMux I__2820 (
            .O(N__15543),
            .I(N__15540));
    LocalMux I__2819 (
            .O(N__15540),
            .I(N__15536));
    InMux I__2818 (
            .O(N__15539),
            .I(N__15533));
    Odrv4 I__2817 (
            .O(N__15536),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    LocalMux I__2816 (
            .O(N__15533),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    InMux I__2815 (
            .O(N__15528),
            .I(N__15525));
    LocalMux I__2814 (
            .O(N__15525),
            .I(N__15522));
    Span4Mux_h I__2813 (
            .O(N__15522),
            .I(N__15519));
    Odrv4 I__2812 (
            .O(N__15519),
            .I(\Lab_UT.dictrl.next_state_RNINV3PZ0Z_2 ));
    CascadeMux I__2811 (
            .O(N__15516),
            .I(N__15510));
    CascadeMux I__2810 (
            .O(N__15515),
            .I(N__15507));
    CascadeMux I__2809 (
            .O(N__15514),
            .I(N__15501));
    CascadeMux I__2808 (
            .O(N__15513),
            .I(N__15498));
    InMux I__2807 (
            .O(N__15510),
            .I(N__15495));
    InMux I__2806 (
            .O(N__15507),
            .I(N__15482));
    InMux I__2805 (
            .O(N__15506),
            .I(N__15482));
    InMux I__2804 (
            .O(N__15505),
            .I(N__15482));
    InMux I__2803 (
            .O(N__15504),
            .I(N__15482));
    InMux I__2802 (
            .O(N__15501),
            .I(N__15482));
    InMux I__2801 (
            .O(N__15498),
            .I(N__15482));
    LocalMux I__2800 (
            .O(N__15495),
            .I(N__15477));
    LocalMux I__2799 (
            .O(N__15482),
            .I(N__15477));
    Span4Mux_s2_v I__2798 (
            .O(N__15477),
            .I(N__15474));
    Odrv4 I__2797 (
            .O(N__15474),
            .I(\Lab_UT.min2_3 ));
    InMux I__2796 (
            .O(N__15471),
            .I(N__15468));
    LocalMux I__2795 (
            .O(N__15468),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__2794 (
            .O(N__15465),
            .I(N__15462));
    LocalMux I__2793 (
            .O(N__15462),
            .I(N__15459));
    Odrv4 I__2792 (
            .O(N__15459),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__2791 (
            .O(N__15456),
            .I(N__15453));
    LocalMux I__2790 (
            .O(N__15453),
            .I(N__15449));
    InMux I__2789 (
            .O(N__15452),
            .I(N__15446));
    Odrv4 I__2788 (
            .O(N__15449),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    LocalMux I__2787 (
            .O(N__15446),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    InMux I__2786 (
            .O(N__15441),
            .I(N__15438));
    LocalMux I__2785 (
            .O(N__15438),
            .I(\Lab_UT.dictrl.N_8 ));
    CascadeMux I__2784 (
            .O(N__15435),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_ ));
    InMux I__2783 (
            .O(N__15432),
            .I(N__15429));
    LocalMux I__2782 (
            .O(N__15429),
            .I(\Lab_UT.dictrl.N_20_0 ));
    CascadeMux I__2781 (
            .O(N__15426),
            .I(\Lab_UT.dictrl.N_18_0_cascade_ ));
    CascadeMux I__2780 (
            .O(N__15423),
            .I(N__15418));
    CascadeMux I__2779 (
            .O(N__15422),
            .I(N__15415));
    InMux I__2778 (
            .O(N__15421),
            .I(N__15401));
    InMux I__2777 (
            .O(N__15418),
            .I(N__15401));
    InMux I__2776 (
            .O(N__15415),
            .I(N__15401));
    InMux I__2775 (
            .O(N__15414),
            .I(N__15401));
    InMux I__2774 (
            .O(N__15413),
            .I(N__15390));
    InMux I__2773 (
            .O(N__15412),
            .I(N__15390));
    InMux I__2772 (
            .O(N__15411),
            .I(N__15390));
    InMux I__2771 (
            .O(N__15410),
            .I(N__15390));
    LocalMux I__2770 (
            .O(N__15401),
            .I(N__15387));
    InMux I__2769 (
            .O(N__15400),
            .I(N__15382));
    InMux I__2768 (
            .O(N__15399),
            .I(N__15382));
    LocalMux I__2767 (
            .O(N__15390),
            .I(N__15377));
    Span4Mux_s2_v I__2766 (
            .O(N__15387),
            .I(N__15377));
    LocalMux I__2765 (
            .O(N__15382),
            .I(N__15374));
    Span4Mux_v I__2764 (
            .O(N__15377),
            .I(N__15371));
    Odrv12 I__2763 (
            .O(N__15374),
            .I(\Lab_UT.dictrl.state_fast_3 ));
    Odrv4 I__2762 (
            .O(N__15371),
            .I(\Lab_UT.dictrl.state_fast_3 ));
    InMux I__2761 (
            .O(N__15366),
            .I(N__15361));
    InMux I__2760 (
            .O(N__15365),
            .I(N__15356));
    InMux I__2759 (
            .O(N__15364),
            .I(N__15356));
    LocalMux I__2758 (
            .O(N__15361),
            .I(N__15353));
    LocalMux I__2757 (
            .O(N__15356),
            .I(N__15348));
    Span4Mux_h I__2756 (
            .O(N__15353),
            .I(N__15348));
    Span4Mux_v I__2755 (
            .O(N__15348),
            .I(N__15345));
    Odrv4 I__2754 (
            .O(N__15345),
            .I(\Lab_UT.dictrl.state_fast_2 ));
    CascadeMux I__2753 (
            .O(N__15342),
            .I(N__15337));
    CascadeMux I__2752 (
            .O(N__15341),
            .I(N__15333));
    CascadeMux I__2751 (
            .O(N__15340),
            .I(N__15330));
    InMux I__2750 (
            .O(N__15337),
            .I(N__15325));
    InMux I__2749 (
            .O(N__15336),
            .I(N__15325));
    InMux I__2748 (
            .O(N__15333),
            .I(N__15320));
    InMux I__2747 (
            .O(N__15330),
            .I(N__15320));
    LocalMux I__2746 (
            .O(N__15325),
            .I(N__15317));
    LocalMux I__2745 (
            .O(N__15320),
            .I(N__15314));
    Odrv4 I__2744 (
            .O(N__15317),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    Odrv4 I__2743 (
            .O(N__15314),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    InMux I__2742 (
            .O(N__15309),
            .I(N__15306));
    LocalMux I__2741 (
            .O(N__15306),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_3_2 ));
    CascadeMux I__2740 (
            .O(N__15303),
            .I(N__15300));
    InMux I__2739 (
            .O(N__15300),
            .I(N__15297));
    LocalMux I__2738 (
            .O(N__15297),
            .I(\Lab_UT.dictrl.N_11_1 ));
    InMux I__2737 (
            .O(N__15294),
            .I(N__15291));
    LocalMux I__2736 (
            .O(N__15291),
            .I(N__15288));
    Span4Mux_v I__2735 (
            .O(N__15288),
            .I(N__15285));
    Odrv4 I__2734 (
            .O(N__15285),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_4_6 ));
    CascadeMux I__2733 (
            .O(N__15282),
            .I(\Lab_UT.dictrl.N_22_0_cascade_ ));
    InMux I__2732 (
            .O(N__15279),
            .I(N__15276));
    LocalMux I__2731 (
            .O(N__15276),
            .I(N__15273));
    Span4Mux_v I__2730 (
            .O(N__15273),
            .I(N__15270));
    Odrv4 I__2729 (
            .O(N__15270),
            .I(\Lab_UT.dictrl.g0_i_m2_0_a7_4_7 ));
    InMux I__2728 (
            .O(N__15267),
            .I(N__15264));
    LocalMux I__2727 (
            .O(N__15264),
            .I(N__15261));
    Odrv4 I__2726 (
            .O(N__15261),
            .I(\Lab_UT.dictrl.N_1110_1 ));
    CascadeMux I__2725 (
            .O(N__15258),
            .I(N__15254));
    CascadeMux I__2724 (
            .O(N__15257),
            .I(N__15250));
    InMux I__2723 (
            .O(N__15254),
            .I(N__15237));
    InMux I__2722 (
            .O(N__15253),
            .I(N__15237));
    InMux I__2721 (
            .O(N__15250),
            .I(N__15237));
    InMux I__2720 (
            .O(N__15249),
            .I(N__15237));
    InMux I__2719 (
            .O(N__15248),
            .I(N__15237));
    LocalMux I__2718 (
            .O(N__15237),
            .I(N__15234));
    Odrv4 I__2717 (
            .O(N__15234),
            .I(\Lab_UT.dictrl.N_1459_1 ));
    InMux I__2716 (
            .O(N__15231),
            .I(N__15228));
    LocalMux I__2715 (
            .O(N__15228),
            .I(\Lab_UT.dictrl.N_40_8 ));
    CascadeMux I__2714 (
            .O(N__15225),
            .I(\Lab_UT.dictrl.N_40_3_cascade_ ));
    InMux I__2713 (
            .O(N__15222),
            .I(N__15219));
    LocalMux I__2712 (
            .O(N__15219),
            .I(\Lab_UT.dictrl.N_1102_2 ));
    InMux I__2711 (
            .O(N__15216),
            .I(N__15213));
    LocalMux I__2710 (
            .O(N__15213),
            .I(N__15210));
    Odrv12 I__2709 (
            .O(N__15210),
            .I(\Lab_UT.dictrl.g2_1_2 ));
    CascadeMux I__2708 (
            .O(N__15207),
            .I(\Lab_UT.dictrl.N_1462_2_cascade_ ));
    InMux I__2707 (
            .O(N__15204),
            .I(N__15201));
    LocalMux I__2706 (
            .O(N__15201),
            .I(N__15197));
    InMux I__2705 (
            .O(N__15200),
            .I(N__15194));
    Span4Mux_v I__2704 (
            .O(N__15197),
            .I(N__15189));
    LocalMux I__2703 (
            .O(N__15194),
            .I(N__15189));
    Odrv4 I__2702 (
            .O(N__15189),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4 ));
    CascadeMux I__2701 (
            .O(N__15186),
            .I(\Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_ ));
    InMux I__2700 (
            .O(N__15183),
            .I(N__15177));
    InMux I__2699 (
            .O(N__15182),
            .I(N__15177));
    LocalMux I__2698 (
            .O(N__15177),
            .I(N__15174));
    Odrv4 I__2697 (
            .O(N__15174),
            .I(\Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3 ));
    CascadeMux I__2696 (
            .O(N__15171),
            .I(\Lab_UT.dictrl.N_11_0_cascade_ ));
    CascadeMux I__2695 (
            .O(N__15168),
            .I(N__15165));
    InMux I__2694 (
            .O(N__15165),
            .I(N__15162));
    LocalMux I__2693 (
            .O(N__15162),
            .I(N__15159));
    Odrv12 I__2692 (
            .O(N__15159),
            .I(\Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1 ));
    InMux I__2691 (
            .O(N__15156),
            .I(N__15138));
    InMux I__2690 (
            .O(N__15155),
            .I(N__15138));
    InMux I__2689 (
            .O(N__15154),
            .I(N__15138));
    InMux I__2688 (
            .O(N__15153),
            .I(N__15138));
    InMux I__2687 (
            .O(N__15152),
            .I(N__15138));
    InMux I__2686 (
            .O(N__15151),
            .I(N__15138));
    LocalMux I__2685 (
            .O(N__15138),
            .I(\Lab_UT.dictrl.m27_1 ));
    InMux I__2684 (
            .O(N__15135),
            .I(N__15125));
    InMux I__2683 (
            .O(N__15134),
            .I(N__15125));
    InMux I__2682 (
            .O(N__15133),
            .I(N__15116));
    InMux I__2681 (
            .O(N__15132),
            .I(N__15116));
    InMux I__2680 (
            .O(N__15131),
            .I(N__15116));
    InMux I__2679 (
            .O(N__15130),
            .I(N__15116));
    LocalMux I__2678 (
            .O(N__15125),
            .I(N__15111));
    LocalMux I__2677 (
            .O(N__15116),
            .I(N__15111));
    Odrv4 I__2676 (
            .O(N__15111),
            .I(\Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83 ));
    InMux I__2675 (
            .O(N__15108),
            .I(N__15105));
    LocalMux I__2674 (
            .O(N__15105),
            .I(N__15102));
    Odrv4 I__2673 (
            .O(N__15102),
            .I(\Lab_UT.dictrl.N_61 ));
    CascadeMux I__2672 (
            .O(N__15099),
            .I(\Lab_UT.dictrl.N_62_cascade_ ));
    CascadeMux I__2671 (
            .O(N__15096),
            .I(N__15093));
    InMux I__2670 (
            .O(N__15093),
            .I(N__15090));
    LocalMux I__2669 (
            .O(N__15090),
            .I(N__15087));
    Span4Mux_h I__2668 (
            .O(N__15087),
            .I(N__15083));
    InMux I__2667 (
            .O(N__15086),
            .I(N__15080));
    Span4Mux_v I__2666 (
            .O(N__15083),
            .I(N__15077));
    LocalMux I__2665 (
            .O(N__15080),
            .I(N__15074));
    Odrv4 I__2664 (
            .O(N__15077),
            .I(\Lab_UT.dictrl.N_9_0 ));
    Odrv4 I__2663 (
            .O(N__15074),
            .I(\Lab_UT.dictrl.N_9_0 ));
    InMux I__2662 (
            .O(N__15069),
            .I(N__15063));
    InMux I__2661 (
            .O(N__15068),
            .I(N__15063));
    LocalMux I__2660 (
            .O(N__15063),
            .I(\Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1 ));
    InMux I__2659 (
            .O(N__15060),
            .I(N__15057));
    LocalMux I__2658 (
            .O(N__15057),
            .I(N__15054));
    Span4Mux_s2_v I__2657 (
            .O(N__15054),
            .I(N__15051));
    Odrv4 I__2656 (
            .O(N__15051),
            .I(\Lab_UT.dictrl.state_fast_1 ));
    InMux I__2655 (
            .O(N__15048),
            .I(N__15033));
    InMux I__2654 (
            .O(N__15047),
            .I(N__15033));
    InMux I__2653 (
            .O(N__15046),
            .I(N__15033));
    InMux I__2652 (
            .O(N__15045),
            .I(N__15033));
    InMux I__2651 (
            .O(N__15044),
            .I(N__15033));
    LocalMux I__2650 (
            .O(N__15033),
            .I(N__15030));
    Span4Mux_h I__2649 (
            .O(N__15030),
            .I(N__15027));
    Span4Mux_h I__2648 (
            .O(N__15027),
            .I(N__15024));
    Odrv4 I__2647 (
            .O(N__15024),
            .I(\Lab_UT.dictrl.N_62_1 ));
    CascadeMux I__2646 (
            .O(N__15021),
            .I(N__15018));
    InMux I__2645 (
            .O(N__15018),
            .I(N__15015));
    LocalMux I__2644 (
            .O(N__15015),
            .I(N__15012));
    Span12Mux_v I__2643 (
            .O(N__15012),
            .I(N__15009));
    Odrv12 I__2642 (
            .O(N__15009),
            .I(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ));
    InMux I__2641 (
            .O(N__15006),
            .I(N__15003));
    LocalMux I__2640 (
            .O(N__15003),
            .I(N__14999));
    InMux I__2639 (
            .O(N__15002),
            .I(N__14996));
    Span4Mux_v I__2638 (
            .O(N__14999),
            .I(N__14993));
    LocalMux I__2637 (
            .O(N__14996),
            .I(N__14990));
    Odrv4 I__2636 (
            .O(N__14993),
            .I(\Lab_UT.dictrl.N_79 ));
    Odrv12 I__2635 (
            .O(N__14990),
            .I(\Lab_UT.dictrl.N_79 ));
    CascadeMux I__2634 (
            .O(N__14985),
            .I(N__14982));
    InMux I__2633 (
            .O(N__14982),
            .I(N__14979));
    LocalMux I__2632 (
            .O(N__14979),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    InMux I__2631 (
            .O(N__14976),
            .I(N__14973));
    LocalMux I__2630 (
            .O(N__14973),
            .I(N__14970));
    Span12Mux_s11_v I__2629 (
            .O(N__14970),
            .I(N__14967));
    Odrv12 I__2628 (
            .O(N__14967),
            .I(\Lab_UT.dictrl.N_99 ));
    InMux I__2627 (
            .O(N__14964),
            .I(N__14961));
    LocalMux I__2626 (
            .O(N__14961),
            .I(N__14954));
    InMux I__2625 (
            .O(N__14960),
            .I(N__14947));
    InMux I__2624 (
            .O(N__14959),
            .I(N__14944));
    InMux I__2623 (
            .O(N__14958),
            .I(N__14941));
    InMux I__2622 (
            .O(N__14957),
            .I(N__14938));
    Span4Mux_v I__2621 (
            .O(N__14954),
            .I(N__14935));
    InMux I__2620 (
            .O(N__14953),
            .I(N__14932));
    InMux I__2619 (
            .O(N__14952),
            .I(N__14929));
    InMux I__2618 (
            .O(N__14951),
            .I(N__14926));
    InMux I__2617 (
            .O(N__14950),
            .I(N__14923));
    LocalMux I__2616 (
            .O(N__14947),
            .I(N__14914));
    LocalMux I__2615 (
            .O(N__14944),
            .I(N__14914));
    LocalMux I__2614 (
            .O(N__14941),
            .I(N__14914));
    LocalMux I__2613 (
            .O(N__14938),
            .I(N__14914));
    Sp12to4 I__2612 (
            .O(N__14935),
            .I(N__14907));
    LocalMux I__2611 (
            .O(N__14932),
            .I(N__14907));
    LocalMux I__2610 (
            .O(N__14929),
            .I(N__14907));
    LocalMux I__2609 (
            .O(N__14926),
            .I(buart__rx_bitcount_3));
    LocalMux I__2608 (
            .O(N__14923),
            .I(buart__rx_bitcount_3));
    Odrv4 I__2607 (
            .O(N__14914),
            .I(buart__rx_bitcount_3));
    Odrv12 I__2606 (
            .O(N__14907),
            .I(buart__rx_bitcount_3));
    InMux I__2605 (
            .O(N__14898),
            .I(N__14895));
    LocalMux I__2604 (
            .O(N__14895),
            .I(N__14890));
    InMux I__2603 (
            .O(N__14894),
            .I(N__14887));
    InMux I__2602 (
            .O(N__14893),
            .I(N__14884));
    Span4Mux_v I__2601 (
            .O(N__14890),
            .I(N__14879));
    LocalMux I__2600 (
            .O(N__14887),
            .I(N__14874));
    LocalMux I__2599 (
            .O(N__14884),
            .I(N__14874));
    InMux I__2598 (
            .O(N__14883),
            .I(N__14869));
    InMux I__2597 (
            .O(N__14882),
            .I(N__14869));
    Span4Mux_h I__2596 (
            .O(N__14879),
            .I(N__14866));
    Span4Mux_h I__2595 (
            .O(N__14874),
            .I(N__14863));
    LocalMux I__2594 (
            .O(N__14869),
            .I(buart__rx_valid_3));
    Odrv4 I__2593 (
            .O(N__14866),
            .I(buart__rx_valid_3));
    Odrv4 I__2592 (
            .O(N__14863),
            .I(buart__rx_valid_3));
    CascadeMux I__2591 (
            .O(N__14856),
            .I(\Lab_UT.dictrl.g0_0_2_1_cascade_ ));
    InMux I__2590 (
            .O(N__14853),
            .I(N__14850));
    LocalMux I__2589 (
            .O(N__14850),
            .I(\Lab_UT.dictrl.g2_1_0 ));
    CascadeMux I__2588 (
            .O(N__14847),
            .I(\Lab_UT.dictrl.g0_0_2_cascade_ ));
    CascadeMux I__2587 (
            .O(N__14844),
            .I(N__14841));
    InMux I__2586 (
            .O(N__14841),
            .I(N__14838));
    LocalMux I__2585 (
            .O(N__14838),
            .I(\Lab_UT.dictrl.g0_12_a6_0_1 ));
    InMux I__2584 (
            .O(N__14835),
            .I(N__14829));
    CascadeMux I__2583 (
            .O(N__14834),
            .I(N__14821));
    InMux I__2582 (
            .O(N__14833),
            .I(N__14818));
    InMux I__2581 (
            .O(N__14832),
            .I(N__14815));
    LocalMux I__2580 (
            .O(N__14829),
            .I(N__14812));
    InMux I__2579 (
            .O(N__14828),
            .I(N__14803));
    InMux I__2578 (
            .O(N__14827),
            .I(N__14803));
    InMux I__2577 (
            .O(N__14826),
            .I(N__14803));
    InMux I__2576 (
            .O(N__14825),
            .I(N__14803));
    InMux I__2575 (
            .O(N__14824),
            .I(N__14798));
    InMux I__2574 (
            .O(N__14821),
            .I(N__14798));
    LocalMux I__2573 (
            .O(N__14818),
            .I(N__14793));
    LocalMux I__2572 (
            .O(N__14815),
            .I(N__14793));
    Span4Mux_s3_v I__2571 (
            .O(N__14812),
            .I(N__14786));
    LocalMux I__2570 (
            .O(N__14803),
            .I(N__14786));
    LocalMux I__2569 (
            .O(N__14798),
            .I(N__14786));
    Span4Mux_h I__2568 (
            .O(N__14793),
            .I(N__14783));
    Span4Mux_v I__2567 (
            .O(N__14786),
            .I(N__14780));
    Odrv4 I__2566 (
            .O(N__14783),
            .I(\Lab_UT.dictrl.state_2_rep1 ));
    Odrv4 I__2565 (
            .O(N__14780),
            .I(\Lab_UT.dictrl.state_2_rep1 ));
    CEMux I__2564 (
            .O(N__14775),
            .I(N__14772));
    LocalMux I__2563 (
            .O(N__14772),
            .I(N__14769));
    Span4Mux_h I__2562 (
            .O(N__14769),
            .I(N__14766));
    Span4Mux_h I__2561 (
            .O(N__14766),
            .I(N__14763));
    Odrv4 I__2560 (
            .O(N__14763),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    CascadeMux I__2559 (
            .O(N__14760),
            .I(\Lab_UT.didp.countrce4.q_5_3_cascade_ ));
    InMux I__2558 (
            .O(N__14757),
            .I(N__14752));
    InMux I__2557 (
            .O(N__14756),
            .I(N__14747));
    InMux I__2556 (
            .O(N__14755),
            .I(N__14747));
    LocalMux I__2555 (
            .O(N__14752),
            .I(\Lab_UT.di_AMtens_3 ));
    LocalMux I__2554 (
            .O(N__14747),
            .I(\Lab_UT.di_AMtens_3 ));
    CascadeMux I__2553 (
            .O(N__14742),
            .I(N__14739));
    InMux I__2552 (
            .O(N__14739),
            .I(N__14736));
    LocalMux I__2551 (
            .O(N__14736),
            .I(\Lab_UT.didp.countrce4.un20_qPone ));
    InMux I__2550 (
            .O(N__14733),
            .I(N__14730));
    LocalMux I__2549 (
            .O(N__14730),
            .I(\uu2.bitmap_pmux_15_ns_1 ));
    InMux I__2548 (
            .O(N__14727),
            .I(N__14723));
    InMux I__2547 (
            .O(N__14726),
            .I(N__14719));
    LocalMux I__2546 (
            .O(N__14723),
            .I(N__14715));
    InMux I__2545 (
            .O(N__14722),
            .I(N__14712));
    LocalMux I__2544 (
            .O(N__14719),
            .I(N__14709));
    InMux I__2543 (
            .O(N__14718),
            .I(N__14706));
    Odrv4 I__2542 (
            .O(N__14715),
            .I(o_One_Sec_Pulse));
    LocalMux I__2541 (
            .O(N__14712),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2540 (
            .O(N__14709),
            .I(o_One_Sec_Pulse));
    LocalMux I__2539 (
            .O(N__14706),
            .I(o_One_Sec_Pulse));
    InMux I__2538 (
            .O(N__14697),
            .I(N__14691));
    InMux I__2537 (
            .O(N__14696),
            .I(N__14691));
    LocalMux I__2536 (
            .O(N__14691),
            .I(N__14688));
    Odrv4 I__2535 (
            .O(N__14688),
            .I(\uu2.bitmapZ0Z_111 ));
    InMux I__2534 (
            .O(N__14685),
            .I(N__14680));
    InMux I__2533 (
            .O(N__14684),
            .I(N__14677));
    InMux I__2532 (
            .O(N__14683),
            .I(N__14674));
    LocalMux I__2531 (
            .O(N__14680),
            .I(N__14671));
    LocalMux I__2530 (
            .O(N__14677),
            .I(N__14668));
    LocalMux I__2529 (
            .O(N__14674),
            .I(N__14662));
    Span4Mux_h I__2528 (
            .O(N__14671),
            .I(N__14662));
    Span4Mux_v I__2527 (
            .O(N__14668),
            .I(N__14659));
    InMux I__2526 (
            .O(N__14667),
            .I(N__14656));
    Span4Mux_v I__2525 (
            .O(N__14662),
            .I(N__14653));
    Odrv4 I__2524 (
            .O(N__14659),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__2523 (
            .O(N__14656),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__2522 (
            .O(N__14653),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__2521 (
            .O(N__14646),
            .I(N__14643));
    LocalMux I__2520 (
            .O(N__14643),
            .I(\uu2.bitmapZ0Z_194 ));
    CascadeMux I__2519 (
            .O(N__14640),
            .I(N__14637));
    InMux I__2518 (
            .O(N__14637),
            .I(N__14634));
    LocalMux I__2517 (
            .O(N__14634),
            .I(N__14631));
    Odrv4 I__2516 (
            .O(N__14631),
            .I(\uu2.bitmapZ0Z_34 ));
    InMux I__2515 (
            .O(N__14628),
            .I(N__14625));
    LocalMux I__2514 (
            .O(N__14625),
            .I(\uu2.bitmapZ0Z_290 ));
    InMux I__2513 (
            .O(N__14622),
            .I(N__14619));
    LocalMux I__2512 (
            .O(N__14619),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__2511 (
            .O(N__14616),
            .I(N__14613));
    InMux I__2510 (
            .O(N__14613),
            .I(N__14610));
    LocalMux I__2509 (
            .O(N__14610),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__2508 (
            .O(N__14607),
            .I(N__14604));
    LocalMux I__2507 (
            .O(N__14604),
            .I(\uu2.N_207 ));
    InMux I__2506 (
            .O(N__14601),
            .I(N__14598));
    LocalMux I__2505 (
            .O(N__14598),
            .I(\uu2.bitmapZ0Z_168 ));
    CascadeMux I__2504 (
            .O(N__14595),
            .I(N__14592));
    InMux I__2503 (
            .O(N__14592),
            .I(N__14589));
    LocalMux I__2502 (
            .O(N__14589),
            .I(N__14586));
    Odrv4 I__2501 (
            .O(N__14586),
            .I(\uu2.N_195 ));
    InMux I__2500 (
            .O(N__14583),
            .I(N__14580));
    LocalMux I__2499 (
            .O(N__14580),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__2498 (
            .O(N__14577),
            .I(N__14574));
    LocalMux I__2497 (
            .O(N__14574),
            .I(N__14571));
    Odrv4 I__2496 (
            .O(N__14571),
            .I(\uu2.bitmapZ0Z_162 ));
    CascadeMux I__2495 (
            .O(N__14568),
            .I(N__14564));
    InMux I__2494 (
            .O(N__14567),
            .I(N__14556));
    InMux I__2493 (
            .O(N__14564),
            .I(N__14556));
    InMux I__2492 (
            .O(N__14563),
            .I(N__14556));
    LocalMux I__2491 (
            .O(N__14556),
            .I(\uu2.N_91 ));
    CascadeMux I__2490 (
            .O(N__14553),
            .I(\uu2.N_28_cascade_ ));
    CascadeMux I__2489 (
            .O(N__14550),
            .I(\uu2.bitmap_pmux_26_i_m2_1_cascade_ ));
    InMux I__2488 (
            .O(N__14547),
            .I(N__14544));
    LocalMux I__2487 (
            .O(N__14544),
            .I(N__14541));
    Odrv4 I__2486 (
            .O(N__14541),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    CascadeMux I__2485 (
            .O(N__14538),
            .I(\uu2.N_55_cascade_ ));
    InMux I__2484 (
            .O(N__14535),
            .I(N__14532));
    LocalMux I__2483 (
            .O(N__14532),
            .I(\uu2.bitmap_pmux_sn_i7_mux_0 ));
    CascadeMux I__2482 (
            .O(N__14529),
            .I(\uu2.N_406_cascade_ ));
    CascadeMux I__2481 (
            .O(N__14526),
            .I(N__14523));
    InMux I__2480 (
            .O(N__14523),
            .I(N__14517));
    InMux I__2479 (
            .O(N__14522),
            .I(N__14517));
    LocalMux I__2478 (
            .O(N__14517),
            .I(\uu2.bitmap_pmux ));
    InMux I__2477 (
            .O(N__14514),
            .I(N__14511));
    LocalMux I__2476 (
            .O(N__14511),
            .I(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ));
    InMux I__2475 (
            .O(N__14508),
            .I(N__14505));
    LocalMux I__2474 (
            .O(N__14505),
            .I(N__14502));
    Odrv4 I__2473 (
            .O(N__14502),
            .I(\Lab_UT.dictrl.next_state_RNO_3Z0Z_0 ));
    CascadeMux I__2472 (
            .O(N__14499),
            .I(\Lab_UT.dictrl.m67_am_1_0_cascade_ ));
    CascadeMux I__2471 (
            .O(N__14496),
            .I(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ));
    InMux I__2470 (
            .O(N__14493),
            .I(N__14490));
    LocalMux I__2469 (
            .O(N__14490),
            .I(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ));
    InMux I__2468 (
            .O(N__14487),
            .I(N__14484));
    LocalMux I__2467 (
            .O(N__14484),
            .I(\Lab_UT.dictrl.G_17_i_a5_0 ));
    InMux I__2466 (
            .O(N__14481),
            .I(N__14477));
    CascadeMux I__2465 (
            .O(N__14480),
            .I(N__14474));
    LocalMux I__2464 (
            .O(N__14477),
            .I(N__14471));
    InMux I__2463 (
            .O(N__14474),
            .I(N__14468));
    Span4Mux_h I__2462 (
            .O(N__14471),
            .I(N__14465));
    LocalMux I__2461 (
            .O(N__14468),
            .I(\Lab_UT.dictrl.N_65 ));
    Odrv4 I__2460 (
            .O(N__14465),
            .I(\Lab_UT.dictrl.N_65 ));
    CascadeMux I__2459 (
            .O(N__14460),
            .I(\Lab_UT.dictrl.N_65_cascade_ ));
    InMux I__2458 (
            .O(N__14457),
            .I(N__14454));
    LocalMux I__2457 (
            .O(N__14454),
            .I(\Lab_UT.dictrl.N_101 ));
    CascadeMux I__2456 (
            .O(N__14451),
            .I(N__14448));
    InMux I__2455 (
            .O(N__14448),
            .I(N__14445));
    LocalMux I__2454 (
            .O(N__14445),
            .I(N__14442));
    Odrv12 I__2453 (
            .O(N__14442),
            .I(\uu2.mem0.w_addr_5 ));
    CascadeMux I__2452 (
            .O(N__14439),
            .I(N__14436));
    InMux I__2451 (
            .O(N__14436),
            .I(N__14433));
    LocalMux I__2450 (
            .O(N__14433),
            .I(N__14430));
    Span4Mux_h I__2449 (
            .O(N__14430),
            .I(N__14427));
    Odrv4 I__2448 (
            .O(N__14427),
            .I(\uu2.mem0.w_addr_6 ));
    InMux I__2447 (
            .O(N__14424),
            .I(N__14421));
    LocalMux I__2446 (
            .O(N__14421),
            .I(N__14417));
    CascadeMux I__2445 (
            .O(N__14420),
            .I(N__14412));
    Span4Mux_s1_v I__2444 (
            .O(N__14417),
            .I(N__14409));
    InMux I__2443 (
            .O(N__14416),
            .I(N__14402));
    InMux I__2442 (
            .O(N__14415),
            .I(N__14402));
    InMux I__2441 (
            .O(N__14412),
            .I(N__14402));
    Odrv4 I__2440 (
            .O(N__14409),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__2439 (
            .O(N__14402),
            .I(\uu2.w_addr_userZ0Z_7 ));
    CascadeMux I__2438 (
            .O(N__14397),
            .I(N__14394));
    InMux I__2437 (
            .O(N__14394),
            .I(N__14391));
    LocalMux I__2436 (
            .O(N__14391),
            .I(N__14388));
    Span4Mux_h I__2435 (
            .O(N__14388),
            .I(N__14385));
    Odrv4 I__2434 (
            .O(N__14385),
            .I(\uu2.mem0.w_addr_7 ));
    InMux I__2433 (
            .O(N__14382),
            .I(N__14379));
    LocalMux I__2432 (
            .O(N__14379),
            .I(\Lab_UT.dictrl.g2_0_3_3 ));
    CascadeMux I__2431 (
            .O(N__14376),
            .I(\Lab_UT.dictrl.g2_0_4_3_cascade_ ));
    InMux I__2430 (
            .O(N__14373),
            .I(N__14363));
    InMux I__2429 (
            .O(N__14372),
            .I(N__14363));
    InMux I__2428 (
            .O(N__14371),
            .I(N__14360));
    InMux I__2427 (
            .O(N__14370),
            .I(N__14357));
    InMux I__2426 (
            .O(N__14369),
            .I(N__14352));
    InMux I__2425 (
            .O(N__14368),
            .I(N__14352));
    LocalMux I__2424 (
            .O(N__14363),
            .I(N__14347));
    LocalMux I__2423 (
            .O(N__14360),
            .I(N__14342));
    LocalMux I__2422 (
            .O(N__14357),
            .I(N__14342));
    LocalMux I__2421 (
            .O(N__14352),
            .I(N__14339));
    InMux I__2420 (
            .O(N__14351),
            .I(N__14334));
    InMux I__2419 (
            .O(N__14350),
            .I(N__14334));
    Span4Mux_v I__2418 (
            .O(N__14347),
            .I(N__14326));
    Span4Mux_h I__2417 (
            .O(N__14342),
            .I(N__14323));
    Span4Mux_v I__2416 (
            .O(N__14339),
            .I(N__14318));
    LocalMux I__2415 (
            .O(N__14334),
            .I(N__14318));
    InMux I__2414 (
            .O(N__14333),
            .I(N__14315));
    InMux I__2413 (
            .O(N__14332),
            .I(N__14306));
    InMux I__2412 (
            .O(N__14331),
            .I(N__14306));
    InMux I__2411 (
            .O(N__14330),
            .I(N__14306));
    InMux I__2410 (
            .O(N__14329),
            .I(N__14306));
    Odrv4 I__2409 (
            .O(N__14326),
            .I(\Lab_UT.dictrl.m12Z0Z_1 ));
    Odrv4 I__2408 (
            .O(N__14323),
            .I(\Lab_UT.dictrl.m12Z0Z_1 ));
    Odrv4 I__2407 (
            .O(N__14318),
            .I(\Lab_UT.dictrl.m12Z0Z_1 ));
    LocalMux I__2406 (
            .O(N__14315),
            .I(\Lab_UT.dictrl.m12Z0Z_1 ));
    LocalMux I__2405 (
            .O(N__14306),
            .I(\Lab_UT.dictrl.m12Z0Z_1 ));
    CascadeMux I__2404 (
            .O(N__14295),
            .I(\Lab_UT.dictrl.N_11_1_cascade_ ));
    InMux I__2403 (
            .O(N__14292),
            .I(N__14289));
    LocalMux I__2402 (
            .O(N__14289),
            .I(\Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0 ));
    CascadeMux I__2401 (
            .O(N__14286),
            .I(\Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_ ));
    InMux I__2400 (
            .O(N__14283),
            .I(N__14273));
    InMux I__2399 (
            .O(N__14282),
            .I(N__14270));
    InMux I__2398 (
            .O(N__14281),
            .I(N__14261));
    InMux I__2397 (
            .O(N__14280),
            .I(N__14261));
    InMux I__2396 (
            .O(N__14279),
            .I(N__14261));
    InMux I__2395 (
            .O(N__14278),
            .I(N__14261));
    InMux I__2394 (
            .O(N__14277),
            .I(N__14258));
    InMux I__2393 (
            .O(N__14276),
            .I(N__14255));
    LocalMux I__2392 (
            .O(N__14273),
            .I(bu_rx_data_fast_6));
    LocalMux I__2391 (
            .O(N__14270),
            .I(bu_rx_data_fast_6));
    LocalMux I__2390 (
            .O(N__14261),
            .I(bu_rx_data_fast_6));
    LocalMux I__2389 (
            .O(N__14258),
            .I(bu_rx_data_fast_6));
    LocalMux I__2388 (
            .O(N__14255),
            .I(bu_rx_data_fast_6));
    CEMux I__2387 (
            .O(N__14244),
            .I(N__14220));
    CEMux I__2386 (
            .O(N__14243),
            .I(N__14220));
    CEMux I__2385 (
            .O(N__14242),
            .I(N__14220));
    CEMux I__2384 (
            .O(N__14241),
            .I(N__14220));
    CEMux I__2383 (
            .O(N__14240),
            .I(N__14220));
    CEMux I__2382 (
            .O(N__14239),
            .I(N__14220));
    CEMux I__2381 (
            .O(N__14238),
            .I(N__14220));
    CEMux I__2380 (
            .O(N__14237),
            .I(N__14220));
    GlobalMux I__2379 (
            .O(N__14220),
            .I(N__14217));
    gio2CtrlBuf I__2378 (
            .O(N__14217),
            .I(\buart.Z_rx.sample_g ));
    InMux I__2377 (
            .O(N__14214),
            .I(N__14211));
    LocalMux I__2376 (
            .O(N__14211),
            .I(N__14208));
    Odrv12 I__2375 (
            .O(N__14208),
            .I(\Lab_UT.dictrl.N_100 ));
    CascadeMux I__2374 (
            .O(N__14205),
            .I(N__14202));
    InMux I__2373 (
            .O(N__14202),
            .I(N__14199));
    LocalMux I__2372 (
            .O(N__14199),
            .I(N__14196));
    Odrv12 I__2371 (
            .O(N__14196),
            .I(\Lab_UT.dictrl.next_state_RNO_8Z0Z_0 ));
    InMux I__2370 (
            .O(N__14193),
            .I(N__14190));
    LocalMux I__2369 (
            .O(N__14190),
            .I(N__14187));
    Odrv4 I__2368 (
            .O(N__14187),
            .I(\Lab_UT.dictrl.m63_d_0_ns_1 ));
    CascadeMux I__2367 (
            .O(N__14184),
            .I(\Lab_UT.dictrl.m59_3_cascade_ ));
    InMux I__2366 (
            .O(N__14181),
            .I(N__14178));
    LocalMux I__2365 (
            .O(N__14178),
            .I(\Lab_UT.dictrl.g2_0_3_4 ));
    CascadeMux I__2364 (
            .O(N__14175),
            .I(\Lab_UT.dictrl.g2_0_4_4_cascade_ ));
    InMux I__2363 (
            .O(N__14172),
            .I(N__14169));
    LocalMux I__2362 (
            .O(N__14169),
            .I(\Lab_UT.dictrl.g2_0_3_2 ));
    CascadeMux I__2361 (
            .O(N__14166),
            .I(\Lab_UT.dictrl.g2_0_4_2_cascade_ ));
    InMux I__2360 (
            .O(N__14163),
            .I(N__14160));
    LocalMux I__2359 (
            .O(N__14160),
            .I(\Lab_UT.dictrl.g2_0_3 ));
    CascadeMux I__2358 (
            .O(N__14157),
            .I(\Lab_UT.dictrl.g2_0_4_cascade_ ));
    InMux I__2357 (
            .O(N__14154),
            .I(N__14140));
    InMux I__2356 (
            .O(N__14153),
            .I(N__14140));
    InMux I__2355 (
            .O(N__14152),
            .I(N__14140));
    InMux I__2354 (
            .O(N__14151),
            .I(N__14140));
    InMux I__2353 (
            .O(N__14150),
            .I(N__14137));
    InMux I__2352 (
            .O(N__14149),
            .I(N__14134));
    LocalMux I__2351 (
            .O(N__14140),
            .I(N__14129));
    LocalMux I__2350 (
            .O(N__14137),
            .I(N__14129));
    LocalMux I__2349 (
            .O(N__14134),
            .I(bu_rx_data_fast_0));
    Odrv4 I__2348 (
            .O(N__14129),
            .I(bu_rx_data_fast_0));
    CascadeMux I__2347 (
            .O(N__14124),
            .I(N__14118));
    CascadeMux I__2346 (
            .O(N__14123),
            .I(N__14115));
    CascadeMux I__2345 (
            .O(N__14122),
            .I(N__14112));
    CascadeMux I__2344 (
            .O(N__14121),
            .I(N__14109));
    InMux I__2343 (
            .O(N__14118),
            .I(N__14098));
    InMux I__2342 (
            .O(N__14115),
            .I(N__14098));
    InMux I__2341 (
            .O(N__14112),
            .I(N__14098));
    InMux I__2340 (
            .O(N__14109),
            .I(N__14098));
    CascadeMux I__2339 (
            .O(N__14108),
            .I(N__14095));
    CascadeMux I__2338 (
            .O(N__14107),
            .I(N__14091));
    LocalMux I__2337 (
            .O(N__14098),
            .I(N__14088));
    InMux I__2336 (
            .O(N__14095),
            .I(N__14085));
    InMux I__2335 (
            .O(N__14094),
            .I(N__14082));
    InMux I__2334 (
            .O(N__14091),
            .I(N__14079));
    Span4Mux_v I__2333 (
            .O(N__14088),
            .I(N__14076));
    LocalMux I__2332 (
            .O(N__14085),
            .I(N__14073));
    LocalMux I__2331 (
            .O(N__14082),
            .I(N__14070));
    LocalMux I__2330 (
            .O(N__14079),
            .I(bu_rx_data_fast_4));
    Odrv4 I__2329 (
            .O(N__14076),
            .I(bu_rx_data_fast_4));
    Odrv4 I__2328 (
            .O(N__14073),
            .I(bu_rx_data_fast_4));
    Odrv4 I__2327 (
            .O(N__14070),
            .I(bu_rx_data_fast_4));
    InMux I__2326 (
            .O(N__14061),
            .I(N__14047));
    InMux I__2325 (
            .O(N__14060),
            .I(N__14047));
    InMux I__2324 (
            .O(N__14059),
            .I(N__14047));
    InMux I__2323 (
            .O(N__14058),
            .I(N__14047));
    InMux I__2322 (
            .O(N__14057),
            .I(N__14042));
    InMux I__2321 (
            .O(N__14056),
            .I(N__14039));
    LocalMux I__2320 (
            .O(N__14047),
            .I(N__14036));
    InMux I__2319 (
            .O(N__14046),
            .I(N__14031));
    InMux I__2318 (
            .O(N__14045),
            .I(N__14031));
    LocalMux I__2317 (
            .O(N__14042),
            .I(N__14026));
    LocalMux I__2316 (
            .O(N__14039),
            .I(N__14026));
    Span4Mux_v I__2315 (
            .O(N__14036),
            .I(N__14023));
    LocalMux I__2314 (
            .O(N__14031),
            .I(N__14018));
    Span4Mux_v I__2313 (
            .O(N__14026),
            .I(N__14018));
    Odrv4 I__2312 (
            .O(N__14023),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__2311 (
            .O(N__14018),
            .I(bu_rx_data_3_rep1));
    CascadeMux I__2310 (
            .O(N__14013),
            .I(N__14010));
    InMux I__2309 (
            .O(N__14010),
            .I(N__14007));
    LocalMux I__2308 (
            .O(N__14007),
            .I(N__14003));
    InMux I__2307 (
            .O(N__14006),
            .I(N__14000));
    Odrv4 I__2306 (
            .O(N__14003),
            .I(\Lab_UT.dictrl.m15Z0Z_1 ));
    LocalMux I__2305 (
            .O(N__14000),
            .I(\Lab_UT.dictrl.m15Z0Z_1 ));
    InMux I__2304 (
            .O(N__13995),
            .I(N__13992));
    LocalMux I__2303 (
            .O(N__13992),
            .I(N__13987));
    InMux I__2302 (
            .O(N__13991),
            .I(N__13984));
    InMux I__2301 (
            .O(N__13990),
            .I(N__13981));
    Odrv4 I__2300 (
            .O(N__13987),
            .I(\Lab_UT.dictrl.N_88_mux ));
    LocalMux I__2299 (
            .O(N__13984),
            .I(\Lab_UT.dictrl.N_88_mux ));
    LocalMux I__2298 (
            .O(N__13981),
            .I(\Lab_UT.dictrl.N_88_mux ));
    CascadeMux I__2297 (
            .O(N__13974),
            .I(\Lab_UT.dictrl.g2_0_4_1_cascade_ ));
    CascadeMux I__2296 (
            .O(N__13971),
            .I(\Lab_UT.dictrl.m53_d_1_2_cascade_ ));
    CascadeMux I__2295 (
            .O(N__13968),
            .I(\Lab_UT.dictrl.N_45_cascade_ ));
    InMux I__2294 (
            .O(N__13965),
            .I(N__13960));
    InMux I__2293 (
            .O(N__13964),
            .I(N__13951));
    InMux I__2292 (
            .O(N__13963),
            .I(N__13948));
    LocalMux I__2291 (
            .O(N__13960),
            .I(N__13945));
    InMux I__2290 (
            .O(N__13959),
            .I(N__13936));
    InMux I__2289 (
            .O(N__13958),
            .I(N__13936));
    InMux I__2288 (
            .O(N__13957),
            .I(N__13936));
    InMux I__2287 (
            .O(N__13956),
            .I(N__13936));
    InMux I__2286 (
            .O(N__13955),
            .I(N__13931));
    InMux I__2285 (
            .O(N__13954),
            .I(N__13931));
    LocalMux I__2284 (
            .O(N__13951),
            .I(N__13928));
    LocalMux I__2283 (
            .O(N__13948),
            .I(N__13919));
    Span4Mux_v I__2282 (
            .O(N__13945),
            .I(N__13919));
    LocalMux I__2281 (
            .O(N__13936),
            .I(N__13919));
    LocalMux I__2280 (
            .O(N__13931),
            .I(N__13916));
    Span4Mux_h I__2279 (
            .O(N__13928),
            .I(N__13913));
    InMux I__2278 (
            .O(N__13927),
            .I(N__13908));
    InMux I__2277 (
            .O(N__13926),
            .I(N__13908));
    Span4Mux_h I__2276 (
            .O(N__13919),
            .I(N__13905));
    Span4Mux_h I__2275 (
            .O(N__13916),
            .I(N__13902));
    Odrv4 I__2274 (
            .O(N__13913),
            .I(bu_rx_data_1_rep2));
    LocalMux I__2273 (
            .O(N__13908),
            .I(bu_rx_data_1_rep2));
    Odrv4 I__2272 (
            .O(N__13905),
            .I(bu_rx_data_1_rep2));
    Odrv4 I__2271 (
            .O(N__13902),
            .I(bu_rx_data_1_rep2));
    InMux I__2270 (
            .O(N__13893),
            .I(N__13890));
    LocalMux I__2269 (
            .O(N__13890),
            .I(\Lab_UT.dictrl.g2_0_3_1 ));
    CascadeMux I__2268 (
            .O(N__13887),
            .I(N__13878));
    CascadeMux I__2267 (
            .O(N__13886),
            .I(N__13872));
    CascadeMux I__2266 (
            .O(N__13885),
            .I(N__13869));
    CascadeMux I__2265 (
            .O(N__13884),
            .I(N__13866));
    InMux I__2264 (
            .O(N__13883),
            .I(N__13863));
    InMux I__2263 (
            .O(N__13882),
            .I(N__13860));
    InMux I__2262 (
            .O(N__13881),
            .I(N__13853));
    InMux I__2261 (
            .O(N__13878),
            .I(N__13853));
    InMux I__2260 (
            .O(N__13877),
            .I(N__13853));
    InMux I__2259 (
            .O(N__13876),
            .I(N__13850));
    InMux I__2258 (
            .O(N__13875),
            .I(N__13847));
    InMux I__2257 (
            .O(N__13872),
            .I(N__13840));
    InMux I__2256 (
            .O(N__13869),
            .I(N__13840));
    InMux I__2255 (
            .O(N__13866),
            .I(N__13840));
    LocalMux I__2254 (
            .O(N__13863),
            .I(N__13835));
    LocalMux I__2253 (
            .O(N__13860),
            .I(N__13830));
    LocalMux I__2252 (
            .O(N__13853),
            .I(N__13830));
    LocalMux I__2251 (
            .O(N__13850),
            .I(N__13827));
    LocalMux I__2250 (
            .O(N__13847),
            .I(N__13824));
    LocalMux I__2249 (
            .O(N__13840),
            .I(N__13821));
    InMux I__2248 (
            .O(N__13839),
            .I(N__13816));
    InMux I__2247 (
            .O(N__13838),
            .I(N__13816));
    Span4Mux_h I__2246 (
            .O(N__13835),
            .I(N__13811));
    Span4Mux_h I__2245 (
            .O(N__13830),
            .I(N__13811));
    Span4Mux_v I__2244 (
            .O(N__13827),
            .I(N__13804));
    Span4Mux_v I__2243 (
            .O(N__13824),
            .I(N__13804));
    Span4Mux_v I__2242 (
            .O(N__13821),
            .I(N__13804));
    LocalMux I__2241 (
            .O(N__13816),
            .I(bu_rx_data_2_rep2));
    Odrv4 I__2240 (
            .O(N__13811),
            .I(bu_rx_data_2_rep2));
    Odrv4 I__2239 (
            .O(N__13804),
            .I(bu_rx_data_2_rep2));
    CascadeMux I__2238 (
            .O(N__13797),
            .I(N__13794));
    InMux I__2237 (
            .O(N__13794),
            .I(N__13791));
    LocalMux I__2236 (
            .O(N__13791),
            .I(N__13787));
    CascadeMux I__2235 (
            .O(N__13790),
            .I(N__13784));
    Span4Mux_v I__2234 (
            .O(N__13787),
            .I(N__13781));
    InMux I__2233 (
            .O(N__13784),
            .I(N__13778));
    Odrv4 I__2232 (
            .O(N__13781),
            .I(Lab_UT_dictrl_m59_1));
    LocalMux I__2231 (
            .O(N__13778),
            .I(Lab_UT_dictrl_m59_1));
    InMux I__2230 (
            .O(N__13773),
            .I(N__13770));
    LocalMux I__2229 (
            .O(N__13770),
            .I(N__13767));
    Odrv4 I__2228 (
            .O(N__13767),
            .I(\Lab_UT.dictrl.g0_12_a6_3_6 ));
    InMux I__2227 (
            .O(N__13764),
            .I(N__13761));
    LocalMux I__2226 (
            .O(N__13761),
            .I(N__13758));
    Odrv4 I__2225 (
            .O(N__13758),
            .I(\Lab_UT.dictrl.N_10 ));
    InMux I__2224 (
            .O(N__13755),
            .I(N__13752));
    LocalMux I__2223 (
            .O(N__13752),
            .I(\Lab_UT.dictrl.g0_12_1 ));
    CascadeMux I__2222 (
            .O(N__13749),
            .I(\Lab_UT.dictrl.m15Z0Z_1_cascade_ ));
    InMux I__2221 (
            .O(N__13746),
            .I(N__13743));
    LocalMux I__2220 (
            .O(N__13743),
            .I(N__13740));
    Odrv4 I__2219 (
            .O(N__13740),
            .I(\Lab_UT.dictrl.N_8_0 ));
    CascadeMux I__2218 (
            .O(N__13737),
            .I(\Lab_UT.dictrl.N_93_cascade_ ));
    CascadeMux I__2217 (
            .O(N__13734),
            .I(N__13731));
    InMux I__2216 (
            .O(N__13731),
            .I(N__13728));
    LocalMux I__2215 (
            .O(N__13728),
            .I(\Lab_UT.dictrl.N_10_0 ));
    CascadeMux I__2214 (
            .O(N__13725),
            .I(N__13722));
    InMux I__2213 (
            .O(N__13722),
            .I(N__13719));
    LocalMux I__2212 (
            .O(N__13719),
            .I(N__13716));
    Span4Mux_h I__2211 (
            .O(N__13716),
            .I(N__13713));
    Odrv4 I__2210 (
            .O(N__13713),
            .I(\Lab_UT.dictrl.g0_i_a4_0_1 ));
    InMux I__2209 (
            .O(N__13710),
            .I(N__13707));
    LocalMux I__2208 (
            .O(N__13707),
            .I(\Lab_UT.dictrl.g0_i_a4_0_3 ));
    InMux I__2207 (
            .O(N__13704),
            .I(N__13692));
    InMux I__2206 (
            .O(N__13703),
            .I(N__13692));
    InMux I__2205 (
            .O(N__13702),
            .I(N__13692));
    InMux I__2204 (
            .O(N__13701),
            .I(N__13689));
    CascadeMux I__2203 (
            .O(N__13700),
            .I(N__13684));
    CascadeMux I__2202 (
            .O(N__13699),
            .I(N__13681));
    LocalMux I__2201 (
            .O(N__13692),
            .I(N__13673));
    LocalMux I__2200 (
            .O(N__13689),
            .I(N__13673));
    CascadeMux I__2199 (
            .O(N__13688),
            .I(N__13668));
    InMux I__2198 (
            .O(N__13687),
            .I(N__13663));
    InMux I__2197 (
            .O(N__13684),
            .I(N__13663));
    InMux I__2196 (
            .O(N__13681),
            .I(N__13658));
    InMux I__2195 (
            .O(N__13680),
            .I(N__13658));
    InMux I__2194 (
            .O(N__13679),
            .I(N__13653));
    InMux I__2193 (
            .O(N__13678),
            .I(N__13653));
    Span4Mux_h I__2192 (
            .O(N__13673),
            .I(N__13650));
    InMux I__2191 (
            .O(N__13672),
            .I(N__13647));
    InMux I__2190 (
            .O(N__13671),
            .I(N__13642));
    InMux I__2189 (
            .O(N__13668),
            .I(N__13642));
    LocalMux I__2188 (
            .O(N__13663),
            .I(N__13639));
    LocalMux I__2187 (
            .O(N__13658),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    LocalMux I__2186 (
            .O(N__13653),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2185 (
            .O(N__13650),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    LocalMux I__2184 (
            .O(N__13647),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    LocalMux I__2183 (
            .O(N__13642),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2182 (
            .O(N__13639),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    InMux I__2181 (
            .O(N__13626),
            .I(N__13623));
    LocalMux I__2180 (
            .O(N__13623),
            .I(\Lab_UT.dispString.b1_m_1 ));
    CascadeMux I__2179 (
            .O(N__13620),
            .I(\Lab_UT.dispString.m67_ns_1_cascade_ ));
    InMux I__2178 (
            .O(N__13617),
            .I(N__13614));
    LocalMux I__2177 (
            .O(N__13614),
            .I(N__13611));
    Odrv4 I__2176 (
            .O(N__13611),
            .I(\Lab_UT.dispString.N_143 ));
    InMux I__2175 (
            .O(N__13608),
            .I(N__13605));
    LocalMux I__2174 (
            .O(N__13605),
            .I(N__13601));
    InMux I__2173 (
            .O(N__13604),
            .I(N__13598));
    Odrv4 I__2172 (
            .O(N__13601),
            .I(\Lab_UT.dispString.N_23_0 ));
    LocalMux I__2171 (
            .O(N__13598),
            .I(\Lab_UT.dispString.N_23_0 ));
    InMux I__2170 (
            .O(N__13593),
            .I(N__13590));
    LocalMux I__2169 (
            .O(N__13590),
            .I(\Lab_UT.dispString.N_158 ));
    CascadeMux I__2168 (
            .O(N__13587),
            .I(\Lab_UT.dispString.m90_ns_1_cascade_ ));
    InMux I__2167 (
            .O(N__13584),
            .I(N__13581));
    LocalMux I__2166 (
            .O(N__13581),
            .I(N__13578));
    Odrv4 I__2165 (
            .O(N__13578),
            .I(\Lab_UT.dispString.N_164 ));
    InMux I__2164 (
            .O(N__13575),
            .I(N__13563));
    InMux I__2163 (
            .O(N__13574),
            .I(N__13563));
    InMux I__2162 (
            .O(N__13573),
            .I(N__13556));
    InMux I__2161 (
            .O(N__13572),
            .I(N__13556));
    InMux I__2160 (
            .O(N__13571),
            .I(N__13556));
    InMux I__2159 (
            .O(N__13570),
            .I(N__13550));
    InMux I__2158 (
            .O(N__13569),
            .I(N__13550));
    InMux I__2157 (
            .O(N__13568),
            .I(N__13547));
    LocalMux I__2156 (
            .O(N__13563),
            .I(N__13530));
    LocalMux I__2155 (
            .O(N__13556),
            .I(N__13530));
    InMux I__2154 (
            .O(N__13555),
            .I(N__13527));
    LocalMux I__2153 (
            .O(N__13550),
            .I(N__13524));
    LocalMux I__2152 (
            .O(N__13547),
            .I(N__13521));
    InMux I__2151 (
            .O(N__13546),
            .I(N__13514));
    InMux I__2150 (
            .O(N__13545),
            .I(N__13514));
    InMux I__2149 (
            .O(N__13544),
            .I(N__13514));
    InMux I__2148 (
            .O(N__13543),
            .I(N__13511));
    InMux I__2147 (
            .O(N__13542),
            .I(N__13508));
    InMux I__2146 (
            .O(N__13541),
            .I(N__13505));
    InMux I__2145 (
            .O(N__13540),
            .I(N__13502));
    InMux I__2144 (
            .O(N__13539),
            .I(N__13493));
    InMux I__2143 (
            .O(N__13538),
            .I(N__13493));
    InMux I__2142 (
            .O(N__13537),
            .I(N__13493));
    InMux I__2141 (
            .O(N__13536),
            .I(N__13493));
    InMux I__2140 (
            .O(N__13535),
            .I(N__13490));
    Span4Mux_h I__2139 (
            .O(N__13530),
            .I(N__13487));
    LocalMux I__2138 (
            .O(N__13527),
            .I(N__13484));
    Span4Mux_v I__2137 (
            .O(N__13524),
            .I(N__13477));
    Span4Mux_v I__2136 (
            .O(N__13521),
            .I(N__13477));
    LocalMux I__2135 (
            .O(N__13514),
            .I(N__13477));
    LocalMux I__2134 (
            .O(N__13511),
            .I(N__13474));
    LocalMux I__2133 (
            .O(N__13508),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2132 (
            .O(N__13505),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2131 (
            .O(N__13502),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2130 (
            .O(N__13493),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2129 (
            .O(N__13490),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2128 (
            .O(N__13487),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2127 (
            .O(N__13484),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2126 (
            .O(N__13477),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2125 (
            .O(N__13474),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    CascadeMux I__2124 (
            .O(N__13455),
            .I(N__13448));
    CascadeMux I__2123 (
            .O(N__13454),
            .I(N__13444));
    CascadeMux I__2122 (
            .O(N__13453),
            .I(N__13441));
    CascadeMux I__2121 (
            .O(N__13452),
            .I(N__13438));
    CascadeMux I__2120 (
            .O(N__13451),
            .I(N__13435));
    InMux I__2119 (
            .O(N__13448),
            .I(N__13426));
    InMux I__2118 (
            .O(N__13447),
            .I(N__13426));
    InMux I__2117 (
            .O(N__13444),
            .I(N__13426));
    InMux I__2116 (
            .O(N__13441),
            .I(N__13423));
    InMux I__2115 (
            .O(N__13438),
            .I(N__13416));
    InMux I__2114 (
            .O(N__13435),
            .I(N__13416));
    InMux I__2113 (
            .O(N__13434),
            .I(N__13416));
    CascadeMux I__2112 (
            .O(N__13433),
            .I(N__13405));
    LocalMux I__2111 (
            .O(N__13426),
            .I(N__13400));
    LocalMux I__2110 (
            .O(N__13423),
            .I(N__13395));
    LocalMux I__2109 (
            .O(N__13416),
            .I(N__13395));
    InMux I__2108 (
            .O(N__13415),
            .I(N__13390));
    InMux I__2107 (
            .O(N__13414),
            .I(N__13390));
    InMux I__2106 (
            .O(N__13413),
            .I(N__13387));
    InMux I__2105 (
            .O(N__13412),
            .I(N__13382));
    InMux I__2104 (
            .O(N__13411),
            .I(N__13382));
    InMux I__2103 (
            .O(N__13410),
            .I(N__13375));
    InMux I__2102 (
            .O(N__13409),
            .I(N__13375));
    InMux I__2101 (
            .O(N__13408),
            .I(N__13375));
    InMux I__2100 (
            .O(N__13405),
            .I(N__13370));
    InMux I__2099 (
            .O(N__13404),
            .I(N__13370));
    InMux I__2098 (
            .O(N__13403),
            .I(N__13367));
    Span4Mux_v I__2097 (
            .O(N__13400),
            .I(N__13360));
    Span4Mux_v I__2096 (
            .O(N__13395),
            .I(N__13360));
    LocalMux I__2095 (
            .O(N__13390),
            .I(N__13360));
    LocalMux I__2094 (
            .O(N__13387),
            .I(N__13357));
    LocalMux I__2093 (
            .O(N__13382),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2092 (
            .O(N__13375),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2091 (
            .O(N__13370),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2090 (
            .O(N__13367),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__2089 (
            .O(N__13360),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__2088 (
            .O(N__13357),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    InMux I__2087 (
            .O(N__13344),
            .I(N__13341));
    LocalMux I__2086 (
            .O(N__13341),
            .I(\Lab_UT.dispString.N_166 ));
    InMux I__2085 (
            .O(N__13338),
            .I(N__13335));
    LocalMux I__2084 (
            .O(N__13335),
            .I(N__13332));
    Odrv4 I__2083 (
            .O(N__13332),
            .I(\Lab_UT.dispString.N_167 ));
    InMux I__2082 (
            .O(N__13329),
            .I(N__13326));
    LocalMux I__2081 (
            .O(N__13326),
            .I(N__13323));
    Odrv4 I__2080 (
            .O(N__13323),
            .I(Lab_UT_dictrl_g1_0_3));
    InMux I__2079 (
            .O(N__13320),
            .I(N__13317));
    LocalMux I__2078 (
            .O(N__13317),
            .I(N__13314));
    Span4Mux_s2_v I__2077 (
            .O(N__13314),
            .I(N__13311));
    Odrv4 I__2076 (
            .O(N__13311),
            .I(\uu2.mem0.w_data_2 ));
    InMux I__2075 (
            .O(N__13308),
            .I(N__13305));
    LocalMux I__2074 (
            .O(N__13305),
            .I(\Lab_UT.dispString.N_145 ));
    CascadeMux I__2073 (
            .O(N__13302),
            .I(\Lab_UT.dispString.N_146_cascade_ ));
    InMux I__2072 (
            .O(N__13299),
            .I(N__13290));
    InMux I__2071 (
            .O(N__13298),
            .I(N__13290));
    InMux I__2070 (
            .O(N__13297),
            .I(N__13290));
    LocalMux I__2069 (
            .O(N__13290),
            .I(L3_tx_data_2));
    InMux I__2068 (
            .O(N__13287),
            .I(N__13283));
    CascadeMux I__2067 (
            .O(N__13286),
            .I(N__13280));
    LocalMux I__2066 (
            .O(N__13283),
            .I(N__13276));
    InMux I__2065 (
            .O(N__13280),
            .I(N__13271));
    InMux I__2064 (
            .O(N__13279),
            .I(N__13271));
    Odrv4 I__2063 (
            .O(N__13276),
            .I(L3_tx_data_0));
    LocalMux I__2062 (
            .O(N__13271),
            .I(L3_tx_data_0));
    InMux I__2061 (
            .O(N__13266),
            .I(N__13262));
    CascadeMux I__2060 (
            .O(N__13265),
            .I(N__13258));
    LocalMux I__2059 (
            .O(N__13262),
            .I(N__13255));
    InMux I__2058 (
            .O(N__13261),
            .I(N__13250));
    InMux I__2057 (
            .O(N__13258),
            .I(N__13250));
    Odrv4 I__2056 (
            .O(N__13255),
            .I(L3_tx_data_6));
    LocalMux I__2055 (
            .O(N__13250),
            .I(L3_tx_data_6));
    CascadeMux I__2054 (
            .O(N__13245),
            .I(\Lab_UT.dispString.m82_ns_1_cascade_ ));
    CascadeMux I__2053 (
            .O(N__13242),
            .I(\Lab_UT.dispString.N_156_cascade_ ));
    CascadeMux I__2052 (
            .O(N__13239),
            .I(N__13235));
    InMux I__2051 (
            .O(N__13238),
            .I(N__13231));
    InMux I__2050 (
            .O(N__13235),
            .I(N__13226));
    InMux I__2049 (
            .O(N__13234),
            .I(N__13226));
    LocalMux I__2048 (
            .O(N__13231),
            .I(N__13223));
    LocalMux I__2047 (
            .O(N__13226),
            .I(N__13220));
    Odrv12 I__2046 (
            .O(N__13223),
            .I(L3_tx_data_3));
    Odrv4 I__2045 (
            .O(N__13220),
            .I(L3_tx_data_3));
    CascadeMux I__2044 (
            .O(N__13215),
            .I(\uu2.un1_w_user_lf_0_cascade_ ));
    InMux I__2043 (
            .O(N__13212),
            .I(N__13209));
    LocalMux I__2042 (
            .O(N__13209),
            .I(\uu2.un1_w_user_lfZ0Z_4 ));
    InMux I__2041 (
            .O(N__13206),
            .I(N__13203));
    LocalMux I__2040 (
            .O(N__13203),
            .I(\uu2.un1_w_user_lf_0 ));
    InMux I__2039 (
            .O(N__13200),
            .I(N__13197));
    LocalMux I__2038 (
            .O(N__13197),
            .I(N__13194));
    Span4Mux_s0_v I__2037 (
            .O(N__13194),
            .I(N__13189));
    InMux I__2036 (
            .O(N__13193),
            .I(N__13184));
    InMux I__2035 (
            .O(N__13192),
            .I(N__13184));
    Odrv4 I__2034 (
            .O(N__13189),
            .I(L3_tx_data_5));
    LocalMux I__2033 (
            .O(N__13184),
            .I(L3_tx_data_5));
    InMux I__2032 (
            .O(N__13179),
            .I(N__13176));
    LocalMux I__2031 (
            .O(N__13176),
            .I(N__13171));
    InMux I__2030 (
            .O(N__13175),
            .I(N__13166));
    InMux I__2029 (
            .O(N__13174),
            .I(N__13166));
    Odrv4 I__2028 (
            .O(N__13171),
            .I(L3_tx_data_1));
    LocalMux I__2027 (
            .O(N__13166),
            .I(L3_tx_data_1));
    InMux I__2026 (
            .O(N__13161),
            .I(N__13158));
    LocalMux I__2025 (
            .O(N__13158),
            .I(N__13153));
    InMux I__2024 (
            .O(N__13157),
            .I(N__13148));
    InMux I__2023 (
            .O(N__13156),
            .I(N__13148));
    Odrv4 I__2022 (
            .O(N__13153),
            .I(L3_tx_data_4));
    LocalMux I__2021 (
            .O(N__13148),
            .I(L3_tx_data_4));
    CascadeMux I__2020 (
            .O(N__13143),
            .I(\uu2.m35Z0Z_4_cascade_ ));
    CascadeMux I__2019 (
            .O(N__13140),
            .I(\uu2.un1_w_user_cr_0_cascade_ ));
    InMux I__2018 (
            .O(N__13137),
            .I(N__13134));
    LocalMux I__2017 (
            .O(N__13134),
            .I(N__13131));
    Odrv4 I__2016 (
            .O(N__13131),
            .I(\uu2.mem0.N_69_i ));
    InMux I__2015 (
            .O(N__13128),
            .I(N__13122));
    InMux I__2014 (
            .O(N__13127),
            .I(N__13122));
    LocalMux I__2013 (
            .O(N__13122),
            .I(\uu2.N_96_mux ));
    InMux I__2012 (
            .O(N__13119),
            .I(N__13116));
    LocalMux I__2011 (
            .O(N__13116),
            .I(N__13113));
    Odrv4 I__2010 (
            .O(N__13113),
            .I(\uu2.mem0.N_71_i ));
    InMux I__2009 (
            .O(N__13110),
            .I(N__13107));
    LocalMux I__2008 (
            .O(N__13107),
            .I(N__13104));
    Odrv4 I__2007 (
            .O(N__13104),
            .I(\uu2.mem0.N_91_mux ));
    InMux I__2006 (
            .O(N__13101),
            .I(N__13098));
    LocalMux I__2005 (
            .O(N__13098),
            .I(N__13095));
    Span4Mux_s3_h I__2004 (
            .O(N__13095),
            .I(N__13092));
    Odrv4 I__2003 (
            .O(N__13092),
            .I(\uu2.mem0.N_50_i ));
    InMux I__2002 (
            .O(N__13089),
            .I(N__13084));
    CascadeMux I__2001 (
            .O(N__13088),
            .I(N__13081));
    CascadeMux I__2000 (
            .O(N__13087),
            .I(N__13078));
    LocalMux I__1999 (
            .O(N__13084),
            .I(N__13074));
    InMux I__1998 (
            .O(N__13081),
            .I(N__13071));
    InMux I__1997 (
            .O(N__13078),
            .I(N__13066));
    InMux I__1996 (
            .O(N__13077),
            .I(N__13066));
    Odrv12 I__1995 (
            .O(N__13074),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1994 (
            .O(N__13071),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1993 (
            .O(N__13066),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__1992 (
            .O(N__13059),
            .I(N__13056));
    InMux I__1991 (
            .O(N__13056),
            .I(N__13053));
    LocalMux I__1990 (
            .O(N__13053),
            .I(N__13050));
    Span4Mux_s1_v I__1989 (
            .O(N__13050),
            .I(N__13047));
    Span4Mux_s3_h I__1988 (
            .O(N__13047),
            .I(N__13044));
    Odrv4 I__1987 (
            .O(N__13044),
            .I(\uu2.mem0.w_addr_3 ));
    CascadeMux I__1986 (
            .O(N__13041),
            .I(N__13038));
    InMux I__1985 (
            .O(N__13038),
            .I(N__13035));
    LocalMux I__1984 (
            .O(N__13035),
            .I(N__13032));
    Span4Mux_s1_v I__1983 (
            .O(N__13032),
            .I(N__13029));
    Odrv4 I__1982 (
            .O(N__13029),
            .I(\uu2.mem0.w_addr_4 ));
    CascadeMux I__1981 (
            .O(N__13026),
            .I(\uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_ ));
    InMux I__1980 (
            .O(N__13023),
            .I(N__13020));
    LocalMux I__1979 (
            .O(N__13020),
            .I(\Lab_UT.dictrl.N_10_1 ));
    CascadeMux I__1978 (
            .O(N__13017),
            .I(\Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_ ));
    InMux I__1977 (
            .O(N__13014),
            .I(N__13011));
    LocalMux I__1976 (
            .O(N__13011),
            .I(\Lab_UT.dictrl.g0_i_m2_1_1 ));
    InMux I__1975 (
            .O(N__13008),
            .I(N__13005));
    LocalMux I__1974 (
            .O(N__13005),
            .I(\Lab_UT.dictrl.g0_i_m2_1_a6_3_2 ));
    InMux I__1973 (
            .O(N__13002),
            .I(N__12997));
    InMux I__1972 (
            .O(N__13001),
            .I(N__12989));
    InMux I__1971 (
            .O(N__13000),
            .I(N__12989));
    LocalMux I__1970 (
            .O(N__12997),
            .I(N__12986));
    InMux I__1969 (
            .O(N__12996),
            .I(N__12979));
    InMux I__1968 (
            .O(N__12995),
            .I(N__12979));
    InMux I__1967 (
            .O(N__12994),
            .I(N__12979));
    LocalMux I__1966 (
            .O(N__12989),
            .I(N__12976));
    Odrv4 I__1965 (
            .O(N__12986),
            .I(bu_rx_data_fast_3));
    LocalMux I__1964 (
            .O(N__12979),
            .I(bu_rx_data_fast_3));
    Odrv4 I__1963 (
            .O(N__12976),
            .I(bu_rx_data_fast_3));
    InMux I__1962 (
            .O(N__12969),
            .I(N__12963));
    InMux I__1961 (
            .O(N__12968),
            .I(N__12963));
    LocalMux I__1960 (
            .O(N__12963),
            .I(\Lab_UT.dictrl.N_7_0 ));
    CascadeMux I__1959 (
            .O(N__12960),
            .I(\Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_ ));
    InMux I__1958 (
            .O(N__12957),
            .I(N__12954));
    LocalMux I__1957 (
            .O(N__12954),
            .I(\Lab_UT.dictrl.G_17_i_a5_1 ));
    InMux I__1956 (
            .O(N__12951),
            .I(N__12948));
    LocalMux I__1955 (
            .O(N__12948),
            .I(N__12945));
    Odrv12 I__1954 (
            .O(N__12945),
            .I(\uu2.mem0.N_66_i ));
    InMux I__1953 (
            .O(N__12942),
            .I(N__12939));
    LocalMux I__1952 (
            .O(N__12939),
            .I(N__12936));
    Span4Mux_h I__1951 (
            .O(N__12936),
            .I(N__12933));
    Odrv4 I__1950 (
            .O(N__12933),
            .I(\uu2.mem0.N_56_i ));
    CascadeMux I__1949 (
            .O(N__12930),
            .I(N__12926));
    InMux I__1948 (
            .O(N__12929),
            .I(N__12921));
    InMux I__1947 (
            .O(N__12926),
            .I(N__12921));
    LocalMux I__1946 (
            .O(N__12921),
            .I(\uu2.N_95_mux ));
    CascadeMux I__1945 (
            .O(N__12918),
            .I(\uu2.N_96_mux_cascade_ ));
    InMux I__1944 (
            .O(N__12915),
            .I(N__12912));
    LocalMux I__1943 (
            .O(N__12912),
            .I(N__12909));
    Span4Mux_v I__1942 (
            .O(N__12909),
            .I(N__12906));
    Odrv4 I__1941 (
            .O(N__12906),
            .I(\uu2.mem0.N_63_i ));
    CascadeMux I__1940 (
            .O(N__12903),
            .I(N__12900));
    InMux I__1939 (
            .O(N__12900),
            .I(N__12897));
    LocalMux I__1938 (
            .O(N__12897),
            .I(N__12894));
    Odrv12 I__1937 (
            .O(N__12894),
            .I(\Lab_UT.dispString.m107_eZ0Z_3 ));
    InMux I__1936 (
            .O(N__12891),
            .I(N__12881));
    InMux I__1935 (
            .O(N__12890),
            .I(N__12881));
    InMux I__1934 (
            .O(N__12889),
            .I(N__12881));
    CascadeMux I__1933 (
            .O(N__12888),
            .I(N__12878));
    LocalMux I__1932 (
            .O(N__12881),
            .I(N__12875));
    InMux I__1931 (
            .O(N__12878),
            .I(N__12872));
    Odrv4 I__1930 (
            .O(N__12875),
            .I(bu_rx_data_fast_5));
    LocalMux I__1929 (
            .O(N__12872),
            .I(bu_rx_data_fast_5));
    CascadeMux I__1928 (
            .O(N__12867),
            .I(\Lab_UT.dictrl.N_10_1_cascade_ ));
    InMux I__1927 (
            .O(N__12864),
            .I(N__12861));
    LocalMux I__1926 (
            .O(N__12861),
            .I(N__12858));
    Span4Mux_v I__1925 (
            .O(N__12858),
            .I(N__12855));
    Odrv4 I__1924 (
            .O(N__12855),
            .I(\Lab_UT.dictrl.N_17_0 ));
    CascadeMux I__1923 (
            .O(N__12852),
            .I(\Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_ ));
    InMux I__1922 (
            .O(N__12849),
            .I(N__12846));
    LocalMux I__1921 (
            .O(N__12846),
            .I(N__12843));
    Odrv4 I__1920 (
            .O(N__12843),
            .I(N_22));
    InMux I__1919 (
            .O(N__12840),
            .I(N__12837));
    LocalMux I__1918 (
            .O(N__12837),
            .I(\Lab_UT.dictrl.N_1105_0 ));
    InMux I__1917 (
            .O(N__12834),
            .I(N__12830));
    CascadeMux I__1916 (
            .O(N__12833),
            .I(N__12824));
    LocalMux I__1915 (
            .O(N__12830),
            .I(N__12821));
    InMux I__1914 (
            .O(N__12829),
            .I(N__12818));
    InMux I__1913 (
            .O(N__12828),
            .I(N__12811));
    InMux I__1912 (
            .O(N__12827),
            .I(N__12811));
    InMux I__1911 (
            .O(N__12824),
            .I(N__12811));
    Odrv4 I__1910 (
            .O(N__12821),
            .I(bu_rx_data_fast_7));
    LocalMux I__1909 (
            .O(N__12818),
            .I(bu_rx_data_fast_7));
    LocalMux I__1908 (
            .O(N__12811),
            .I(bu_rx_data_fast_7));
    InMux I__1907 (
            .O(N__12804),
            .I(N__12801));
    LocalMux I__1906 (
            .O(N__12801),
            .I(\buart.Z_rx.G_17_i_a5_2_5 ));
    InMux I__1905 (
            .O(N__12798),
            .I(N__12795));
    LocalMux I__1904 (
            .O(N__12795),
            .I(N__12792));
    Span4Mux_v I__1903 (
            .O(N__12792),
            .I(N__12789));
    Odrv4 I__1902 (
            .O(N__12789),
            .I(\buart.Z_rx.G_17_i_a5_2_4 ));
    CascadeMux I__1901 (
            .O(N__12786),
            .I(G_17_i_a5_2_6_cascade_));
    InMux I__1900 (
            .O(N__12783),
            .I(N__12770));
    InMux I__1899 (
            .O(N__12782),
            .I(N__12770));
    InMux I__1898 (
            .O(N__12781),
            .I(N__12770));
    InMux I__1897 (
            .O(N__12780),
            .I(N__12770));
    InMux I__1896 (
            .O(N__12779),
            .I(N__12767));
    LocalMux I__1895 (
            .O(N__12770),
            .I(bu_rx_data_fast_1));
    LocalMux I__1894 (
            .O(N__12767),
            .I(bu_rx_data_fast_1));
    CascadeMux I__1893 (
            .O(N__12762),
            .I(N__12758));
    CascadeMux I__1892 (
            .O(N__12761),
            .I(N__12755));
    InMux I__1891 (
            .O(N__12758),
            .I(N__12743));
    InMux I__1890 (
            .O(N__12755),
            .I(N__12743));
    InMux I__1889 (
            .O(N__12754),
            .I(N__12743));
    InMux I__1888 (
            .O(N__12753),
            .I(N__12743));
    InMux I__1887 (
            .O(N__12752),
            .I(N__12740));
    LocalMux I__1886 (
            .O(N__12743),
            .I(bu_rx_data_fast_2));
    LocalMux I__1885 (
            .O(N__12740),
            .I(bu_rx_data_fast_2));
    CascadeMux I__1884 (
            .O(N__12735),
            .I(\Lab_UT.dictrl.g2_0_3_0_cascade_ ));
    InMux I__1883 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__1882 (
            .O(N__12729),
            .I(\Lab_UT.dictrl.g2_0_4_0 ));
    CascadeMux I__1881 (
            .O(N__12726),
            .I(N__12722));
    InMux I__1880 (
            .O(N__12725),
            .I(N__12718));
    InMux I__1879 (
            .O(N__12722),
            .I(N__12713));
    InMux I__1878 (
            .O(N__12721),
            .I(N__12713));
    LocalMux I__1877 (
            .O(N__12718),
            .I(N__12705));
    LocalMux I__1876 (
            .O(N__12713),
            .I(N__12702));
    InMux I__1875 (
            .O(N__12712),
            .I(N__12691));
    InMux I__1874 (
            .O(N__12711),
            .I(N__12691));
    InMux I__1873 (
            .O(N__12710),
            .I(N__12691));
    InMux I__1872 (
            .O(N__12709),
            .I(N__12691));
    InMux I__1871 (
            .O(N__12708),
            .I(N__12691));
    Odrv4 I__1870 (
            .O(N__12705),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__1869 (
            .O(N__12702),
            .I(bu_rx_data_1_rep1));
    LocalMux I__1868 (
            .O(N__12691),
            .I(bu_rx_data_1_rep1));
    CascadeMux I__1867 (
            .O(N__12684),
            .I(N__12679));
    CascadeMux I__1866 (
            .O(N__12683),
            .I(N__12674));
    CascadeMux I__1865 (
            .O(N__12682),
            .I(N__12671));
    InMux I__1864 (
            .O(N__12679),
            .I(N__12661));
    InMux I__1863 (
            .O(N__12678),
            .I(N__12661));
    InMux I__1862 (
            .O(N__12677),
            .I(N__12661));
    InMux I__1861 (
            .O(N__12674),
            .I(N__12650));
    InMux I__1860 (
            .O(N__12671),
            .I(N__12650));
    InMux I__1859 (
            .O(N__12670),
            .I(N__12650));
    InMux I__1858 (
            .O(N__12669),
            .I(N__12650));
    InMux I__1857 (
            .O(N__12668),
            .I(N__12650));
    LocalMux I__1856 (
            .O(N__12661),
            .I(N__12647));
    LocalMux I__1855 (
            .O(N__12650),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__1854 (
            .O(N__12647),
            .I(bu_rx_data_2_rep1));
    InMux I__1853 (
            .O(N__12642),
            .I(N__12639));
    LocalMux I__1852 (
            .O(N__12639),
            .I(\Lab_UT.dictrl.m27_d_1 ));
    CascadeMux I__1851 (
            .O(N__12636),
            .I(\Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_ ));
    InMux I__1850 (
            .O(N__12633),
            .I(N__12630));
    LocalMux I__1849 (
            .O(N__12630),
            .I(N__12627));
    Odrv4 I__1848 (
            .O(N__12627),
            .I(\Lab_UT.dictrl.G_17_i_a5_0_0 ));
    CascadeMux I__1847 (
            .O(N__12624),
            .I(N__12621));
    InMux I__1846 (
            .O(N__12621),
            .I(N__12618));
    LocalMux I__1845 (
            .O(N__12618),
            .I(\Lab_UT.dictrl.m71Z0Z_0 ));
    InMux I__1844 (
            .O(N__12615),
            .I(N__12599));
    InMux I__1843 (
            .O(N__12614),
            .I(N__12599));
    InMux I__1842 (
            .O(N__12613),
            .I(N__12599));
    InMux I__1841 (
            .O(N__12612),
            .I(N__12599));
    InMux I__1840 (
            .O(N__12611),
            .I(N__12590));
    InMux I__1839 (
            .O(N__12610),
            .I(N__12590));
    InMux I__1838 (
            .O(N__12609),
            .I(N__12590));
    InMux I__1837 (
            .O(N__12608),
            .I(N__12590));
    LocalMux I__1836 (
            .O(N__12599),
            .I(N__12585));
    LocalMux I__1835 (
            .O(N__12590),
            .I(N__12585));
    Span4Mux_h I__1834 (
            .O(N__12585),
            .I(N__12582));
    Odrv4 I__1833 (
            .O(N__12582),
            .I(N_105_mux));
    InMux I__1832 (
            .O(N__12579),
            .I(N__12576));
    LocalMux I__1831 (
            .O(N__12576),
            .I(\Lab_UT.dispString.N_186 ));
    InMux I__1830 (
            .O(N__12573),
            .I(N__12570));
    LocalMux I__1829 (
            .O(N__12570),
            .I(\Lab_UT.dictrl.g0_12_a6_3Z0Z_7 ));
    CascadeMux I__1828 (
            .O(N__12567),
            .I(\Lab_UT.dictrl.g0_12_a6_3_8_cascade_ ));
    InMux I__1827 (
            .O(N__12564),
            .I(N__12561));
    LocalMux I__1826 (
            .O(N__12561),
            .I(\Lab_UT.dictrl.N_16 ));
    InMux I__1825 (
            .O(N__12558),
            .I(N__12555));
    LocalMux I__1824 (
            .O(N__12555),
            .I(N_10_2));
    InMux I__1823 (
            .O(N__12552),
            .I(N__12549));
    LocalMux I__1822 (
            .O(N__12549),
            .I(\Lab_UT.dictrl.N_97_mux_0_0_0 ));
    CascadeMux I__1821 (
            .O(N__12546),
            .I(\Lab_UT.dictrl.g0_10_1_cascade_ ));
    CascadeMux I__1820 (
            .O(N__12543),
            .I(N__12540));
    InMux I__1819 (
            .O(N__12540),
            .I(N__12537));
    LocalMux I__1818 (
            .O(N__12537),
            .I(N__12534));
    Span4Mux_v I__1817 (
            .O(N__12534),
            .I(N__12531));
    Odrv4 I__1816 (
            .O(N__12531),
            .I(\Lab_UT.dictrl.m63_d_0_ns_1_1 ));
    InMux I__1815 (
            .O(N__12528),
            .I(N__12524));
    InMux I__1814 (
            .O(N__12527),
            .I(N__12521));
    LocalMux I__1813 (
            .O(N__12524),
            .I(N__12518));
    LocalMux I__1812 (
            .O(N__12521),
            .I(N__12515));
    Odrv4 I__1811 (
            .O(N__12518),
            .I(\Lab_UT.dispString.N_112_mux ));
    Odrv4 I__1810 (
            .O(N__12515),
            .I(\Lab_UT.dispString.N_112_mux ));
    InMux I__1809 (
            .O(N__12510),
            .I(N__12507));
    LocalMux I__1808 (
            .O(N__12507),
            .I(\uu0.sec_clkDZ0 ));
    CascadeMux I__1807 (
            .O(N__12504),
            .I(\Lab_UT.alarmstate_1_0_i_1_cascade_ ));
    CascadeMux I__1806 (
            .O(N__12501),
            .I(G_215_cascade_));
    InMux I__1805 (
            .O(N__12498),
            .I(N__12495));
    LocalMux I__1804 (
            .O(N__12495),
            .I(G_214));
    InMux I__1803 (
            .O(N__12492),
            .I(N__12486));
    InMux I__1802 (
            .O(N__12491),
            .I(N__12486));
    LocalMux I__1801 (
            .O(N__12486),
            .I(G_216));
    CascadeMux I__1800 (
            .O(N__12483),
            .I(G_214_cascade_));
    InMux I__1799 (
            .O(N__12480),
            .I(N__12477));
    LocalMux I__1798 (
            .O(N__12477),
            .I(\Lab_UT.m57 ));
    CascadeMux I__1797 (
            .O(N__12474),
            .I(N__12470));
    CascadeMux I__1796 (
            .O(N__12473),
            .I(N__12464));
    InMux I__1795 (
            .O(N__12470),
            .I(N__12455));
    InMux I__1794 (
            .O(N__12469),
            .I(N__12455));
    InMux I__1793 (
            .O(N__12468),
            .I(N__12455));
    InMux I__1792 (
            .O(N__12467),
            .I(N__12455));
    InMux I__1791 (
            .O(N__12464),
            .I(N__12447));
    LocalMux I__1790 (
            .O(N__12455),
            .I(N__12444));
    InMux I__1789 (
            .O(N__12454),
            .I(N__12441));
    InMux I__1788 (
            .O(N__12453),
            .I(N__12432));
    InMux I__1787 (
            .O(N__12452),
            .I(N__12432));
    InMux I__1786 (
            .O(N__12451),
            .I(N__12432));
    InMux I__1785 (
            .O(N__12450),
            .I(N__12432));
    LocalMux I__1784 (
            .O(N__12447),
            .I(G_213));
    Odrv4 I__1783 (
            .O(N__12444),
            .I(G_213));
    LocalMux I__1782 (
            .O(N__12441),
            .I(G_213));
    LocalMux I__1781 (
            .O(N__12432),
            .I(G_213));
    InMux I__1780 (
            .O(N__12423),
            .I(N__12409));
    InMux I__1779 (
            .O(N__12422),
            .I(N__12409));
    InMux I__1778 (
            .O(N__12421),
            .I(N__12409));
    InMux I__1777 (
            .O(N__12420),
            .I(N__12409));
    CascadeMux I__1776 (
            .O(N__12419),
            .I(N__12403));
    InMux I__1775 (
            .O(N__12418),
            .I(N__12399));
    LocalMux I__1774 (
            .O(N__12409),
            .I(N__12396));
    InMux I__1773 (
            .O(N__12408),
            .I(N__12393));
    InMux I__1772 (
            .O(N__12407),
            .I(N__12384));
    InMux I__1771 (
            .O(N__12406),
            .I(N__12384));
    InMux I__1770 (
            .O(N__12403),
            .I(N__12384));
    InMux I__1769 (
            .O(N__12402),
            .I(N__12384));
    LocalMux I__1768 (
            .O(N__12399),
            .I(G_215));
    Odrv4 I__1767 (
            .O(N__12396),
            .I(G_215));
    LocalMux I__1766 (
            .O(N__12393),
            .I(G_215));
    LocalMux I__1765 (
            .O(N__12384),
            .I(G_215));
    CascadeMux I__1764 (
            .O(N__12375),
            .I(G_213_cascade_));
    InMux I__1763 (
            .O(N__12372),
            .I(N__12365));
    InMux I__1762 (
            .O(N__12371),
            .I(N__12365));
    InMux I__1761 (
            .O(N__12370),
            .I(N__12362));
    LocalMux I__1760 (
            .O(N__12365),
            .I(N__12359));
    LocalMux I__1759 (
            .O(N__12362),
            .I(\uu0.un88_ci_3 ));
    Odrv12 I__1758 (
            .O(N__12359),
            .I(\uu0.un88_ci_3 ));
    InMux I__1757 (
            .O(N__12354),
            .I(N__12351));
    LocalMux I__1756 (
            .O(N__12351),
            .I(N__12347));
    InMux I__1755 (
            .O(N__12350),
            .I(N__12342));
    Span4Mux_h I__1754 (
            .O(N__12347),
            .I(N__12339));
    InMux I__1753 (
            .O(N__12346),
            .I(N__12334));
    InMux I__1752 (
            .O(N__12345),
            .I(N__12334));
    LocalMux I__1751 (
            .O(N__12342),
            .I(N__12331));
    Odrv4 I__1750 (
            .O(N__12339),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__1749 (
            .O(N__12334),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1748 (
            .O(N__12331),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__1747 (
            .O(N__12324),
            .I(N__12321));
    LocalMux I__1746 (
            .O(N__12321),
            .I(N__12318));
    Odrv4 I__1745 (
            .O(N__12318),
            .I(\uu0.un99_ci_0 ));
    CascadeMux I__1744 (
            .O(N__12315),
            .I(N__12312));
    InMux I__1743 (
            .O(N__12312),
            .I(N__12309));
    LocalMux I__1742 (
            .O(N__12309),
            .I(\Lab_UT.dispString.dOutP_0_iv_2_tz_1 ));
    CascadeMux I__1741 (
            .O(N__12306),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_ ));
    InMux I__1740 (
            .O(N__12303),
            .I(N__12300));
    LocalMux I__1739 (
            .O(N__12300),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_1_1 ));
    CascadeMux I__1738 (
            .O(N__12297),
            .I(N__12294));
    InMux I__1737 (
            .O(N__12294),
            .I(N__12291));
    LocalMux I__1736 (
            .O(N__12291),
            .I(\Lab_UT.dispString.m74_ns_1 ));
    InMux I__1735 (
            .O(N__12288),
            .I(N__12285));
    LocalMux I__1734 (
            .O(N__12285),
            .I(\Lab_UT.dispString.m77_ns_1 ));
    InMux I__1733 (
            .O(N__12282),
            .I(N__12278));
    InMux I__1732 (
            .O(N__12281),
            .I(N__12275));
    LocalMux I__1731 (
            .O(N__12278),
            .I(N__12270));
    LocalMux I__1730 (
            .O(N__12275),
            .I(N__12270));
    Odrv4 I__1729 (
            .O(N__12270),
            .I(\Lab_UT.dispString.N_30_i ));
    InMux I__1728 (
            .O(N__12267),
            .I(N__12264));
    LocalMux I__1727 (
            .O(N__12264),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_1 ));
    InMux I__1726 (
            .O(N__12261),
            .I(N__12258));
    LocalMux I__1725 (
            .O(N__12258),
            .I(N__12254));
    InMux I__1724 (
            .O(N__12257),
            .I(N__12250));
    Span4Mux_h I__1723 (
            .O(N__12254),
            .I(N__12247));
    InMux I__1722 (
            .O(N__12253),
            .I(N__12244));
    LocalMux I__1721 (
            .O(N__12250),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv4 I__1720 (
            .O(N__12247),
            .I(\uu0.l_countZ0Z_5 ));
    LocalMux I__1719 (
            .O(N__12244),
            .I(\uu0.l_countZ0Z_5 ));
    InMux I__1718 (
            .O(N__12237),
            .I(N__12233));
    InMux I__1717 (
            .O(N__12236),
            .I(N__12230));
    LocalMux I__1716 (
            .O(N__12233),
            .I(N__12227));
    LocalMux I__1715 (
            .O(N__12230),
            .I(N__12222));
    Span4Mux_h I__1714 (
            .O(N__12227),
            .I(N__12219));
    InMux I__1713 (
            .O(N__12226),
            .I(N__12214));
    InMux I__1712 (
            .O(N__12225),
            .I(N__12214));
    Odrv12 I__1711 (
            .O(N__12222),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__1710 (
            .O(N__12219),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__1709 (
            .O(N__12214),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__1708 (
            .O(N__12207),
            .I(N__12201));
    InMux I__1707 (
            .O(N__12206),
            .I(N__12201));
    LocalMux I__1706 (
            .O(N__12201),
            .I(\uu2.un284_ci ));
    CascadeMux I__1705 (
            .O(N__12198),
            .I(N__12195));
    InMux I__1704 (
            .O(N__12195),
            .I(N__12186));
    InMux I__1703 (
            .O(N__12194),
            .I(N__12186));
    InMux I__1702 (
            .O(N__12193),
            .I(N__12179));
    InMux I__1701 (
            .O(N__12192),
            .I(N__12179));
    InMux I__1700 (
            .O(N__12191),
            .I(N__12179));
    LocalMux I__1699 (
            .O(N__12186),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1698 (
            .O(N__12179),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__1697 (
            .O(N__12174),
            .I(N__12162));
    InMux I__1696 (
            .O(N__12173),
            .I(N__12162));
    InMux I__1695 (
            .O(N__12172),
            .I(N__12162));
    InMux I__1694 (
            .O(N__12171),
            .I(N__12159));
    InMux I__1693 (
            .O(N__12170),
            .I(N__12154));
    InMux I__1692 (
            .O(N__12169),
            .I(N__12154));
    LocalMux I__1691 (
            .O(N__12162),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1690 (
            .O(N__12159),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1689 (
            .O(N__12154),
            .I(\uu2.l_countZ0Z_0 ));
    CEMux I__1688 (
            .O(N__12147),
            .I(N__12144));
    LocalMux I__1687 (
            .O(N__12144),
            .I(N__12141));
    Odrv4 I__1686 (
            .O(N__12141),
            .I(\uu2.un28_w_addr_user_i_0 ));
    InMux I__1685 (
            .O(N__12138),
            .I(N__12134));
    InMux I__1684 (
            .O(N__12137),
            .I(N__12131));
    LocalMux I__1683 (
            .O(N__12134),
            .I(\uu2.un1_l_count_1_0 ));
    LocalMux I__1682 (
            .O(N__12131),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1681 (
            .O(N__12126),
            .I(N__12099));
    InMux I__1680 (
            .O(N__12125),
            .I(N__12099));
    InMux I__1679 (
            .O(N__12124),
            .I(N__12099));
    InMux I__1678 (
            .O(N__12123),
            .I(N__12099));
    InMux I__1677 (
            .O(N__12122),
            .I(N__12099));
    InMux I__1676 (
            .O(N__12121),
            .I(N__12099));
    InMux I__1675 (
            .O(N__12120),
            .I(N__12099));
    CascadeMux I__1674 (
            .O(N__12119),
            .I(N__12095));
    InMux I__1673 (
            .O(N__12118),
            .I(N__12084));
    InMux I__1672 (
            .O(N__12117),
            .I(N__12084));
    InMux I__1671 (
            .O(N__12116),
            .I(N__12084));
    InMux I__1670 (
            .O(N__12115),
            .I(N__12084));
    CascadeMux I__1669 (
            .O(N__12114),
            .I(N__12081));
    LocalMux I__1668 (
            .O(N__12099),
            .I(N__12078));
    InMux I__1667 (
            .O(N__12098),
            .I(N__12069));
    InMux I__1666 (
            .O(N__12095),
            .I(N__12069));
    InMux I__1665 (
            .O(N__12094),
            .I(N__12069));
    InMux I__1664 (
            .O(N__12093),
            .I(N__12069));
    LocalMux I__1663 (
            .O(N__12084),
            .I(N__12066));
    InMux I__1662 (
            .O(N__12081),
            .I(N__12063));
    Span4Mux_h I__1661 (
            .O(N__12078),
            .I(N__12056));
    LocalMux I__1660 (
            .O(N__12069),
            .I(N__12056));
    Span4Mux_h I__1659 (
            .O(N__12066),
            .I(N__12056));
    LocalMux I__1658 (
            .O(N__12063),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1657 (
            .O(N__12056),
            .I(vbuf_tx_data_rdy));
    CascadeMux I__1656 (
            .O(N__12051),
            .I(\uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ));
    CascadeMux I__1655 (
            .O(N__12048),
            .I(N__12044));
    InMux I__1654 (
            .O(N__12047),
            .I(N__12028));
    InMux I__1653 (
            .O(N__12044),
            .I(N__12028));
    InMux I__1652 (
            .O(N__12043),
            .I(N__12028));
    InMux I__1651 (
            .O(N__12042),
            .I(N__12028));
    InMux I__1650 (
            .O(N__12041),
            .I(N__12028));
    InMux I__1649 (
            .O(N__12040),
            .I(N__12023));
    InMux I__1648 (
            .O(N__12039),
            .I(N__12023));
    LocalMux I__1647 (
            .O(N__12028),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1646 (
            .O(N__12023),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__1645 (
            .O(N__12018),
            .I(\uu2.un426_ci_3_cascade_ ));
    CascadeMux I__1644 (
            .O(N__12015),
            .I(N__12011));
    InMux I__1643 (
            .O(N__12014),
            .I(N__12008));
    InMux I__1642 (
            .O(N__12011),
            .I(N__12002));
    LocalMux I__1641 (
            .O(N__12008),
            .I(N__11999));
    InMux I__1640 (
            .O(N__12007),
            .I(N__11996));
    InMux I__1639 (
            .O(N__12006),
            .I(N__11991));
    InMux I__1638 (
            .O(N__12005),
            .I(N__11991));
    LocalMux I__1637 (
            .O(N__12002),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1636 (
            .O(N__11999),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1635 (
            .O(N__11996),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1634 (
            .O(N__11991),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__1633 (
            .O(N__11982),
            .I(N__11979));
    LocalMux I__1632 (
            .O(N__11979),
            .I(N__11973));
    InMux I__1631 (
            .O(N__11978),
            .I(N__11970));
    InMux I__1630 (
            .O(N__11977),
            .I(N__11965));
    InMux I__1629 (
            .O(N__11976),
            .I(N__11965));
    Odrv4 I__1628 (
            .O(N__11973),
            .I(\uu2.un404_ci_0 ));
    LocalMux I__1627 (
            .O(N__11970),
            .I(\uu2.un404_ci_0 ));
    LocalMux I__1626 (
            .O(N__11965),
            .I(\uu2.un404_ci_0 ));
    InMux I__1625 (
            .O(N__11958),
            .I(N__11951));
    InMux I__1624 (
            .O(N__11957),
            .I(N__11942));
    InMux I__1623 (
            .O(N__11956),
            .I(N__11942));
    InMux I__1622 (
            .O(N__11955),
            .I(N__11942));
    InMux I__1621 (
            .O(N__11954),
            .I(N__11942));
    LocalMux I__1620 (
            .O(N__11951),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__1619 (
            .O(N__11942),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__1618 (
            .O(N__11937),
            .I(N__11934));
    InMux I__1617 (
            .O(N__11934),
            .I(N__11931));
    LocalMux I__1616 (
            .O(N__11931),
            .I(N__11925));
    CascadeMux I__1615 (
            .O(N__11930),
            .I(N__11922));
    InMux I__1614 (
            .O(N__11929),
            .I(N__11917));
    InMux I__1613 (
            .O(N__11928),
            .I(N__11917));
    Span4Mux_s2_v I__1612 (
            .O(N__11925),
            .I(N__11914));
    InMux I__1611 (
            .O(N__11922),
            .I(N__11911));
    LocalMux I__1610 (
            .O(N__11917),
            .I(N__11908));
    Odrv4 I__1609 (
            .O(N__11914),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1608 (
            .O(N__11911),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__1607 (
            .O(N__11908),
            .I(\uu2.r_addrZ0Z_5 ));
    InMux I__1606 (
            .O(N__11901),
            .I(N__11898));
    LocalMux I__1605 (
            .O(N__11898),
            .I(\Lab_UT.dictrl.g1_5_0 ));
    InMux I__1604 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__1603 (
            .O(N__11892),
            .I(\Lab_UT.dictrl.N_97_mux_0 ));
    CascadeMux I__1602 (
            .O(N__11889),
            .I(\Lab_UT.dictrl.g0_16_2_cascade_ ));
    InMux I__1601 (
            .O(N__11886),
            .I(N__11883));
    LocalMux I__1600 (
            .O(N__11883),
            .I(N__11880));
    Span4Mux_v I__1599 (
            .O(N__11880),
            .I(N__11877));
    Odrv4 I__1598 (
            .O(N__11877),
            .I(\Lab_UT.dictrl.N_2446_1 ));
    CascadeMux I__1597 (
            .O(N__11874),
            .I(N__11871));
    InMux I__1596 (
            .O(N__11871),
            .I(N__11868));
    LocalMux I__1595 (
            .O(N__11868),
            .I(N__11865));
    Odrv4 I__1594 (
            .O(N__11865),
            .I(\uu2.mem0.w_addr_0 ));
    IoInMux I__1593 (
            .O(N__11862),
            .I(N__11859));
    LocalMux I__1592 (
            .O(N__11859),
            .I(N__11856));
    Span12Mux_s9_v I__1591 (
            .O(N__11856),
            .I(N__11852));
    InMux I__1590 (
            .O(N__11855),
            .I(N__11849));
    Odrv12 I__1589 (
            .O(N__11852),
            .I(clk));
    LocalMux I__1588 (
            .O(N__11849),
            .I(clk));
    SRMux I__1587 (
            .O(N__11844),
            .I(N__11841));
    LocalMux I__1586 (
            .O(N__11841),
            .I(N__11837));
    CEMux I__1585 (
            .O(N__11840),
            .I(N__11834));
    Span4Mux_h I__1584 (
            .O(N__11837),
            .I(N__11831));
    LocalMux I__1583 (
            .O(N__11834),
            .I(N__11828));
    Odrv4 I__1582 (
            .O(N__11831),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    Odrv4 I__1581 (
            .O(N__11828),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1580 (
            .O(N__11823),
            .I(N__11820));
    InMux I__1579 (
            .O(N__11820),
            .I(N__11817));
    LocalMux I__1578 (
            .O(N__11817),
            .I(N__11814));
    Odrv4 I__1577 (
            .O(N__11814),
            .I(\uu2.mem0.w_addr_1 ));
    CascadeMux I__1576 (
            .O(N__11811),
            .I(N__11808));
    InMux I__1575 (
            .O(N__11808),
            .I(N__11805));
    LocalMux I__1574 (
            .O(N__11805),
            .I(N__11802));
    Odrv12 I__1573 (
            .O(N__11802),
            .I(\uu2.mem0.w_addr_2 ));
    CascadeMux I__1572 (
            .O(N__11799),
            .I(\Lab_UT.dictrl.m40Z0Z_1_cascade_ ));
    InMux I__1571 (
            .O(N__11796),
            .I(N__11793));
    LocalMux I__1570 (
            .O(N__11793),
            .I(N__11790));
    Span4Mux_h I__1569 (
            .O(N__11790),
            .I(N__11787));
    Odrv4 I__1568 (
            .O(N__11787),
            .I(\Lab_UT.dictrl.N_10_3 ));
    CascadeMux I__1567 (
            .O(N__11784),
            .I(\Lab_UT.dictrl.N_5_0_cascade_ ));
    CascadeMux I__1566 (
            .O(N__11781),
            .I(N__11778));
    InMux I__1565 (
            .O(N__11778),
            .I(N__11775));
    LocalMux I__1564 (
            .O(N__11775),
            .I(\Lab_UT.dictrl.g0_9Z0Z_3 ));
    InMux I__1563 (
            .O(N__11772),
            .I(N__11769));
    LocalMux I__1562 (
            .O(N__11769),
            .I(N__11766));
    Odrv12 I__1561 (
            .O(N__11766),
            .I(\Lab_UT.dictrl.g1_4 ));
    CascadeMux I__1560 (
            .O(N__11763),
            .I(\Lab_UT.dictrl.N_97_mux_0_cascade_ ));
    InMux I__1559 (
            .O(N__11760),
            .I(N__11757));
    LocalMux I__1558 (
            .O(N__11757),
            .I(N__11754));
    Span4Mux_s3_h I__1557 (
            .O(N__11754),
            .I(N__11751));
    Odrv4 I__1556 (
            .O(N__11751),
            .I(\Lab_UT.dictrl.N_2435_0 ));
    InMux I__1555 (
            .O(N__11748),
            .I(N__11745));
    LocalMux I__1554 (
            .O(N__11745),
            .I(N__11742));
    Span4Mux_h I__1553 (
            .O(N__11742),
            .I(N__11737));
    InMux I__1552 (
            .O(N__11741),
            .I(N__11730));
    InMux I__1551 (
            .O(N__11740),
            .I(N__11730));
    Span4Mux_v I__1550 (
            .O(N__11737),
            .I(N__11727));
    InMux I__1549 (
            .O(N__11736),
            .I(N__11722));
    InMux I__1548 (
            .O(N__11735),
            .I(N__11722));
    LocalMux I__1547 (
            .O(N__11730),
            .I(N__11719));
    Odrv4 I__1546 (
            .O(N__11727),
            .I(buart__rx_hh_1));
    LocalMux I__1545 (
            .O(N__11722),
            .I(buart__rx_hh_1));
    Odrv4 I__1544 (
            .O(N__11719),
            .I(buart__rx_hh_1));
    CascadeMux I__1543 (
            .O(N__11712),
            .I(\Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_ ));
    InMux I__1542 (
            .O(N__11709),
            .I(N__11706));
    LocalMux I__1541 (
            .O(N__11706),
            .I(\Lab_UT.dictrl.g0_12_o6_2_2 ));
    CascadeMux I__1540 (
            .O(N__11703),
            .I(\Lab_UT.dictrl.N_13_0_cascade_ ));
    InMux I__1539 (
            .O(N__11700),
            .I(N__11697));
    LocalMux I__1538 (
            .O(N__11697),
            .I(\Lab_UT.dictrl.g0_10Z0Z_3 ));
    InMux I__1537 (
            .O(N__11694),
            .I(N__11691));
    LocalMux I__1536 (
            .O(N__11691),
            .I(\Lab_UT.dictrl.m34_4Z0Z_2 ));
    CascadeMux I__1535 (
            .O(N__11688),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    CascadeMux I__1534 (
            .O(N__11685),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ));
    CascadeMux I__1533 (
            .O(N__11682),
            .I(N__11677));
    InMux I__1532 (
            .O(N__11681),
            .I(N__11672));
    InMux I__1531 (
            .O(N__11680),
            .I(N__11672));
    InMux I__1530 (
            .O(N__11677),
            .I(N__11669));
    LocalMux I__1529 (
            .O(N__11672),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__1528 (
            .O(N__11669),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__1527 (
            .O(N__11664),
            .I(N__11660));
    InMux I__1526 (
            .O(N__11663),
            .I(N__11649));
    InMux I__1525 (
            .O(N__11660),
            .I(N__11649));
    InMux I__1524 (
            .O(N__11659),
            .I(N__11649));
    InMux I__1523 (
            .O(N__11658),
            .I(N__11649));
    LocalMux I__1522 (
            .O(N__11649),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__1521 (
            .O(N__11646),
            .I(N__11639));
    InMux I__1520 (
            .O(N__11645),
            .I(N__11636));
    InMux I__1519 (
            .O(N__11644),
            .I(N__11629));
    InMux I__1518 (
            .O(N__11643),
            .I(N__11629));
    InMux I__1517 (
            .O(N__11642),
            .I(N__11629));
    LocalMux I__1516 (
            .O(N__11639),
            .I(N__11626));
    LocalMux I__1515 (
            .O(N__11636),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__1514 (
            .O(N__11629),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    Odrv4 I__1513 (
            .O(N__11626),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    InMux I__1512 (
            .O(N__11619),
            .I(N__11604));
    InMux I__1511 (
            .O(N__11618),
            .I(N__11604));
    InMux I__1510 (
            .O(N__11617),
            .I(N__11604));
    InMux I__1509 (
            .O(N__11616),
            .I(N__11604));
    InMux I__1508 (
            .O(N__11615),
            .I(N__11604));
    LocalMux I__1507 (
            .O(N__11604),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__1506 (
            .O(N__11601),
            .I(N__11588));
    InMux I__1505 (
            .O(N__11600),
            .I(N__11588));
    InMux I__1504 (
            .O(N__11599),
            .I(N__11588));
    InMux I__1503 (
            .O(N__11598),
            .I(N__11578));
    InMux I__1502 (
            .O(N__11597),
            .I(N__11578));
    InMux I__1501 (
            .O(N__11596),
            .I(N__11573));
    InMux I__1500 (
            .O(N__11595),
            .I(N__11573));
    LocalMux I__1499 (
            .O(N__11588),
            .I(N__11570));
    InMux I__1498 (
            .O(N__11587),
            .I(N__11563));
    InMux I__1497 (
            .O(N__11586),
            .I(N__11563));
    InMux I__1496 (
            .O(N__11585),
            .I(N__11563));
    InMux I__1495 (
            .O(N__11584),
            .I(N__11558));
    InMux I__1494 (
            .O(N__11583),
            .I(N__11558));
    LocalMux I__1493 (
            .O(N__11578),
            .I(N__11555));
    LocalMux I__1492 (
            .O(N__11573),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1491 (
            .O(N__11570),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1490 (
            .O(N__11563),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1489 (
            .O(N__11558),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1488 (
            .O(N__11555),
            .I(\uu0.un4_l_count_0 ));
    IoInMux I__1487 (
            .O(N__11544),
            .I(N__11541));
    LocalMux I__1486 (
            .O(N__11541),
            .I(N__11538));
    IoSpan4Mux I__1485 (
            .O(N__11538),
            .I(N__11535));
    Span4Mux_s0_h I__1484 (
            .O(N__11535),
            .I(N__11532));
    Odrv4 I__1483 (
            .O(N__11532),
            .I(\uu0.un11_l_count_i ));
    InMux I__1482 (
            .O(N__11529),
            .I(N__11523));
    InMux I__1481 (
            .O(N__11528),
            .I(N__11523));
    LocalMux I__1480 (
            .O(N__11523),
            .I(N__11520));
    Span4Mux_h I__1479 (
            .O(N__11520),
            .I(N__11517));
    Odrv4 I__1478 (
            .O(N__11517),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__1477 (
            .O(N__11514),
            .I(N__11511));
    LocalMux I__1476 (
            .O(N__11511),
            .I(\uu0.delay_lineZ0Z_1 ));
    CascadeMux I__1475 (
            .O(N__11508),
            .I(\buart.Z_tx.un1_bitcount_c3_cascade_ ));
    InMux I__1474 (
            .O(N__11505),
            .I(N__11499));
    InMux I__1473 (
            .O(N__11504),
            .I(N__11499));
    LocalMux I__1472 (
            .O(N__11499),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__1471 (
            .O(N__11496),
            .I(N__11493));
    LocalMux I__1470 (
            .O(N__11493),
            .I(\buart.Z_tx.uart_busy_0_0 ));
    InMux I__1469 (
            .O(N__11490),
            .I(N__11484));
    InMux I__1468 (
            .O(N__11489),
            .I(N__11477));
    InMux I__1467 (
            .O(N__11488),
            .I(N__11477));
    InMux I__1466 (
            .O(N__11487),
            .I(N__11477));
    LocalMux I__1465 (
            .O(N__11484),
            .I(N__11474));
    LocalMux I__1464 (
            .O(N__11477),
            .I(\buart.Z_tx.ser_clk ));
    Odrv4 I__1463 (
            .O(N__11474),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__1462 (
            .O(N__11469),
            .I(N__11466));
    InMux I__1461 (
            .O(N__11466),
            .I(N__11463));
    LocalMux I__1460 (
            .O(N__11463),
            .I(\uu2.un1_l_count_1_2_0 ));
    InMux I__1459 (
            .O(N__11460),
            .I(N__11455));
    InMux I__1458 (
            .O(N__11459),
            .I(N__11452));
    InMux I__1457 (
            .O(N__11458),
            .I(N__11449));
    LocalMux I__1456 (
            .O(N__11455),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__1455 (
            .O(N__11452),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__1454 (
            .O(N__11449),
            .I(\uu2.l_countZ0Z_5 ));
    CascadeMux I__1453 (
            .O(N__11442),
            .I(\uu2.vbuf_count.un328_ci_3_cascade_ ));
    InMux I__1452 (
            .O(N__11439),
            .I(N__11436));
    LocalMux I__1451 (
            .O(N__11436),
            .I(N__11431));
    InMux I__1450 (
            .O(N__11435),
            .I(N__11428));
    InMux I__1449 (
            .O(N__11434),
            .I(N__11425));
    Span4Mux_s3_h I__1448 (
            .O(N__11431),
            .I(N__11422));
    LocalMux I__1447 (
            .O(N__11428),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__1446 (
            .O(N__11425),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__1445 (
            .O(N__11422),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__1444 (
            .O(N__11415),
            .I(\uu2.un350_ci_cascade_ ));
    CascadeMux I__1443 (
            .O(N__11412),
            .I(N__11405));
    InMux I__1442 (
            .O(N__11411),
            .I(N__11400));
    InMux I__1441 (
            .O(N__11410),
            .I(N__11400));
    InMux I__1440 (
            .O(N__11409),
            .I(N__11393));
    InMux I__1439 (
            .O(N__11408),
            .I(N__11393));
    InMux I__1438 (
            .O(N__11405),
            .I(N__11393));
    LocalMux I__1437 (
            .O(N__11400),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__1436 (
            .O(N__11393),
            .I(\uu2.l_countZ0Z_4 ));
    CascadeMux I__1435 (
            .O(N__11388),
            .I(N__11383));
    InMux I__1434 (
            .O(N__11387),
            .I(N__11376));
    InMux I__1433 (
            .O(N__11386),
            .I(N__11376));
    InMux I__1432 (
            .O(N__11383),
            .I(N__11376));
    LocalMux I__1431 (
            .O(N__11376),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__1430 (
            .O(N__11373),
            .I(N__11370));
    LocalMux I__1429 (
            .O(N__11370),
            .I(\uu2.un1_l_count_2_2 ));
    CascadeMux I__1428 (
            .O(N__11367),
            .I(N__11364));
    InMux I__1427 (
            .O(N__11364),
            .I(N__11358));
    InMux I__1426 (
            .O(N__11363),
            .I(N__11351));
    InMux I__1425 (
            .O(N__11362),
            .I(N__11351));
    InMux I__1424 (
            .O(N__11361),
            .I(N__11351));
    LocalMux I__1423 (
            .O(N__11358),
            .I(\uu2.un306_ci ));
    LocalMux I__1422 (
            .O(N__11351),
            .I(\uu2.un306_ci ));
    InMux I__1421 (
            .O(N__11346),
            .I(N__11340));
    InMux I__1420 (
            .O(N__11345),
            .I(N__11340));
    LocalMux I__1419 (
            .O(N__11340),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    CascadeMux I__1418 (
            .O(N__11337),
            .I(N__11334));
    InMux I__1417 (
            .O(N__11334),
            .I(N__11319));
    InMux I__1416 (
            .O(N__11333),
            .I(N__11319));
    InMux I__1415 (
            .O(N__11332),
            .I(N__11319));
    InMux I__1414 (
            .O(N__11331),
            .I(N__11319));
    InMux I__1413 (
            .O(N__11330),
            .I(N__11319));
    LocalMux I__1412 (
            .O(N__11319),
            .I(\uu2.l_countZ0Z_6 ));
    InMux I__1411 (
            .O(N__11316),
            .I(N__11309));
    InMux I__1410 (
            .O(N__11315),
            .I(N__11309));
    InMux I__1409 (
            .O(N__11314),
            .I(N__11306));
    LocalMux I__1408 (
            .O(N__11309),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__1407 (
            .O(N__11306),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__1406 (
            .O(N__11301),
            .I(N__11298));
    LocalMux I__1405 (
            .O(N__11298),
            .I(\uu2.un350_ci ));
    InMux I__1404 (
            .O(N__11295),
            .I(N__11290));
    InMux I__1403 (
            .O(N__11294),
            .I(N__11287));
    InMux I__1402 (
            .O(N__11293),
            .I(N__11284));
    LocalMux I__1401 (
            .O(N__11290),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1400 (
            .O(N__11287),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__1399 (
            .O(N__11284),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__1398 (
            .O(N__11277),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    CascadeMux I__1397 (
            .O(N__11274),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__1396 (
            .O(N__11271),
            .I(N__11268));
    LocalMux I__1395 (
            .O(N__11268),
            .I(\uu2.un1_l_count_1_3 ));
    CascadeMux I__1394 (
            .O(N__11265),
            .I(N__11260));
    InMux I__1393 (
            .O(N__11264),
            .I(N__11255));
    InMux I__1392 (
            .O(N__11263),
            .I(N__11255));
    InMux I__1391 (
            .O(N__11260),
            .I(N__11252));
    LocalMux I__1390 (
            .O(N__11255),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__1389 (
            .O(N__11252),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__1388 (
            .O(N__11247),
            .I(N__11240));
    InMux I__1387 (
            .O(N__11246),
            .I(N__11229));
    InMux I__1386 (
            .O(N__11245),
            .I(N__11229));
    InMux I__1385 (
            .O(N__11244),
            .I(N__11229));
    InMux I__1384 (
            .O(N__11243),
            .I(N__11229));
    InMux I__1383 (
            .O(N__11240),
            .I(N__11229));
    LocalMux I__1382 (
            .O(N__11229),
            .I(\uu2.l_countZ0Z_2 ));
    CascadeMux I__1381 (
            .O(N__11226),
            .I(\uu2.un306_ci_cascade_ ));
    CascadeMux I__1380 (
            .O(N__11223),
            .I(\uu2.un404_ci_0_cascade_ ));
    CascadeMux I__1379 (
            .O(N__11220),
            .I(N__11217));
    InMux I__1378 (
            .O(N__11217),
            .I(N__11211));
    InMux I__1377 (
            .O(N__11216),
            .I(N__11204));
    InMux I__1376 (
            .O(N__11215),
            .I(N__11204));
    InMux I__1375 (
            .O(N__11214),
            .I(N__11204));
    LocalMux I__1374 (
            .O(N__11211),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1373 (
            .O(N__11204),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1372 (
            .O(N__11199),
            .I(N__11194));
    CascadeMux I__1371 (
            .O(N__11198),
            .I(N__11191));
    CascadeMux I__1370 (
            .O(N__11197),
            .I(N__11188));
    InMux I__1369 (
            .O(N__11194),
            .I(N__11185));
    InMux I__1368 (
            .O(N__11191),
            .I(N__11180));
    InMux I__1367 (
            .O(N__11188),
            .I(N__11180));
    LocalMux I__1366 (
            .O(N__11185),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1365 (
            .O(N__11180),
            .I(\uu2.r_addrZ0Z_3 ));
    CascadeMux I__1364 (
            .O(N__11175),
            .I(N__11171));
    CascadeMux I__1363 (
            .O(N__11174),
            .I(N__11168));
    InMux I__1362 (
            .O(N__11171),
            .I(N__11163));
    InMux I__1361 (
            .O(N__11168),
            .I(N__11160));
    InMux I__1360 (
            .O(N__11167),
            .I(N__11155));
    InMux I__1359 (
            .O(N__11166),
            .I(N__11155));
    LocalMux I__1358 (
            .O(N__11163),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1357 (
            .O(N__11160),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1356 (
            .O(N__11155),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1355 (
            .O(N__11148),
            .I(N__11145));
    InMux I__1354 (
            .O(N__11145),
            .I(N__11142));
    LocalMux I__1353 (
            .O(N__11142),
            .I(N__11135));
    InMux I__1352 (
            .O(N__11141),
            .I(N__11130));
    InMux I__1351 (
            .O(N__11140),
            .I(N__11130));
    InMux I__1350 (
            .O(N__11139),
            .I(N__11125));
    InMux I__1349 (
            .O(N__11138),
            .I(N__11125));
    Odrv4 I__1348 (
            .O(N__11135),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1347 (
            .O(N__11130),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1346 (
            .O(N__11125),
            .I(\uu2.r_addrZ0Z_1 ));
    CEMux I__1345 (
            .O(N__11118),
            .I(N__11115));
    LocalMux I__1344 (
            .O(N__11115),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__1343 (
            .O(N__11112),
            .I(\uu2.trig_rd_is_det_cascade_ ));
    CascadeMux I__1342 (
            .O(N__11109),
            .I(N__11105));
    CascadeMux I__1341 (
            .O(N__11108),
            .I(N__11101));
    InMux I__1340 (
            .O(N__11105),
            .I(N__11095));
    InMux I__1339 (
            .O(N__11104),
            .I(N__11088));
    InMux I__1338 (
            .O(N__11101),
            .I(N__11088));
    InMux I__1337 (
            .O(N__11100),
            .I(N__11088));
    InMux I__1336 (
            .O(N__11099),
            .I(N__11083));
    InMux I__1335 (
            .O(N__11098),
            .I(N__11083));
    LocalMux I__1334 (
            .O(N__11095),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1333 (
            .O(N__11088),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1332 (
            .O(N__11083),
            .I(\uu2.r_addrZ0Z_0 ));
    InMux I__1331 (
            .O(N__11076),
            .I(N__11073));
    LocalMux I__1330 (
            .O(N__11073),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1329 (
            .O(N__11070),
            .I(N__11064));
    InMux I__1328 (
            .O(N__11069),
            .I(N__11064));
    LocalMux I__1327 (
            .O(N__11064),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    CascadeMux I__1326 (
            .O(N__11061),
            .I(N__11058));
    InMux I__1325 (
            .O(N__11058),
            .I(N__11055));
    LocalMux I__1324 (
            .O(N__11055),
            .I(N__11052));
    Odrv4 I__1323 (
            .O(N__11052),
            .I(\Lab_UT.dictrl.g1_6_0 ));
    InMux I__1322 (
            .O(N__11049),
            .I(N__11046));
    LocalMux I__1321 (
            .O(N__11046),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__1320 (
            .O(N__11043),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1319 (
            .O(N__11040),
            .I(N__11037));
    InMux I__1318 (
            .O(N__11037),
            .I(N__11033));
    InMux I__1317 (
            .O(N__11036),
            .I(N__11030));
    LocalMux I__1316 (
            .O(N__11033),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1315 (
            .O(N__11030),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__1314 (
            .O(N__11025),
            .I(N__11021));
    CascadeMux I__1313 (
            .O(N__11024),
            .I(N__11018));
    InMux I__1312 (
            .O(N__11021),
            .I(N__11014));
    InMux I__1311 (
            .O(N__11018),
            .I(N__11009));
    InMux I__1310 (
            .O(N__11017),
            .I(N__11009));
    LocalMux I__1309 (
            .O(N__11014),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1308 (
            .O(N__11009),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__1307 (
            .O(N__11004),
            .I(N__11001));
    LocalMux I__1306 (
            .O(N__11001),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    CascadeMux I__1305 (
            .O(N__10998),
            .I(\Lab_UT.dictrl.N_1792_1_cascade_ ));
    InMux I__1304 (
            .O(N__10995),
            .I(N__10992));
    LocalMux I__1303 (
            .O(N__10992),
            .I(\Lab_UT.dictrl.N_1451_0 ));
    CascadeMux I__1302 (
            .O(N__10989),
            .I(\Lab_UT.dictrl.g0_i_a5_2_4_cascade_ ));
    InMux I__1301 (
            .O(N__10986),
            .I(N__10983));
    LocalMux I__1300 (
            .O(N__10983),
            .I(\Lab_UT.dictrl.g0_i_a5_2_5 ));
    CascadeMux I__1299 (
            .O(N__10980),
            .I(N__10977));
    InMux I__1298 (
            .O(N__10977),
            .I(N__10974));
    LocalMux I__1297 (
            .O(N__10974),
            .I(\Lab_UT.dictrl.g0_5_3 ));
    InMux I__1296 (
            .O(N__10971),
            .I(N__10968));
    LocalMux I__1295 (
            .O(N__10968),
            .I(N__10965));
    Odrv4 I__1294 (
            .O(N__10965),
            .I(\Lab_UT.dictrl.g0_5_4 ));
    CascadeMux I__1293 (
            .O(N__10962),
            .I(\Lab_UT.dictrl.g0_69_1_cascade_ ));
    InMux I__1292 (
            .O(N__10959),
            .I(N__10956));
    LocalMux I__1291 (
            .O(N__10956),
            .I(\Lab_UT.dictrl.g1_0_3_1 ));
    CascadeMux I__1290 (
            .O(N__10953),
            .I(\Lab_UT.dictrl.g1_5_1_cascade_ ));
    InMux I__1289 (
            .O(N__10950),
            .I(N__10947));
    LocalMux I__1288 (
            .O(N__10947),
            .I(\Lab_UT.dictrl.N_61_1 ));
    InMux I__1287 (
            .O(N__10944),
            .I(N__10941));
    LocalMux I__1286 (
            .O(N__10941),
            .I(\Lab_UT.dictrl.g1_7_0 ));
    InMux I__1285 (
            .O(N__10938),
            .I(N__10935));
    LocalMux I__1284 (
            .O(N__10935),
            .I(N_107));
    CascadeMux I__1283 (
            .O(N__10932),
            .I(m72_cascade_));
    InMux I__1282 (
            .O(N__10929),
            .I(N__10923));
    InMux I__1281 (
            .O(N__10928),
            .I(N__10923));
    LocalMux I__1280 (
            .O(N__10923),
            .I(N_105));
    InMux I__1279 (
            .O(N__10920),
            .I(N__10914));
    InMux I__1278 (
            .O(N__10919),
            .I(N__10914));
    LocalMux I__1277 (
            .O(N__10914),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__1276 (
            .O(N__10911),
            .I(N__10906));
    InMux I__1275 (
            .O(N__10910),
            .I(N__10898));
    InMux I__1274 (
            .O(N__10909),
            .I(N__10898));
    InMux I__1273 (
            .O(N__10906),
            .I(N__10891));
    InMux I__1272 (
            .O(N__10905),
            .I(N__10891));
    InMux I__1271 (
            .O(N__10904),
            .I(N__10891));
    InMux I__1270 (
            .O(N__10903),
            .I(N__10888));
    LocalMux I__1269 (
            .O(N__10898),
            .I(resetGen_reset_count_4));
    LocalMux I__1268 (
            .O(N__10891),
            .I(resetGen_reset_count_4));
    LocalMux I__1267 (
            .O(N__10888),
            .I(resetGen_reset_count_4));
    CascadeMux I__1266 (
            .O(N__10881),
            .I(N__10876));
    CascadeMux I__1265 (
            .O(N__10880),
            .I(N__10872));
    CascadeMux I__1264 (
            .O(N__10879),
            .I(N__10869));
    InMux I__1263 (
            .O(N__10876),
            .I(N__10863));
    InMux I__1262 (
            .O(N__10875),
            .I(N__10863));
    InMux I__1261 (
            .O(N__10872),
            .I(N__10856));
    InMux I__1260 (
            .O(N__10869),
            .I(N__10856));
    InMux I__1259 (
            .O(N__10868),
            .I(N__10856));
    LocalMux I__1258 (
            .O(N__10863),
            .I(resetGen_reset_count_0));
    LocalMux I__1257 (
            .O(N__10856),
            .I(resetGen_reset_count_0));
    InMux I__1256 (
            .O(N__10851),
            .I(N__10848));
    LocalMux I__1255 (
            .O(N__10848),
            .I(N__10843));
    InMux I__1254 (
            .O(N__10847),
            .I(N__10838));
    InMux I__1253 (
            .O(N__10846),
            .I(N__10838));
    Odrv4 I__1252 (
            .O(N__10843),
            .I(buart__rx_hh_0));
    LocalMux I__1251 (
            .O(N__10838),
            .I(buart__rx_hh_0));
    InMux I__1250 (
            .O(N__10833),
            .I(N__10830));
    LocalMux I__1249 (
            .O(N__10830),
            .I(N__10827));
    Odrv12 I__1248 (
            .O(N__10827),
            .I(vbuf_tx_data_6));
    InMux I__1247 (
            .O(N__10824),
            .I(N__10821));
    LocalMux I__1246 (
            .O(N__10821),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__1245 (
            .O(N__10818),
            .I(N__10815));
    LocalMux I__1244 (
            .O(N__10815),
            .I(N__10812));
    Odrv12 I__1243 (
            .O(N__10812),
            .I(vbuf_tx_data_7));
    InMux I__1242 (
            .O(N__10809),
            .I(N__10806));
    LocalMux I__1241 (
            .O(N__10806),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__1240 (
            .O(N__10803),
            .I(N__10800));
    LocalMux I__1239 (
            .O(N__10800),
            .I(N__10797));
    Span4Mux_s1_v I__1238 (
            .O(N__10797),
            .I(N__10793));
    CEMux I__1237 (
            .O(N__10796),
            .I(N__10790));
    Odrv4 I__1236 (
            .O(N__10793),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    LocalMux I__1235 (
            .O(N__10790),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1234 (
            .O(N__10785),
            .I(N__10781));
    InMux I__1233 (
            .O(N__10784),
            .I(N__10778));
    LocalMux I__1232 (
            .O(N__10781),
            .I(\uu0.l_countZ0Z_13 ));
    LocalMux I__1231 (
            .O(N__10778),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__1230 (
            .O(N__10773),
            .I(N__10767));
    InMux I__1229 (
            .O(N__10772),
            .I(N__10760));
    InMux I__1228 (
            .O(N__10771),
            .I(N__10760));
    InMux I__1227 (
            .O(N__10770),
            .I(N__10760));
    LocalMux I__1226 (
            .O(N__10767),
            .I(N__10757));
    LocalMux I__1225 (
            .O(N__10760),
            .I(N__10752));
    Span4Mux_s1_h I__1224 (
            .O(N__10757),
            .I(N__10752));
    Odrv4 I__1223 (
            .O(N__10752),
            .I(\uu0.un4_l_count_0_8 ));
    InMux I__1222 (
            .O(N__10749),
            .I(N__10746));
    LocalMux I__1221 (
            .O(N__10746),
            .I(N__10740));
    CascadeMux I__1220 (
            .O(N__10745),
            .I(N__10737));
    CascadeMux I__1219 (
            .O(N__10744),
            .I(N__10734));
    InMux I__1218 (
            .O(N__10743),
            .I(N__10731));
    Span4Mux_h I__1217 (
            .O(N__10740),
            .I(N__10728));
    InMux I__1216 (
            .O(N__10737),
            .I(N__10723));
    InMux I__1215 (
            .O(N__10734),
            .I(N__10723));
    LocalMux I__1214 (
            .O(N__10731),
            .I(\uu0.un154_ci_9 ));
    Odrv4 I__1213 (
            .O(N__10728),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__1212 (
            .O(N__10723),
            .I(\uu0.un154_ci_9 ));
    InMux I__1211 (
            .O(N__10716),
            .I(N__10709));
    InMux I__1210 (
            .O(N__10715),
            .I(N__10709));
    InMux I__1209 (
            .O(N__10714),
            .I(N__10706));
    LocalMux I__1208 (
            .O(N__10709),
            .I(N__10703));
    LocalMux I__1207 (
            .O(N__10706),
            .I(\uu0.l_countZ0Z_12 ));
    Odrv4 I__1206 (
            .O(N__10703),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__1205 (
            .O(N__10698),
            .I(N__10695));
    LocalMux I__1204 (
            .O(N__10695),
            .I(\uu0.un165_ci_0 ));
    InMux I__1203 (
            .O(N__10692),
            .I(N__10686));
    InMux I__1202 (
            .O(N__10691),
            .I(N__10679));
    InMux I__1201 (
            .O(N__10690),
            .I(N__10679));
    InMux I__1200 (
            .O(N__10689),
            .I(N__10679));
    LocalMux I__1199 (
            .O(N__10686),
            .I(resetGen_reset_count_1));
    LocalMux I__1198 (
            .O(N__10679),
            .I(resetGen_reset_count_1));
    InMux I__1197 (
            .O(N__10674),
            .I(N__10671));
    LocalMux I__1196 (
            .O(N__10671),
            .I(\uu0.un44_ci ));
    CascadeMux I__1195 (
            .O(N__10668),
            .I(N__10665));
    InMux I__1194 (
            .O(N__10665),
            .I(N__10662));
    LocalMux I__1193 (
            .O(N__10662),
            .I(N__10656));
    InMux I__1192 (
            .O(N__10661),
            .I(N__10651));
    InMux I__1191 (
            .O(N__10660),
            .I(N__10651));
    InMux I__1190 (
            .O(N__10659),
            .I(N__10648));
    Odrv4 I__1189 (
            .O(N__10656),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__1188 (
            .O(N__10651),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__1187 (
            .O(N__10648),
            .I(\uu0.l_countZ0Z_2 ));
    InMux I__1186 (
            .O(N__10641),
            .I(N__10636));
    InMux I__1185 (
            .O(N__10640),
            .I(N__10631));
    InMux I__1184 (
            .O(N__10639),
            .I(N__10631));
    LocalMux I__1183 (
            .O(N__10636),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__1182 (
            .O(N__10631),
            .I(\uu0.l_countZ0Z_3 ));
    CascadeMux I__1181 (
            .O(N__10626),
            .I(N__10620));
    CascadeMux I__1180 (
            .O(N__10625),
            .I(N__10617));
    InMux I__1179 (
            .O(N__10624),
            .I(N__10614));
    InMux I__1178 (
            .O(N__10623),
            .I(N__10611));
    InMux I__1177 (
            .O(N__10620),
            .I(N__10608));
    InMux I__1176 (
            .O(N__10617),
            .I(N__10605));
    LocalMux I__1175 (
            .O(N__10614),
            .I(\uu0.un66_ci ));
    LocalMux I__1174 (
            .O(N__10611),
            .I(\uu0.un66_ci ));
    LocalMux I__1173 (
            .O(N__10608),
            .I(\uu0.un66_ci ));
    LocalMux I__1172 (
            .O(N__10605),
            .I(\uu0.un66_ci ));
    InMux I__1171 (
            .O(N__10596),
            .I(N__10591));
    InMux I__1170 (
            .O(N__10595),
            .I(N__10586));
    InMux I__1169 (
            .O(N__10594),
            .I(N__10586));
    LocalMux I__1168 (
            .O(N__10591),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__1167 (
            .O(N__10586),
            .I(\uu0.l_countZ0Z_7 ));
    InMux I__1166 (
            .O(N__10581),
            .I(N__10578));
    LocalMux I__1165 (
            .O(N__10578),
            .I(\uu0.un220_ci ));
    CascadeMux I__1164 (
            .O(N__10575),
            .I(N__10572));
    InMux I__1163 (
            .O(N__10572),
            .I(N__10569));
    LocalMux I__1162 (
            .O(N__10569),
            .I(\uu0.un143_ci_0 ));
    CascadeMux I__1161 (
            .O(N__10566),
            .I(N__10563));
    InMux I__1160 (
            .O(N__10563),
            .I(N__10558));
    InMux I__1159 (
            .O(N__10562),
            .I(N__10553));
    InMux I__1158 (
            .O(N__10561),
            .I(N__10553));
    LocalMux I__1157 (
            .O(N__10558),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__1156 (
            .O(N__10553),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__1155 (
            .O(N__10548),
            .I(N__10544));
    CascadeMux I__1154 (
            .O(N__10547),
            .I(N__10541));
    InMux I__1153 (
            .O(N__10544),
            .I(N__10536));
    InMux I__1152 (
            .O(N__10541),
            .I(N__10536));
    LocalMux I__1151 (
            .O(N__10536),
            .I(\uu0.l_countZ0Z_18 ));
    InMux I__1150 (
            .O(N__10533),
            .I(N__10530));
    LocalMux I__1149 (
            .O(N__10530),
            .I(\uu0.un4_l_count_11 ));
    InMux I__1148 (
            .O(N__10527),
            .I(N__10524));
    LocalMux I__1147 (
            .O(N__10524),
            .I(N__10521));
    Odrv4 I__1146 (
            .O(N__10521),
            .I(\uu0.un4_l_count_12 ));
    InMux I__1145 (
            .O(N__10518),
            .I(N__10515));
    LocalMux I__1144 (
            .O(N__10515),
            .I(\uu0.un4_l_count_13 ));
    CascadeMux I__1143 (
            .O(N__10512),
            .I(\uu0.un4_l_count_16_cascade_ ));
    InMux I__1142 (
            .O(N__10509),
            .I(N__10506));
    LocalMux I__1141 (
            .O(N__10506),
            .I(N__10503));
    Odrv4 I__1140 (
            .O(N__10503),
            .I(\uu0.un4_l_count_18 ));
    InMux I__1139 (
            .O(N__10500),
            .I(N__10489));
    InMux I__1138 (
            .O(N__10499),
            .I(N__10489));
    CascadeMux I__1137 (
            .O(N__10498),
            .I(N__10484));
    CascadeMux I__1136 (
            .O(N__10497),
            .I(N__10481));
    InMux I__1135 (
            .O(N__10496),
            .I(N__10477));
    InMux I__1134 (
            .O(N__10495),
            .I(N__10472));
    InMux I__1133 (
            .O(N__10494),
            .I(N__10472));
    LocalMux I__1132 (
            .O(N__10489),
            .I(N__10469));
    InMux I__1131 (
            .O(N__10488),
            .I(N__10466));
    InMux I__1130 (
            .O(N__10487),
            .I(N__10457));
    InMux I__1129 (
            .O(N__10484),
            .I(N__10457));
    InMux I__1128 (
            .O(N__10481),
            .I(N__10457));
    InMux I__1127 (
            .O(N__10480),
            .I(N__10457));
    LocalMux I__1126 (
            .O(N__10477),
            .I(\uu0.un110_ci ));
    LocalMux I__1125 (
            .O(N__10472),
            .I(\uu0.un110_ci ));
    Odrv12 I__1124 (
            .O(N__10469),
            .I(\uu0.un110_ci ));
    LocalMux I__1123 (
            .O(N__10466),
            .I(\uu0.un110_ci ));
    LocalMux I__1122 (
            .O(N__10457),
            .I(\uu0.un110_ci ));
    CascadeMux I__1121 (
            .O(N__10446),
            .I(\uu0.un4_l_count_0_cascade_ ));
    CEMux I__1120 (
            .O(N__10443),
            .I(N__10428));
    CEMux I__1119 (
            .O(N__10442),
            .I(N__10428));
    CEMux I__1118 (
            .O(N__10441),
            .I(N__10428));
    CEMux I__1117 (
            .O(N__10440),
            .I(N__10428));
    CEMux I__1116 (
            .O(N__10439),
            .I(N__10428));
    GlobalMux I__1115 (
            .O(N__10428),
            .I(N__10425));
    gio2CtrlBuf I__1114 (
            .O(N__10425),
            .I(\uu0.un11_l_count_i_g ));
    InMux I__1113 (
            .O(N__10422),
            .I(N__10419));
    LocalMux I__1112 (
            .O(N__10419),
            .I(N__10416));
    Odrv12 I__1111 (
            .O(N__10416),
            .I(vbuf_tx_data_5));
    InMux I__1110 (
            .O(N__10413),
            .I(N__10410));
    LocalMux I__1109 (
            .O(N__10410),
            .I(N__10407));
    Odrv12 I__1108 (
            .O(N__10407),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__1107 (
            .O(N__10404),
            .I(N__10391));
    InMux I__1106 (
            .O(N__10403),
            .I(N__10391));
    InMux I__1105 (
            .O(N__10402),
            .I(N__10391));
    InMux I__1104 (
            .O(N__10401),
            .I(N__10391));
    InMux I__1103 (
            .O(N__10400),
            .I(N__10388));
    LocalMux I__1102 (
            .O(N__10391),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__1101 (
            .O(N__10388),
            .I(\uu0.l_countZ0Z_0 ));
    CascadeMux I__1100 (
            .O(N__10383),
            .I(N__10378));
    InMux I__1099 (
            .O(N__10382),
            .I(N__10370));
    InMux I__1098 (
            .O(N__10381),
            .I(N__10370));
    InMux I__1097 (
            .O(N__10378),
            .I(N__10370));
    InMux I__1096 (
            .O(N__10377),
            .I(N__10367));
    LocalMux I__1095 (
            .O(N__10370),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__1094 (
            .O(N__10367),
            .I(\uu0.l_countZ0Z_1 ));
    CascadeMux I__1093 (
            .O(N__10362),
            .I(\uu0.un66_ci_cascade_ ));
    CascadeMux I__1092 (
            .O(N__10359),
            .I(\uu0.un110_ci_cascade_ ));
    InMux I__1091 (
            .O(N__10356),
            .I(N__10350));
    InMux I__1090 (
            .O(N__10355),
            .I(N__10345));
    InMux I__1089 (
            .O(N__10354),
            .I(N__10345));
    InMux I__1088 (
            .O(N__10353),
            .I(N__10342));
    LocalMux I__1087 (
            .O(N__10350),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__1086 (
            .O(N__10345),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__1085 (
            .O(N__10342),
            .I(\uu0.l_countZ0Z_10 ));
    CascadeMux I__1084 (
            .O(N__10335),
            .I(N__10330));
    InMux I__1083 (
            .O(N__10334),
            .I(N__10323));
    InMux I__1082 (
            .O(N__10333),
            .I(N__10323));
    InMux I__1081 (
            .O(N__10330),
            .I(N__10318));
    InMux I__1080 (
            .O(N__10329),
            .I(N__10318));
    InMux I__1079 (
            .O(N__10328),
            .I(N__10314));
    LocalMux I__1078 (
            .O(N__10323),
            .I(N__10311));
    LocalMux I__1077 (
            .O(N__10318),
            .I(N__10308));
    InMux I__1076 (
            .O(N__10317),
            .I(N__10305));
    LocalMux I__1075 (
            .O(N__10314),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1074 (
            .O(N__10311),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__1073 (
            .O(N__10308),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1072 (
            .O(N__10305),
            .I(\uu0.l_countZ0Z_8 ));
    InMux I__1071 (
            .O(N__10296),
            .I(N__10287));
    InMux I__1070 (
            .O(N__10295),
            .I(N__10287));
    InMux I__1069 (
            .O(N__10294),
            .I(N__10280));
    InMux I__1068 (
            .O(N__10293),
            .I(N__10280));
    InMux I__1067 (
            .O(N__10292),
            .I(N__10280));
    LocalMux I__1066 (
            .O(N__10287),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1065 (
            .O(N__10280),
            .I(\uu0.l_countZ0Z_9 ));
    CascadeMux I__1064 (
            .O(N__10275),
            .I(N__10270));
    InMux I__1063 (
            .O(N__10274),
            .I(N__10263));
    InMux I__1062 (
            .O(N__10273),
            .I(N__10263));
    InMux I__1061 (
            .O(N__10270),
            .I(N__10263));
    LocalMux I__1060 (
            .O(N__10263),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__1059 (
            .O(N__10260),
            .I(N__10255));
    InMux I__1058 (
            .O(N__10259),
            .I(N__10248));
    InMux I__1057 (
            .O(N__10258),
            .I(N__10248));
    InMux I__1056 (
            .O(N__10255),
            .I(N__10248));
    LocalMux I__1055 (
            .O(N__10248),
            .I(\uu0.un198_ci_2 ));
    InMux I__1054 (
            .O(N__10245),
            .I(N__10235));
    InMux I__1053 (
            .O(N__10244),
            .I(N__10235));
    InMux I__1052 (
            .O(N__10243),
            .I(N__10235));
    InMux I__1051 (
            .O(N__10242),
            .I(N__10232));
    LocalMux I__1050 (
            .O(N__10235),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1049 (
            .O(N__10232),
            .I(\uu0.l_countZ0Z_16 ));
    InMux I__1048 (
            .O(N__10227),
            .I(N__10224));
    LocalMux I__1047 (
            .O(N__10224),
            .I(vbuf_tx_data_1));
    InMux I__1046 (
            .O(N__10221),
            .I(N__10218));
    LocalMux I__1045 (
            .O(N__10218),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__1044 (
            .O(N__10215),
            .I(N__10212));
    LocalMux I__1043 (
            .O(N__10212),
            .I(vbuf_tx_data_2));
    InMux I__1042 (
            .O(N__10209),
            .I(N__10206));
    LocalMux I__1041 (
            .O(N__10206),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__1040 (
            .O(N__10203),
            .I(N__10200));
    LocalMux I__1039 (
            .O(N__10200),
            .I(vbuf_tx_data_3));
    InMux I__1038 (
            .O(N__10197),
            .I(N__10194));
    LocalMux I__1037 (
            .O(N__10194),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1036 (
            .O(N__10191),
            .I(N__10188));
    LocalMux I__1035 (
            .O(N__10188),
            .I(vbuf_tx_data_4));
    InMux I__1034 (
            .O(N__10185),
            .I(N__10182));
    LocalMux I__1033 (
            .O(N__10182),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    CascadeMux I__1032 (
            .O(N__10179),
            .I(\uu0.un44_ci_cascade_ ));
    InMux I__1031 (
            .O(N__10176),
            .I(N__10173));
    LocalMux I__1030 (
            .O(N__10173),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1029 (
            .O(N__10170),
            .I(N__10167));
    LocalMux I__1028 (
            .O(N__10167),
            .I(\uu2.r_data_wire_3 ));
    InMux I__1027 (
            .O(N__10164),
            .I(N__10161));
    LocalMux I__1026 (
            .O(N__10161),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1025 (
            .O(N__10158),
            .I(N__10155));
    LocalMux I__1024 (
            .O(N__10155),
            .I(\uu2.r_data_wire_5 ));
    InMux I__1023 (
            .O(N__10152),
            .I(N__10149));
    LocalMux I__1022 (
            .O(N__10149),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1021 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__1020 (
            .O(N__10143),
            .I(\uu2.r_data_wire_7 ));
    InMux I__1019 (
            .O(N__10140),
            .I(N__10137));
    LocalMux I__1018 (
            .O(N__10137),
            .I(vbuf_tx_data_0));
    InMux I__1017 (
            .O(N__10134),
            .I(N__10131));
    LocalMux I__1016 (
            .O(N__10131),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1015 (
            .O(N__10128),
            .I(N__10125));
    LocalMux I__1014 (
            .O(N__10125),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1013 (
            .O(N__10122),
            .I(N__10119));
    LocalMux I__1012 (
            .O(N__10119),
            .I(N__10116));
    Span12Mux_s1_h I__1011 (
            .O(N__10116),
            .I(N__10113));
    Odrv12 I__1010 (
            .O(N__10113),
            .I(o_serial_data_c));
    InMux I__1009 (
            .O(N__10110),
            .I(N__10105));
    InMux I__1008 (
            .O(N__10109),
            .I(N__10100));
    InMux I__1007 (
            .O(N__10108),
            .I(N__10100));
    LocalMux I__1006 (
            .O(N__10105),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1005 (
            .O(N__10100),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__1004 (
            .O(N__10095),
            .I(N__10092));
    InMux I__1003 (
            .O(N__10092),
            .I(N__10086));
    InMux I__1002 (
            .O(N__10091),
            .I(N__10079));
    InMux I__1001 (
            .O(N__10090),
            .I(N__10079));
    InMux I__1000 (
            .O(N__10089),
            .I(N__10079));
    LocalMux I__999 (
            .O(N__10086),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__998 (
            .O(N__10079),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__997 (
            .O(N__10074),
            .I(N__10069));
    InMux I__996 (
            .O(N__10073),
            .I(N__10064));
    InMux I__995 (
            .O(N__10072),
            .I(N__10064));
    LocalMux I__994 (
            .O(N__10069),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__993 (
            .O(N__10064),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__992 (
            .O(N__10059),
            .I(N__10056));
    InMux I__991 (
            .O(N__10056),
            .I(N__10053));
    LocalMux I__990 (
            .O(N__10053),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__989 (
            .O(N__10050),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__988 (
            .O(N__10047),
            .I(N__10043));
    InMux I__987 (
            .O(N__10046),
            .I(N__10040));
    LocalMux I__986 (
            .O(N__10043),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__985 (
            .O(N__10040),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__984 (
            .O(N__10035),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    CascadeMux I__983 (
            .O(N__10032),
            .I(N__10028));
    CascadeMux I__982 (
            .O(N__10031),
            .I(N__10024));
    InMux I__981 (
            .O(N__10028),
            .I(N__10021));
    InMux I__980 (
            .O(N__10027),
            .I(N__10018));
    InMux I__979 (
            .O(N__10024),
            .I(N__10015));
    LocalMux I__978 (
            .O(N__10021),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__977 (
            .O(N__10018),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__976 (
            .O(N__10015),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__975 (
            .O(N__10008),
            .I(N__10005));
    LocalMux I__974 (
            .O(N__10005),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__973 (
            .O(N__10002),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__972 (
            .O(N__9999),
            .I(N__9990));
    InMux I__971 (
            .O(N__9998),
            .I(N__9990));
    InMux I__970 (
            .O(N__9997),
            .I(N__9985));
    InMux I__969 (
            .O(N__9996),
            .I(N__9985));
    InMux I__968 (
            .O(N__9995),
            .I(N__9982));
    LocalMux I__967 (
            .O(N__9990),
            .I(N__9979));
    LocalMux I__966 (
            .O(N__9985),
            .I(buart__rx_ser_clk));
    LocalMux I__965 (
            .O(N__9982),
            .I(buart__rx_ser_clk));
    Odrv4 I__964 (
            .O(N__9979),
            .I(buart__rx_ser_clk));
    InMux I__963 (
            .O(N__9972),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__962 (
            .O(N__9969),
            .I(N__9966));
    InMux I__961 (
            .O(N__9966),
            .I(N__9962));
    InMux I__960 (
            .O(N__9965),
            .I(N__9959));
    LocalMux I__959 (
            .O(N__9962),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__958 (
            .O(N__9959),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__957 (
            .O(N__9954),
            .I(N__9951));
    LocalMux I__956 (
            .O(N__9951),
            .I(\uu2.r_data_wire_0 ));
    InMux I__955 (
            .O(N__9948),
            .I(N__9945));
    LocalMux I__954 (
            .O(N__9945),
            .I(\uu2.r_data_wire_1 ));
    InMux I__953 (
            .O(N__9942),
            .I(N__9939));
    LocalMux I__952 (
            .O(N__9939),
            .I(uart_RXD));
    CascadeMux I__951 (
            .O(N__9936),
            .I(N__9932));
    InMux I__950 (
            .O(N__9935),
            .I(N__9927));
    InMux I__949 (
            .O(N__9932),
            .I(N__9927));
    LocalMux I__948 (
            .O(N__9927),
            .I(\Lab_UT.dispString.N_115_mux ));
    CascadeMux I__947 (
            .O(N__9924),
            .I(\Lab_UT.dispString.N_115_mux_cascade_ ));
    InMux I__946 (
            .O(N__9921),
            .I(N__9914));
    InMux I__945 (
            .O(N__9920),
            .I(N__9911));
    InMux I__944 (
            .O(N__9919),
            .I(N__9904));
    InMux I__943 (
            .O(N__9918),
            .I(N__9904));
    InMux I__942 (
            .O(N__9917),
            .I(N__9904));
    LocalMux I__941 (
            .O(N__9914),
            .I(buart__rx_bitcount_1));
    LocalMux I__940 (
            .O(N__9911),
            .I(buart__rx_bitcount_1));
    LocalMux I__939 (
            .O(N__9904),
            .I(buart__rx_bitcount_1));
    CascadeMux I__938 (
            .O(N__9897),
            .I(N__9892));
    CascadeMux I__937 (
            .O(N__9896),
            .I(N__9888));
    CascadeMux I__936 (
            .O(N__9895),
            .I(N__9885));
    InMux I__935 (
            .O(N__9892),
            .I(N__9878));
    InMux I__934 (
            .O(N__9891),
            .I(N__9878));
    InMux I__933 (
            .O(N__9888),
            .I(N__9878));
    InMux I__932 (
            .O(N__9885),
            .I(N__9875));
    LocalMux I__931 (
            .O(N__9878),
            .I(N__9872));
    LocalMux I__930 (
            .O(N__9875),
            .I(buart__rx_bitcount_4));
    Odrv4 I__929 (
            .O(N__9872),
            .I(buart__rx_bitcount_4));
    CascadeMux I__928 (
            .O(N__9867),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    InMux I__927 (
            .O(N__9864),
            .I(N__9861));
    LocalMux I__926 (
            .O(N__9861),
            .I(\Lab_UT.dispString.N_177 ));
    CascadeMux I__925 (
            .O(N__9858),
            .I(buart__rx_ser_clk_cascade_));
    InMux I__924 (
            .O(N__9855),
            .I(N__9851));
    InMux I__923 (
            .O(N__9854),
            .I(N__9845));
    LocalMux I__922 (
            .O(N__9851),
            .I(N__9842));
    InMux I__921 (
            .O(N__9850),
            .I(N__9839));
    InMux I__920 (
            .O(N__9849),
            .I(N__9834));
    InMux I__919 (
            .O(N__9848),
            .I(N__9834));
    LocalMux I__918 (
            .O(N__9845),
            .I(buart__rx_bitcount_0));
    Odrv4 I__917 (
            .O(N__9842),
            .I(buart__rx_bitcount_0));
    LocalMux I__916 (
            .O(N__9839),
            .I(buart__rx_bitcount_0));
    LocalMux I__915 (
            .O(N__9834),
            .I(buart__rx_bitcount_0));
    IoInMux I__914 (
            .O(N__9825),
            .I(N__9822));
    LocalMux I__913 (
            .O(N__9822),
            .I(N__9819));
    IoSpan4Mux I__912 (
            .O(N__9819),
            .I(N__9816));
    Span4Mux_s0_v I__911 (
            .O(N__9816),
            .I(N__9813));
    Span4Mux_v I__910 (
            .O(N__9813),
            .I(N__9810));
    Odrv4 I__909 (
            .O(N__9810),
            .I(buart__rx_sample));
    CascadeMux I__908 (
            .O(N__9807),
            .I(N__9804));
    InMux I__907 (
            .O(N__9804),
            .I(N__9801));
    LocalMux I__906 (
            .O(N__9801),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    InMux I__905 (
            .O(N__9798),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__904 (
            .O(N__9795),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__903 (
            .O(N__9792),
            .I(Lab_UT_dispString_m103_ns_1_cascade_));
    InMux I__902 (
            .O(N__9789),
            .I(N__9786));
    LocalMux I__901 (
            .O(N__9786),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    CascadeMux I__900 (
            .O(N__9783),
            .I(buart__rx_N_27_0_i_cascade_));
    InMux I__899 (
            .O(N__9780),
            .I(N__9777));
    LocalMux I__898 (
            .O(N__9777),
            .I(N__9774));
    Odrv4 I__897 (
            .O(N__9774),
            .I(N_179));
    InMux I__896 (
            .O(N__9771),
            .I(N__9765));
    InMux I__895 (
            .O(N__9770),
            .I(N__9758));
    InMux I__894 (
            .O(N__9769),
            .I(N__9758));
    InMux I__893 (
            .O(N__9768),
            .I(N__9758));
    LocalMux I__892 (
            .O(N__9765),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__891 (
            .O(N__9758),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__890 (
            .O(N__9753),
            .I(resetGen_reset_count_2_2_cascade_));
    CascadeMux I__889 (
            .O(N__9750),
            .I(N__9744));
    InMux I__888 (
            .O(N__9749),
            .I(N__9735));
    InMux I__887 (
            .O(N__9748),
            .I(N__9735));
    InMux I__886 (
            .O(N__9747),
            .I(N__9735));
    InMux I__885 (
            .O(N__9744),
            .I(N__9735));
    LocalMux I__884 (
            .O(N__9735),
            .I(resetGen_reset_count_2));
    InMux I__883 (
            .O(N__9732),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__882 (
            .O(N__9729),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__881 (
            .O(N__9726),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__880 (
            .O(N__9723),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__879 (
            .O(N__9720),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__878 (
            .O(N__9717),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__877 (
            .O(N__9714),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    InMux I__876 (
            .O(N__9711),
            .I(N__9705));
    InMux I__875 (
            .O(N__9710),
            .I(N__9705));
    LocalMux I__874 (
            .O(N__9705),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    InMux I__873 (
            .O(N__9702),
            .I(N__9696));
    InMux I__872 (
            .O(N__9701),
            .I(N__9696));
    LocalMux I__871 (
            .O(N__9696),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__870 (
            .O(N__9693),
            .I(N__9689));
    CascadeMux I__869 (
            .O(N__9692),
            .I(N__9686));
    InMux I__868 (
            .O(N__9689),
            .I(N__9681));
    InMux I__867 (
            .O(N__9686),
            .I(N__9681));
    LocalMux I__866 (
            .O(N__9681),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__865 (
            .O(N__9678),
            .I(N__9672));
    InMux I__864 (
            .O(N__9677),
            .I(N__9672));
    LocalMux I__863 (
            .O(N__9672),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__862 (
            .O(N__9669),
            .I(N__9665));
    InMux I__861 (
            .O(N__9668),
            .I(N__9662));
    InMux I__860 (
            .O(N__9665),
            .I(N__9659));
    LocalMux I__859 (
            .O(N__9662),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__858 (
            .O(N__9659),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__857 (
            .O(N__9654),
            .I(N__9651));
    LocalMux I__856 (
            .O(N__9651),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__855 (
            .O(N__9648),
            .I(N__9645));
    InMux I__854 (
            .O(N__9645),
            .I(N__9640));
    InMux I__853 (
            .O(N__9644),
            .I(N__9635));
    InMux I__852 (
            .O(N__9643),
            .I(N__9635));
    LocalMux I__851 (
            .O(N__9640),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__850 (
            .O(N__9635),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__849 (
            .O(N__9630),
            .I(N__9627));
    InMux I__848 (
            .O(N__9627),
            .I(N__9615));
    InMux I__847 (
            .O(N__9626),
            .I(N__9615));
    InMux I__846 (
            .O(N__9625),
            .I(N__9615));
    InMux I__845 (
            .O(N__9624),
            .I(N__9610));
    InMux I__844 (
            .O(N__9623),
            .I(N__9610));
    InMux I__843 (
            .O(N__9622),
            .I(N__9607));
    LocalMux I__842 (
            .O(N__9615),
            .I(N__9602));
    LocalMux I__841 (
            .O(N__9610),
            .I(N__9602));
    LocalMux I__840 (
            .O(N__9607),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__839 (
            .O(N__9602),
            .I(\uu0.l_precountZ0Z_0 ));
    CascadeMux I__838 (
            .O(N__9597),
            .I(\uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__837 (
            .O(N__9594),
            .I(\uu0.un154_ci_9_cascade_ ));
    CascadeMux I__836 (
            .O(N__9591),
            .I(\uu0.un187_ci_1_cascade_ ));
    InMux I__835 (
            .O(N__9588),
            .I(N__9576));
    InMux I__834 (
            .O(N__9587),
            .I(N__9576));
    InMux I__833 (
            .O(N__9586),
            .I(N__9576));
    InMux I__832 (
            .O(N__9585),
            .I(N__9576));
    LocalMux I__831 (
            .O(N__9576),
            .I(\uu0.l_countZ0Z_14 ));
    CascadeMux I__830 (
            .O(N__9573),
            .I(N__9568));
    InMux I__829 (
            .O(N__9572),
            .I(N__9561));
    InMux I__828 (
            .O(N__9571),
            .I(N__9561));
    InMux I__827 (
            .O(N__9568),
            .I(N__9561));
    LocalMux I__826 (
            .O(N__9561),
            .I(\uu0.l_countZ0Z_15 ));
    CascadeMux I__825 (
            .O(N__9558),
            .I(N__9553));
    CascadeMux I__824 (
            .O(N__9557),
            .I(N__9550));
    InMux I__823 (
            .O(N__9556),
            .I(N__9543));
    InMux I__822 (
            .O(N__9553),
            .I(N__9543));
    InMux I__821 (
            .O(N__9550),
            .I(N__9543));
    LocalMux I__820 (
            .O(N__9543),
            .I(\uu0.l_precountZ0Z_3 ));
    InMux I__819 (
            .O(N__9540),
            .I(N__9525));
    InMux I__818 (
            .O(N__9539),
            .I(N__9525));
    InMux I__817 (
            .O(N__9538),
            .I(N__9525));
    InMux I__816 (
            .O(N__9537),
            .I(N__9525));
    InMux I__815 (
            .O(N__9536),
            .I(N__9525));
    LocalMux I__814 (
            .O(N__9525),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__813 (
            .O(N__9522),
            .I(N__9516));
    InMux I__812 (
            .O(N__9521),
            .I(N__9507));
    InMux I__811 (
            .O(N__9520),
            .I(N__9507));
    InMux I__810 (
            .O(N__9519),
            .I(N__9507));
    InMux I__809 (
            .O(N__9516),
            .I(N__9507));
    LocalMux I__808 (
            .O(N__9507),
            .I(\uu0.l_precountZ0Z_2 ));
    IoInMux I__807 (
            .O(N__9504),
            .I(N__9501));
    LocalMux I__806 (
            .O(N__9501),
            .I(N__9498));
    IoSpan4Mux I__805 (
            .O(N__9498),
            .I(N__9495));
    Odrv4 I__804 (
            .O(N__9495),
            .I(clk_in_c));
    INV \INVuu2.bitmap_84C  (
            .O(\INVuu2.bitmap_84C_net ),
            .I(N__26194));
    INV \INVuu2.bitmap_212C  (
            .O(\INVuu2.bitmap_212C_net ),
            .I(N__26200));
    INV \INVuu2.w_addr_displaying_0C  (
            .O(\INVuu2.w_addr_displaying_0C_net ),
            .I(N__26204));
    INV \INVuu2.bitmap_87C  (
            .O(\INVuu2.bitmap_87C_net ),
            .I(N__26186));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__26193));
    INV \INVuu2.w_addr_user_5C  (
            .O(\INVuu2.w_addr_user_5C_net ),
            .I(N__26203));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__26178));
    INV \INVuu2.bitmap_215C  (
            .O(\INVuu2.bitmap_215C_net ),
            .I(N__26185));
    INV \INVuu2.w_addr_displaying_3C  (
            .O(\INVuu2.w_addr_displaying_3C_net ),
            .I(N__26192));
    INV \INVuu2.w_addr_displaying_nesr_5C  (
            .O(\INVuu2.w_addr_displaying_nesr_5C_net ),
            .I(N__26199));
    INV \INVuu2.bitmap_197C  (
            .O(\INVuu2.bitmap_197C_net ),
            .I(N__26177));
    INV \INVuu2.w_addr_displaying_1C  (
            .O(\INVuu2.w_addr_displaying_1C_net ),
            .I(N__26184));
    INV \INVuu2.bitmap_203C  (
            .O(\INVuu2.bitmap_203C_net ),
            .I(N__26191));
    INV \INVuu2.bitmap_111C  (
            .O(\INVuu2.bitmap_111C_net ),
            .I(N__26152));
    INV \INVuu2.bitmap_66C  (
            .O(\INVuu2.bitmap_66C_net ),
            .I(N__26160));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__26169));
    INV \INVuu2.w_addr_displaying_4C  (
            .O(\INVuu2.w_addr_displaying_4C_net ),
            .I(N__26163));
    INV \INVuu2.w_addr_user_nesr_8C  (
            .O(\INVuu2.w_addr_user_nesr_8C_net ),
            .I(N__26176));
    INV \INVuu2.w_addr_user_1C  (
            .O(\INVuu2.w_addr_user_1C_net ),
            .I(N__26183));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__26202));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_13_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__11862),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB bu_rx_data_rdy_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__25611),
            .GLOBALBUFFEROUTPUT(bu_rx_data_rdy_0_g));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__11544),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    ICE_GB \buart.Z_rx.sample_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__9825),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__16693),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.vram_rd_clk_LC_1_1_0 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_1_1_0 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_1_1_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_1_1_0  (
            .in0(_gnd_net_),
            .in1(N__14667),
            .in2(_gnd_net_),
            .in3(N__11439),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(),
            .sr(N__25833));
    defparam \uu0.l_precount_0_LC_1_1_1 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_1_1_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_1_1_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_1_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9622),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26205),
            .ce(),
            .sr(N__25833));
    defparam \uu0.l_count_5_LC_1_2_0 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_1_2_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_1_2_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu0.l_count_5_LC_1_2_0  (
            .in0(N__10624),
            .in1(N__12257),
            .in2(_gnd_net_),
            .in3(N__12236),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__10442),
            .sr(N__25830));
    defparam \uu0.l_count_8_LC_1_2_1 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_2_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_count_8_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__10488),
            .in2(_gnd_net_),
            .in3(N__10328),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26201),
            .ce(N__10442),
            .sr(N__25830));
    defparam \uu0.delay_line_0_LC_1_3_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_3_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_3_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_3_0  (
            .in0(N__9537),
            .in1(N__9625),
            .in2(N__9558),
            .in3(N__9519),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26195),
            .ce(),
            .sr(N__25827));
    defparam \uu0.l_precount_3_LC_1_3_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_3_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_3_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_3_1  (
            .in0(N__9521),
            .in1(N__9556),
            .in2(N__9630),
            .in3(N__9540),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26195),
            .ce(),
            .sr(N__25827));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_3_2 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_3_2  (
            .in0(N__9536),
            .in1(N__12253),
            .in2(N__9557),
            .in3(N__10377),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_1_LC_1_3_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_3_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_3_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_precount_1_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__9624),
            .in2(_gnd_net_),
            .in3(N__9538),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26195),
            .ce(),
            .sr(N__25827));
    defparam \uu0.l_precount_2_LC_1_3_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_3_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_3_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_1_3_4  (
            .in0(N__9539),
            .in1(N__9626),
            .in2(_gnd_net_),
            .in3(N__9520),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26195),
            .ce(),
            .sr(N__25827));
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_3_5 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI3Q7K1_2_LC_1_3_5  (
            .in0(N__10317),
            .in1(N__10659),
            .in2(N__9522),
            .in3(N__10400),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIO2782_16_LC_1_3_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNIO2782_16_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIO2782_16_LC_1_3_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNIO2782_16_LC_1_3_6  (
            .in0(N__9623),
            .in1(N__10242),
            .in2(N__9597),
            .in3(N__10773),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_4_0 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_4_0  (
            .in0(N__10770),
            .in1(N__9571),
            .in2(N__10744),
            .in3(N__9586),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_4_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_4_1  (
            .in0(N__10354),
            .in1(N__10329),
            .in2(N__10566),
            .in3(N__10295),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_4_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_4_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_4_2  (
            .in0(N__10771),
            .in1(_gnd_net_),
            .in2(N__9594),
            .in3(N__9587),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_4_3 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_4_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_4_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_15_LC_1_4_3  (
            .in0(N__9572),
            .in1(N__10496),
            .in2(N__9591),
            .in3(N__11595),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26188),
            .ce(N__10439),
            .sr(N__25824));
    defparam \uu0.l_count_14_LC_1_4_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_4_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_4_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_14_LC_1_4_4  (
            .in0(N__10772),
            .in1(N__10494),
            .in2(N__10745),
            .in3(N__9588),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26188),
            .ce(N__10439),
            .sr(N__25824));
    defparam \uu0.l_count_4_LC_1_4_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_4_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_4_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu0.l_count_4_LC_1_4_5  (
            .in0(N__10623),
            .in1(N__12226),
            .in2(_gnd_net_),
            .in3(N__11596),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26188),
            .ce(N__10439),
            .sr(N__25824));
    defparam \uu0.l_count_10_LC_1_4_6 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_4_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_4_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_10_LC_1_4_6  (
            .in0(N__10296),
            .in1(N__10495),
            .in2(N__10335),
            .in3(N__10355),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26188),
            .ce(N__10439),
            .sr(N__25824));
    defparam \uu0.l_count_RNIGTCU_15_LC_1_4_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_4_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu0.l_count_RNIGTCU_15_LC_1_4_7  (
            .in0(N__9585),
            .in1(N__10353),
            .in2(N__9573),
            .in3(N__12225),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_5_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__9771),
            .in2(N__9648),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_5_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_5_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_1_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_1_5_1  (
            .in0(_gnd_net_),
            .in1(N__9678),
            .in2(_gnd_net_),
            .in3(N__9726),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__26180),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_5_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_5_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_1_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_1_5_2  (
            .in0(N__11488),
            .in1(N__9668),
            .in2(_gnd_net_),
            .in3(N__9723),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__26180),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_5_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_1_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(N__9702),
            .in2(_gnd_net_),
            .in3(N__9720),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__26180),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_5_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_1_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_1_5_4  (
            .in0(N__11489),
            .in1(N__9711),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__26180),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_5_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_5_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_1_5_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__11487),
            .in2(N__9693),
            .in3(N__9714),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26180),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_1_5_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_1_5_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_1_5_7  (
            .in0(N__9710),
            .in1(N__9701),
            .in2(N__9692),
            .in3(N__9677),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_0  (
            .in0(N__9643),
            .in1(N__9768),
            .in2(N__9669),
            .in3(N__9654),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_6_4 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_6_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_1_6_4  (
            .in0(N__9644),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9770),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26173),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_6_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_1_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9769),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26173),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m75_LC_1_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m75_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m75_LC_1_7_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.m75_LC_1_7_2  (
            .in0(N__10689),
            .in1(N__10868),
            .in2(N__9750),
            .in3(N__12608),
            .lcout(N_105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m82_LC_1_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m82_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m82_LC_1_7_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.dictrl.m82_LC_1_7_3  (
            .in0(N__12610),
            .in1(N__10691),
            .in2(N__10880),
            .in3(N__9747),
            .lcout(),
            .ltout(resetGen_reset_count_2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_1_7_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_1_7_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_1_7_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \resetGen.reset_count_2_LC_1_7_4  (
            .in0(N__9749),
            .in1(N__10909),
            .in2(N__9753),
            .in3(N__12611),
            .lcout(resetGen_reset_count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26165),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m78_LC_1_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m78_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m78_LC_1_7_5 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Lab_UT.dictrl.m78_LC_1_7_5  (
            .in0(N__12609),
            .in1(N__10690),
            .in2(N__10879),
            .in3(N__9748),
            .lcout(N_107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_1_7_6 .C_ON=1'b0;
    defparam \resetGen.rst_LC_1_7_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_1_7_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10910),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26165),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_1_8_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_8_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_8_7 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_1_8_7  (
            .in0(N__16250),
            .in1(N__16181),
            .in2(N__9807),
            .in3(N__14951),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26156),
            .ce(N__16081),
            .sr(N__25817));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_9_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__9850),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_9_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(N__9920),
            .in2(_gnd_net_),
            .in3(N__9732),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_9_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__16131),
            .in2(_gnd_net_),
            .in3(N__9729),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_9_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__14950),
            .in2(_gnd_net_),
            .in3(N__9798),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_1_9_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_9_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_9_4 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_1_9_4  (
            .in0(N__16249),
            .in1(N__16174),
            .in2(N__9895),
            .in3(N__9795),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26150),
            .ce(N__16085),
            .sr(N__25818));
    defparam \Lab_UT.dispString.m103_ns_1_LC_1_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m103_ns_1_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m103_ns_1_LC_1_10_0 .LUT_INIT=16'b0010111000111111;
    LogicCell40 \Lab_UT.dispString.m103_ns_1_LC_1_10_0  (
            .in0(N__9998),
            .in1(N__14958),
            .in2(N__9936),
            .in3(N__14882),
            .lcout(),
            .ltout(Lab_UT_dispString_m103_ns_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_1_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_1_10_1 .LUT_INIT=16'b1101101111001010;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_1_10_1  (
            .in0(N__9780),
            .in1(N__9999),
            .in2(N__9792),
            .in3(N__25924),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_1_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_1_10_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_1_10_4 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_1_10_4  (
            .in0(N__16238),
            .in1(N__16173),
            .in2(N__16959),
            .in3(N__9854),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26144),
            .ce(N__16077),
            .sr(N__25819));
    defparam \Lab_UT.dispString.N_27_0_i_LC_1_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.N_27_0_i_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.N_27_0_i_LC_1_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.dispString.N_27_0_i_LC_1_10_5  (
            .in0(N__14883),
            .in1(N__9935),
            .in2(_gnd_net_),
            .in3(N__14959),
            .lcout(buart__rx_N_27_0_i),
            .ltout(buart__rx_N_27_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_1_LC_1_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_10_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_10_6 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_1_10_6  (
            .in0(N__16239),
            .in1(N__9789),
            .in2(N__9783),
            .in3(N__9921),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26144),
            .ce(N__16077),
            .sr(N__25819));
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_1_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_1_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_1_11_0  (
            .in0(N__16128),
            .in1(N__9917),
            .in2(N__9896),
            .in3(N__9848),
            .lcout(buart__rx_valid_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m103_e_LC_1_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m103_e_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m103_e_LC_1_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dispString.m103_e_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__11740),
            .in2(_gnd_net_),
            .in3(N__10846),
            .lcout(N_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_1_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_11_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9942),
            .lcout(buart__rx_hh_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26135),
            .ce(),
            .sr(N__25821));
    defparam \Lab_UT.dispString.m8_LC_1_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m8_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m8_LC_1_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dispString.m8_LC_1_11_4  (
            .in0(N__16129),
            .in1(N__9919),
            .in2(N__9897),
            .in3(N__9849),
            .lcout(\Lab_UT.dispString.N_115_mux ),
            .ltout(\Lab_UT.dispString.N_115_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m11_LC_1_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m11_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m11_LC_1_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dispString.m11_LC_1_11_5  (
            .in0(N__14960),
            .in1(N__10847),
            .in2(N__9924),
            .in3(N__11741),
            .lcout(buart__rx_startbit),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m97_e_LC_1_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m97_e_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m97_e_LC_1_11_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dispString.m97_e_LC_1_11_7  (
            .in0(N__9918),
            .in1(N__9891),
            .in2(_gnd_net_),
            .in3(N__14957),
            .lcout(\Lab_UT.dispString.N_177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_1_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_1_12_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_1_12_0  (
            .in0(N__10073),
            .in1(N__16241),
            .in2(N__10059),
            .in3(N__9996),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26131),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_12_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_12_1  (
            .in0(N__10046),
            .in1(N__10072),
            .in2(N__10031),
            .in3(N__10108),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_12_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_12_2  (
            .in0(_gnd_net_),
            .in1(N__9965),
            .in2(N__9867),
            .in3(N__10089),
            .lcout(buart__rx_ser_clk),
            .ltout(buart__rx_ser_clk_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m98_LC_1_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m98_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m98_LC_1_12_3 .LUT_INIT=16'b1101000000000000;
    LogicCell40 \Lab_UT.dispString.m98_LC_1_12_3  (
            .in0(N__9864),
            .in1(N__16130),
            .in2(N__9858),
            .in3(N__9855),
            .lcout(buart__rx_sample),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_12_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_1_12_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_1_12_4  (
            .in0(N__10008),
            .in1(N__16242),
            .in2(N__10032),
            .in3(N__9997),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26131),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_12_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_1_12_5 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_1_12_5  (
            .in0(N__10091),
            .in1(_gnd_net_),
            .in2(N__16253),
            .in3(N__10109),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26131),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_1_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_1_12_6  (
            .in0(_gnd_net_),
            .in1(N__16240),
            .in2(_gnd_net_),
            .in3(N__10090),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26131),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_13_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__10110),
            .in2(N__10095),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_13_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_13_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(N__10074),
            .in2(_gnd_net_),
            .in3(N__10050),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_13_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_1_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_1_13_2  (
            .in0(N__16252),
            .in1(N__10047),
            .in2(_gnd_net_),
            .in3(N__10035),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__26128),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_13_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_13_3  (
            .in0(_gnd_net_),
            .in1(N__10027),
            .in2(_gnd_net_),
            .in3(N__10002),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_1_13_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_1_13_4  (
            .in0(N__9995),
            .in1(N__16251),
            .in2(N__9969),
            .in3(N__9972),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26128),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_0_LC_2_1_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_0_LC_2_1_0  (
            .in0(N__9954),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_1_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_1_LC_2_1_1  (
            .in0(N__9948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_1_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_2_LC_2_1_2  (
            .in0(N__10176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_1_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_3_LC_2_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10170),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_1_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10164),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_1_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10158),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_1_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10152),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_1_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_7_LC_2_1_7  (
            .in0(N__10146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__16011),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_2_0  (
            .in0(N__12122),
            .in1(N__10221),
            .in2(_gnd_net_),
            .in3(N__10140),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__10134),
            .in2(_gnd_net_),
            .in3(N__12120),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_2_2  (
            .in0(N__12121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10128),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_2_3  (
            .in0(N__10209),
            .in1(N__12123),
            .in2(_gnd_net_),
            .in3(N__10227),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_2_4  (
            .in0(N__12124),
            .in1(N__10197),
            .in2(_gnd_net_),
            .in3(N__10215),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_2_5  (
            .in0(N__10185),
            .in1(N__12125),
            .in2(_gnd_net_),
            .in3(N__10203),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_2_6  (
            .in0(N__12126),
            .in1(N__10413),
            .in2(_gnd_net_),
            .in3(N__10191),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26196),
            .ce(N__10803),
            .sr(N__25834));
    defparam \uu0.l_count_6_LC_2_3_0 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_2_3_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_2_3_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_6_LC_2_3_0  (
            .in0(N__12372),
            .in1(N__12346),
            .in2(N__10625),
            .in3(N__11601),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26189),
            .ce(N__10443),
            .sr(N__25832));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_3_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_3_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_3_1  (
            .in0(N__10381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10402),
            .lcout(\uu0.un44_ci ),
            .ltout(\uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_2_3_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_2_3_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_2_3_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu0.l_count_2_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10179),
            .in3(N__10661),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26189),
            .ce(N__10443),
            .sr(N__25832));
    defparam \uu0.l_count_1_LC_2_3_3 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_2_3_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_2_3_3  (
            .in0(N__10382),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10404),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26189),
            .ce(N__10443),
            .sr(N__25832));
    defparam \uu0.l_count_0_LC_2_3_4 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_2_3_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_2_3_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_2_3_4  (
            .in0(N__10403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11599),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26189),
            .ce(N__10443),
            .sr(N__25832));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_3_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_3_5  (
            .in0(N__10660),
            .in1(N__10401),
            .in2(N__10383),
            .in3(N__10641),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_3_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_3_6  (
            .in0(N__12371),
            .in1(N__12345),
            .in2(N__10362),
            .in3(N__10596),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_12_LC_2_3_7 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_2_3_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_2_3_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_12_LC_2_3_7  (
            .in0(N__11600),
            .in1(N__10743),
            .in2(N__10359),
            .in3(N__10714),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26189),
            .ce(N__10443),
            .sr(N__25832));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_4_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_4_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_4_0  (
            .in0(N__10292),
            .in1(N__10594),
            .in2(N__10275),
            .in3(N__10639),
            .lcout(\uu0.un4_l_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_4_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_4_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_4_1  (
            .in0(N__10333),
            .in1(N__10356),
            .in2(_gnd_net_),
            .in3(N__10293),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_9_LC_2_4_2 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_2_4_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_2_4_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu0.l_count_9_LC_2_4_2  (
            .in0(N__10294),
            .in1(N__10487),
            .in2(_gnd_net_),
            .in3(N__10334),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26181),
            .ce(N__10441),
            .sr(N__25828));
    defparam \uu0.l_count_17_LC_2_4_3 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_4_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_17_LC_2_4_3  (
            .in0(N__10245),
            .in1(N__10259),
            .in2(N__10498),
            .in3(N__10274),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26181),
            .ce(N__10441),
            .sr(N__25828));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_4_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_4_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_4_4  (
            .in0(N__10273),
            .in1(N__10480),
            .in2(N__10260),
            .in3(N__10243),
            .lcout(\uu0.un220_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_2_4_5 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_2_4_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_2_4_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_16_LC_2_4_5  (
            .in0(N__10244),
            .in1(N__10258),
            .in2(N__10497),
            .in3(N__11585),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26181),
            .ce(N__10441),
            .sr(N__25828));
    defparam \uu0.l_count_3_LC_2_4_6 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_2_4_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_3_LC_2_4_6  (
            .in0(N__11587),
            .in1(N__10674),
            .in2(N__10668),
            .in3(N__10640),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26181),
            .ce(N__10441),
            .sr(N__25828));
    defparam \uu0.l_count_7_LC_2_4_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_2_4_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_7_LC_2_4_7  (
            .in0(N__10595),
            .in1(N__12324),
            .in2(N__10626),
            .in3(N__11586),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26181),
            .ce(N__10441),
            .sr(N__25828));
    defparam \uu0.l_count_18_LC_2_5_0 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_5_0 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \uu0.l_count_18_LC_2_5_0  (
            .in0(N__11584),
            .in1(_gnd_net_),
            .in2(N__10548),
            .in3(N__10581),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26174),
            .ce(N__10440),
            .sr(N__25825));
    defparam \uu0.l_count_11_LC_2_5_1 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_2_5_1 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_11_LC_2_5_1  (
            .in0(N__10499),
            .in1(N__10562),
            .in2(N__10575),
            .in3(N__11583),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26174),
            .ce(N__10440),
            .sr(N__25825));
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_5_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIOIDD2_18_LC_2_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNIOIDD2_18_LC_2_5_2  (
            .in0(N__10561),
            .in1(N__12350),
            .in2(N__10547),
            .in3(N__10533),
            .lcout(),
            .ltout(\uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_5_3 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_15_LC_2_5_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_15_LC_2_5_3  (
            .in0(N__10527),
            .in1(N__10518),
            .in2(N__10512),
            .in3(N__10509),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_13_LC_2_5_4 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_2_5_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uu0.l_count_13_LC_2_5_4  (
            .in0(N__10698),
            .in1(N__10500),
            .in2(N__10446),
            .in3(N__10785),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26174),
            .ce(N__10440),
            .sr(N__25825));
    defparam \buart.Z_tx.shifter_6_LC_2_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_6_0  (
            .in0(N__12117),
            .in1(N__10824),
            .in2(_gnd_net_),
            .in3(N__10422),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26166),
            .ce(N__10796),
            .sr(N__25823));
    defparam \buart.Z_tx.shifter_7_LC_2_6_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_6_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_6_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_6_1  (
            .in0(N__10833),
            .in1(N__10809),
            .in2(_gnd_net_),
            .in3(N__12118),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26166),
            .ce(N__10796),
            .sr(N__25823));
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_6_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_6_2  (
            .in0(N__12116),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10818),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26166),
            .ce(N__10796),
            .sr(N__25823));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__12115),
            .in2(_gnd_net_),
            .in3(N__11646),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_6_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_6_4  (
            .in0(_gnd_net_),
            .in1(N__25876),
            .in2(_gnd_net_),
            .in3(N__16635),
            .lcout(\Lab_UT.didp.regrce2.LdAStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_2_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_2_6_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_2_6_5  (
            .in0(N__25877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16665),
            .lcout(\Lab_UT.didp.regrce4.LdAMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_6_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_2_6_6  (
            .in0(N__10715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10784),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_6_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__10749),
            .in2(_gnd_net_),
            .in3(N__10716),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_2_7_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_2_7_1 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_2_7_1  (
            .in0(N__12614),
            .in1(N__10905),
            .in2(N__10881),
            .in3(N__10692),
            .lcout(resetGen_reset_count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26157),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m72_LC_2_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m72_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m72_LC_2_7_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.m72_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(N__10903),
            .in2(_gnd_net_),
            .in3(N__12612),
            .lcout(),
            .ltout(m72_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_2_7_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_2_7_3 .LUT_INIT=16'b1010110110101000;
    LogicCell40 \resetGen.reset_count_3_LC_2_7_3  (
            .in0(N__10919),
            .in1(N__10938),
            .in2(N__10932),
            .in3(N__10928),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26157),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_2_7_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_2_7_4 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \resetGen.reset_count_4_LC_2_7_4  (
            .in0(N__10929),
            .in1(N__10920),
            .in2(N__10911),
            .in3(N__12615),
            .lcout(resetGen_reset_count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26157),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_2_7_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_2_7_6 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_2_7_6  (
            .in0(N__10904),
            .in1(N__10875),
            .in2(_gnd_net_),
            .in3(N__12613),
            .lcout(resetGen_reset_count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26157),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_1_LC_2_9_2 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_2_9_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_2_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10851),
            .lcout(buart__rx_hh_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26145),
            .ce(),
            .sr(N__25820));
    defparam \buart.Z_rx.shifter_2_rep2_LC_2_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep2_LC_2_10_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep2_LC_2_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep2_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26389),
            .lcout(bu_rx_data_2_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_3_rep1_LC_2_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_2_10_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_2_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18875),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_4_LC_2_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_2_10_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_2_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19047),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_3_rep2_LC_2_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_LC_2_10_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep2_LC_2_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18876),
            .lcout(bu_rx_data_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_5_rep1_LC_2_10_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_rep1_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_rep1_LC_2_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_rep1_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19212),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_7_rep1_LC_2_10_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_2_10_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_2_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_2_10_5  (
            .in0(N__11736),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_7_LC_2_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_2_10_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_2_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11735),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \buart.Z_rx.shifter_1_rep2_LC_2_10_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep2_LC_2_10_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep2_LC_2_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_rep2_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26651),
            .lcout(bu_rx_data_1_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26136),
            .ce(N__14244),
            .sr(N__25822));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIEGPT_LC_2_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIEGPT_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIEGPT_LC_2_11_0 .LUT_INIT=16'b0100000001110011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIEGPT_LC_2_11_0  (
            .in0(N__18586),
            .in1(N__18339),
            .in2(N__20503),
            .in3(N__19729),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_69_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIDS133_LC_2_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIDS133_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIDS133_LC_2_11_1 .LUT_INIT=16'b1000010100000101;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIDS133_LC_2_11_1  (
            .in0(N__18340),
            .in1(N__10959),
            .in2(N__10962),
            .in3(N__14370),
            .lcout(\Lab_UT.dictrl.N_61_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_1_LC_2_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_1_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_1_LC_2_11_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_1_LC_2_11_2  (
            .in0(N__13927),
            .in1(N__13839),
            .in2(N__18724),
            .in3(N__17117),
            .lcout(\Lab_UT.dictrl.g1_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_10_LC_2_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_10_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_10_LC_2_11_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \Lab_UT.dictrl.g1_10_LC_2_11_3  (
            .in0(N__13838),
            .in1(N__20489),
            .in2(N__18725),
            .in3(N__13926),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_9_LC_2_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_9_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_9_LC_2_11_4 .LUT_INIT=16'b1111001111111111;
    LogicCell40 \Lab_UT.dictrl.g1_9_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__19191),
            .in2(N__10953),
            .in3(N__19036),
            .lcout(\Lab_UT.dictrl.g1_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNII0HP5_2_LC_2_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNII0HP5_2_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNII0HP5_2_LC_2_12_0 .LUT_INIT=16'b1101110111011000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNII0HP5_2_LC_2_12_0  (
            .in0(N__22813),
            .in1(N__10950),
            .in2(N__11061),
            .in3(N__10944),
            .lcout(\Lab_UT.dictrl.N_62_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_5_LC_2_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_5_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_5_LC_2_12_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_5_LC_2_12_1  (
            .in0(N__24317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22814),
            .lcout(\Lab_UT.dictrl.g2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_3_LC_2_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_3_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_3_LC_2_12_2 .LUT_INIT=16'b0100111100001011;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_3_LC_2_12_2  (
            .in0(N__22816),
            .in1(N__24318),
            .in2(N__12543),
            .in3(N__11886),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1792_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_2_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_2_12_3 .LUT_INIT=16'b1111100101100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_2_12_3  (
            .in0(N__24319),
            .in1(N__22817),
            .in2(N__10998),
            .in3(N__10995),
            .lcout(\Lab_UT.dictrl.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIE5JQ_2_LC_2_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIE5JQ_2_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIE5JQ_2_LC_2_12_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIE5JQ_2_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__22812),
            .in2(_gnd_net_),
            .in3(N__24316),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_2_LC_2_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_2_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_2_LC_2_12_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_2_LC_2_12_5  (
            .in0(N__10971),
            .in1(N__22815),
            .in2(N__10980),
            .in3(N__11760),
            .lcout(\Lab_UT.dictrl.N_1451_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_2_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_2_13_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_2_13_0  (
            .in0(N__26616),
            .in1(N__24062),
            .in2(N__19737),
            .in3(N__21710),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_a5_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_2_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_2_13_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__10986),
            .in2(N__10989),
            .in3(N__14373),
            .lcout(\Lab_UT.dictrl.N_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_2_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_2_13_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_2_13_2  (
            .in0(N__26359),
            .in1(N__18854),
            .in2(N__25439),
            .in3(N__19209),
            .lcout(\Lab_UT.dictrl.g0_i_a5_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_8_LC_2_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_8_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_8_LC_2_13_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_8_LC_2_13_3  (
            .in0(N__21709),
            .in1(N__26358),
            .in2(N__18892),
            .in3(N__26615),
            .lcout(\Lab_UT.dictrl.g0_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_9_LC_2_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_9_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_9_LC_2_13_4 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_9_LC_2_13_4  (
            .in0(N__14372),
            .in1(N__19208),
            .in2(N__25440),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.g0_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_2_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_2_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_2_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25408),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26124),
            .ce(N__14242),
            .sr(N__25831));
    defparam \buart.Z_rx.shifter_1_LC_2_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_2_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_2_13_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_LC_2_13_6  (
            .in0(N__26617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26124),
            .ce(N__14242),
            .sr(N__25831));
    defparam \buart.Z_rx.shifter_2_LC_2_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_2_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_2_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_2_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26360),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26124),
            .ce(N__14242),
            .sr(N__25831));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI1TO01_LC_2_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI1TO01_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI1TO01_LC_2_14_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNI1TO01_LC_2_14_3  (
            .in0(N__18853),
            .in1(N__18234),
            .in2(N__18152),
            .in3(N__19730),
            .lcout(\Lab_UT.dictrl.g1_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_rep2_LC_2_15_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep2_LC_2_15_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep2_LC_2_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep2_LC_2_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18129),
            .lcout(bu_rx_data_6_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26119),
            .ce(N__14239),
            .sr(N__25837));
    defparam \uu2.r_addr_esr_7_LC_4_1_0 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_1_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_1_0  (
            .in0(N__11215),
            .in1(N__11049),
            .in2(N__11024),
            .in3(N__11977),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26190),
            .ce(N__11118),
            .sr(N__25812));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1  (
            .in0(N__11928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12005),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_1_2  (
            .in0(N__11036),
            .in1(N__11004),
            .in2(N__11043),
            .in3(N__11976),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26190),
            .ce(N__11118),
            .sr(N__25812));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_3 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_3  (
            .in0(_gnd_net_),
            .in1(N__11017),
            .in2(_gnd_net_),
            .in3(N__11214),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4  (
            .in0(N__11166),
            .in1(N__11138),
            .in2(N__11197),
            .in3(N__11098),
            .lcout(\uu2.un404_ci_0 ),
            .ltout(\uu2.un404_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_1_5  (
            .in0(N__11929),
            .in1(N__11216),
            .in2(N__11223),
            .in3(N__12006),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26190),
            .ce(N__11118),
            .sr(N__25812));
    defparam \uu2.r_addr_esr_3_LC_4_1_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_1_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_1_6  (
            .in0(N__11167),
            .in1(N__11139),
            .in2(N__11198),
            .in3(N__11099),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26190),
            .ce(N__11118),
            .sr(N__25812));
    defparam \uu2.r_addr_2_LC_4_2_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_4_2_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_4_2_0  (
            .in0(N__11141),
            .in1(N__11104),
            .in2(N__11174),
            .in3(N__11957),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.r_addr_1_LC_4_2_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_4_2_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.r_addr_1_LC_4_2_1  (
            .in0(N__11955),
            .in1(_gnd_net_),
            .in2(N__11108),
            .in3(N__11140),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_2  (
            .in0(_gnd_net_),
            .in1(N__11954),
            .in2(_gnd_net_),
            .in3(N__25880),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_3  (
            .in0(_gnd_net_),
            .in1(N__11076),
            .in2(_gnd_net_),
            .in3(N__11069),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(\uu2.trig_rd_is_det_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_0_LC_4_2_4 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_2_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.r_addr_0_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11112),
            .in3(N__11100),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.trig_rd_det_1_LC_4_2_5 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_4_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_4_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11070),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.trig_rd_det_0_LC_4_2_6 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_4_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_4_2_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_4_2_6  (
            .in0(_gnd_net_),
            .in1(N__14683),
            .in2(_gnd_net_),
            .in3(N__12137),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.r_addr_4_LC_4_2_7 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_2_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_4_LC_4_2_7  (
            .in0(N__11956),
            .in1(N__12007),
            .in2(_gnd_net_),
            .in3(N__11978),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26182),
            .ce(),
            .sr(N__25805));
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_4_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_4_3_0  (
            .in0(N__11314),
            .in1(N__11458),
            .in2(N__11265),
            .in3(N__11293),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_4_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_4_3_1  (
            .in0(N__11244),
            .in1(N__12193),
            .in2(N__11277),
            .in3(N__11373),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_3_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_4_3_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_4_3_2 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uu2.l_count_3_LC_4_3_2  (
            .in0(N__12207),
            .in1(N__11246),
            .in2(N__11274),
            .in3(N__11264),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26175),
            .ce(),
            .sr(N__25839));
    defparam \uu2.l_count_2_LC_4_3_3 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_4_3_3 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_4_3_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_2_LC_4_3_3  (
            .in0(N__11245),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12206),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26175),
            .ce(),
            .sr(N__25839));
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_3_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_4_3_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_4_3_4  (
            .in0(N__12192),
            .in1(N__11271),
            .in2(N__11469),
            .in3(N__11243),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_3_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_3_5  (
            .in0(N__11263),
            .in1(N__12191),
            .in2(N__11247),
            .in3(N__12171),
            .lcout(\uu2.un306_ci ),
            .ltout(\uu2.un306_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_4_3_6 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_4_3_6 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_4_3_6 .LUT_INIT=16'b0001001000010010;
    LogicCell40 \uu2.l_count_4_LC_4_3_6  (
            .in0(N__11411),
            .in1(N__11434),
            .in2(N__11226),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26175),
            .ce(),
            .sr(N__25839));
    defparam \uu2.l_count_5_LC_4_3_7 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_4_3_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_4_3_7 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \uu2.l_count_5_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__11410),
            .in2(N__11367),
            .in3(N__11460),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26175),
            .ce(),
            .sr(N__25839));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_4_4_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_4_4_0  (
            .in0(N__11330),
            .in1(N__11408),
            .in2(N__11388),
            .in3(N__12169),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_6_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_4_4_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_4_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.l_count_6_LC_4_4_1  (
            .in0(N__11345),
            .in1(N__11333),
            .in2(_gnd_net_),
            .in3(N__11362),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26167),
            .ce(),
            .sr(N__25836));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__11459),
            .in2(_gnd_net_),
            .in3(N__11409),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(\uu2.vbuf_count.un328_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_4_3  (
            .in0(N__11315),
            .in1(N__11332),
            .in2(N__11442),
            .in3(N__11361),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_4_4_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_4_4_4 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uu2.l_count_9_LC_4_4_4  (
            .in0(N__11387),
            .in1(N__11435),
            .in2(N__11415),
            .in3(N__11295),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26167),
            .ce(),
            .sr(N__25836));
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_4_4_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_4_4_5  (
            .in0(N__12170),
            .in1(N__11331),
            .in2(N__11412),
            .in3(N__11386),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_7_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_4_4_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_4_4_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.l_count_7_LC_4_4_6  (
            .in0(N__11363),
            .in1(N__11346),
            .in2(N__11337),
            .in3(N__11316),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26167),
            .ce(),
            .sr(N__25836));
    defparam \uu2.l_count_8_LC_4_4_7 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_4_4_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_4_4_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__11294),
            .in2(_gnd_net_),
            .in3(N__11301),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26167),
            .ce(),
            .sr(N__25836));
    defparam \Lab_UT.dispString.cnt_0_LC_4_5_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_4_5_2 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_4_5_2  (
            .in0(N__13680),
            .in1(N__13411),
            .in2(N__22070),
            .in3(N__13541),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26158),
            .ce(),
            .sr(N__25800));
    defparam \Lab_UT.dispString.cnt_1_LC_4_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_4_5_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_4_5_3  (
            .in0(N__13412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13540),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26158),
            .ce(),
            .sr(N__25800));
    defparam \Lab_UT.dispString.cnt_2_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_4_5_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_4_5_4  (
            .in0(N__12282),
            .in1(_gnd_net_),
            .in2(N__13699),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26158),
            .ce(),
            .sr(N__25800));
    defparam \uu0.sec_clk_LC_4_5_5 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_4_5_5 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_4_5_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.sec_clk_LC_4_5_5  (
            .in0(N__11598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14722),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26158),
            .ce(),
            .sr(N__25800));
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_5_6 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_4_5_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_4_5_6  (
            .in0(N__11514),
            .in1(N__11528),
            .in2(_gnd_net_),
            .in3(N__11597),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_1_LC_4_5_7 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_4_5_7 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_4_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.delay_line_1_LC_4_5_7  (
            .in0(N__11529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26158),
            .ce(),
            .sr(N__25800));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_6_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_6_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__11504),
            .in2(_gnd_net_),
            .in3(N__11615),
            .lcout(\buart.Z_tx.uart_busy_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_6_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_6_1 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_4_6_1  (
            .in0(N__11617),
            .in1(N__11681),
            .in2(N__11664),
            .in3(N__11642),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_4_6_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_4_6_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_4_6_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_4_6_2  (
            .in0(N__12098),
            .in1(N__11645),
            .in2(N__11508),
            .in3(N__11505),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26151),
            .ce(),
            .sr(N__25829));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_6_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_6_3 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_6_3  (
            .in0(N__11658),
            .in1(N__11496),
            .in2(N__11682),
            .in3(N__11490),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_6_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_6_4 .LUT_INIT=16'b1010101010011010;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_4_6_4  (
            .in0(N__11680),
            .in1(N__11659),
            .in2(N__11688),
            .in3(N__11616),
            .lcout(),
            .ltout(\buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_4_6_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_4_6_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_4_6_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11685),
            .in3(N__12093),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26151),
            .ce(),
            .sr(N__25829));
    defparam \buart.Z_tx.bitcount_1_LC_4_6_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_4_6_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_4_6_6 .LUT_INIT=16'b1111110011110110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_4_6_6  (
            .in0(N__11643),
            .in1(N__11663),
            .in2(N__12119),
            .in3(N__11619),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26151),
            .ce(),
            .sr(N__25829));
    defparam \buart.Z_tx.bitcount_0_LC_4_6_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_4_6_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_4_6_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_4_6_7  (
            .in0(N__11618),
            .in1(N__12094),
            .in2(_gnd_net_),
            .in3(N__11644),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26151),
            .ce(),
            .sr(N__25829));
    defparam \buart.Z_rx.shifter_2_rep2_RNICDH61_LC_4_7_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep2_RNICDH61_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_2_rep2_RNICDH61_LC_4_7_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep2_RNICDH61_LC_4_7_0  (
            .in0(N__18891),
            .in1(N__21779),
            .in2(N__18141),
            .in3(N__13883),
            .lcout(\buart.Z_rx.G_17_i_a5_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__13413),
            .in2(_gnd_net_),
            .in3(N__13543),
            .lcout(\Lab_UT.dispString.N_30_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m4_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m4_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m4_LC_4_8_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dispString.m4_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(N__14953),
            .in2(_gnd_net_),
            .in3(N__14894),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m71_0_LC_4_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m71_0_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m71_0_LC_4_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.m71_0_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(N__18910),
            .in2(_gnd_net_),
            .in3(N__25503),
            .lcout(\Lab_UT.dictrl.m71Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_12_a6_3_7_LC_4_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_12_a6_3_7_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_12_a6_3_7_LC_4_9_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_12_a6_3_7_LC_4_9_0  (
            .in0(N__19017),
            .in1(N__21749),
            .in2(N__19190),
            .in3(N__26348),
            .lcout(\Lab_UT.dictrl.g0_12_a6_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIH0Q52_5_LC_4_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIH0Q52_5_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIH0Q52_5_LC_4_9_1 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \buart.Z_rx.shifter_RNIH0Q52_5_LC_4_9_1  (
            .in0(N__19157),
            .in1(N__13329),
            .in2(N__13790),
            .in3(N__19018),
            .lcout(N_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_25_LC_4_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_25_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_25_LC_4_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_25_LC_4_9_3  (
            .in0(N__26349),
            .in1(N__19019),
            .in2(N__19192),
            .in3(N__11700),
            .lcout(\Lab_UT.dictrl.N_97_mux_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF4VT_0_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF4VT_0_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF4VT_0_LC_4_10_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIF4VT_0_LC_4_10_0  (
            .in0(N__19423),
            .in1(N__20360),
            .in2(N__18585),
            .in3(N__16592),
            .lcout(\Lab_UT.dictrl.g0_12_o6_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIMFOD2_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIMFOD2_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIMFOD2_LC_4_10_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIMFOD2_LC_4_10_1  (
            .in0(N__14832),
            .in1(N__17096),
            .in2(_gnd_net_),
            .in3(N__19917),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_13_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIJT0P3_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIJT0P3_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIJT0P3_LC_4_10_2 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNIJT0P3_LC_4_10_2  (
            .in0(N__11709),
            .in1(N__19710),
            .in2(N__11703),
            .in3(N__16829),
            .lcout(\Lab_UT.dictrl.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIOEMF_0_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIOEMF_0_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIOEMF_0_LC_4_10_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIOEMF_0_LC_4_10_3  (
            .in0(N__16593),
            .in1(N__14833),
            .in2(N__12684),
            .in3(N__12725),
            .lcout(\Lab_UT.dictrl.N_17_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m34_4_2_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m34_4_2_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m34_4_2_LC_4_10_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.m34_4_2_LC_4_10_4  (
            .in0(N__17094),
            .in1(N__12677),
            .in2(_gnd_net_),
            .in3(N__14045),
            .lcout(\Lab_UT.dictrl.m34_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m59_1_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m59_1_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m59_1_LC_4_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m59_1_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(N__12721),
            .in2(_gnd_net_),
            .in3(N__14046),
            .lcout(Lab_UT_dictrl_m59_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_10_3_LC_4_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_10_3_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_10_3_LC_4_10_7 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \Lab_UT.dictrl.g0_10_3_LC_4_10_7  (
            .in0(N__12678),
            .in1(N__17095),
            .in2(N__12726),
            .in3(N__19424),
            .lcout(\Lab_UT.dictrl.g0_10Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIOIIC1_LC_4_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIOIIC1_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIOIIC1_LC_4_11_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIOIIC1_LC_4_11_0  (
            .in0(N__13963),
            .in1(N__11694),
            .in2(N__20488),
            .in3(N__15636),
            .lcout(\Lab_UT.dictrl.m34_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_12_o3_2_LC_4_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_12_o3_2_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_12_o3_2_LC_4_11_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g0_12_o3_2_LC_4_11_2  (
            .in0(N__18729),
            .in1(N__13877),
            .in2(_gnd_net_),
            .in3(N__13956),
            .lcout(\Lab_UT.dictrl.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_17_LC_4_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_17_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_17_LC_4_11_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_17_LC_4_11_3  (
            .in0(N__13957),
            .in1(N__18730),
            .in2(N__13887),
            .in3(N__20267),
            .lcout(\Lab_UT.dictrl.g1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_4_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_4_11_4 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_13_LC_4_11_4  (
            .in0(N__20268),
            .in1(N__13881),
            .in2(N__18752),
            .in3(N__13959),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_4_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_4_11_5 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_6_LC_4_11_5  (
            .in0(N__19149),
            .in1(N__21770),
            .in2(N__11712),
            .in3(N__14371),
            .lcout(\Lab_UT.dictrl.N_15_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_4_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_4_11_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_8_LC_4_11_6  (
            .in0(N__13882),
            .in1(N__13958),
            .in2(N__18751),
            .in3(N__24011),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_a7_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep2_RNIDJQN_LC_4_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep2_RNIDJQN_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep2_RNIDJQN_LC_4_12_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \buart.Z_rx.shifter_1_rep2_RNIDJQN_LC_4_12_0  (
            .in0(N__18994),
            .in1(N__18750),
            .in2(N__19150),
            .in3(N__13964),
            .lcout(\buart.Z_rx.G_17_i_a5_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_5_1_LC_4_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_5_1_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_5_1_LC_4_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_5_1_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__19115),
            .in2(_gnd_net_),
            .in3(N__18995),
            .lcout(\Lab_UT.dictrl.g0_i_a4_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_LC_4_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_4_12_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_4_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_5_LC_4_12_2  (
            .in0(N__19116),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_6_LC_4_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_4_12_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18137),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_fast_5_LC_4_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_4_12_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_4_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_4_12_4  (
            .in0(N__19117),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_fast_4_LC_4_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_4_12_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_4_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18998),
            .lcout(bu_rx_data_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_12_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_rep1_LC_4_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_4_rep1_LC_4_12_6  (
            .in0(N__18996),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_4_rep2_LC_4_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep2_LC_4_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_rep2_LC_4_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_rep2_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18997),
            .lcout(bu_rx_data_4_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26122),
            .ce(N__14241),
            .sr(N__25835));
    defparam \buart.Z_rx.shifter_0_rep1_LC_4_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_LC_4_13_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_rep1_LC_4_13_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_LC_4_13_0  (
            .in0(N__25457),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_fast_0_LC_4_13_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_4_13_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(N__25456),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_13_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_4_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26649),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_fast_1_LC_4_13_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_4_13_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_4_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_4_13_3  (
            .in0(N__26650),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_fast_7_LC_4_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_4_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_4_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11748),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_4_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_4_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26330),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_3_LC_4_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_4_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_4_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18933),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \buart.Z_rx.shifter_fast_2_LC_4_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_4_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26331),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26120),
            .ce(N__14240),
            .sr(N__25838));
    defparam \Lab_UT.dictrl.g0_9_3_LC_4_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_9_3_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_9_3_LC_4_14_0 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \Lab_UT.dictrl.g0_9_3_LC_4_14_0  (
            .in0(N__12783),
            .in1(N__12829),
            .in2(N__12762),
            .in3(N__12996),
            .lcout(\Lab_UT.dictrl.g0_9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_LC_4_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_LC_4_14_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.g0_i_m2_1_o6_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__12754),
            .in2(_gnd_net_),
            .in3(N__12781),
            .lcout(\Lab_UT.dictrl.N_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m23_a0_LC_4_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m23_a0_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m23_a0_LC_4_14_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \Lab_UT.dictrl.m23_a0_LC_4_14_2  (
            .in0(N__12782),
            .in1(_gnd_net_),
            .in2(N__12761),
            .in3(N__12995),
            .lcout(\Lab_UT.dictrl.m23_aZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m40_1_LC_4_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m40_1_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m40_1_LC_4_14_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.dictrl.m40_1_LC_4_14_3  (
            .in0(N__12994),
            .in1(N__12753),
            .in2(N__14108),
            .in3(N__12780),
            .lcout(\Lab_UT.dictrl.m40Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.m40Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_4_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_4_14_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_4_14_4  (
            .in0(N__18931),
            .in1(N__22819),
            .in2(N__11799),
            .in3(N__20577),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_4_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_4_14_5 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_4_14_5  (
            .in0(N__11796),
            .in1(N__17238),
            .in2(N__11784),
            .in3(N__19473),
            .lcout(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_3_LC_4_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_4_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_4_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_4_14_6  (
            .in0(N__18932),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26118),
            .ce(N__14238),
            .sr(N__25840));
    defparam \Lab_UT.dictrl.g0_8_LC_4_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_8_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_8_LC_4_15_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_8_LC_4_15_0  (
            .in0(N__20296),
            .in1(N__18595),
            .in2(N__11781),
            .in3(N__20406),
            .lcout(\Lab_UT.dictrl.N_97_mux_0 ),
            .ltout(\Lab_UT.dictrl.N_97_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_10_LC_4_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_10_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_10_LC_4_15_1 .LUT_INIT=16'b0000111111101110;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_10_LC_4_15_1  (
            .in0(N__11901),
            .in1(N__11772),
            .in2(N__11763),
            .in3(N__19735),
            .lcout(\Lab_UT.dictrl.N_2435_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_18_LC_4_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_18_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_18_LC_4_15_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_18_LC_4_15_2  (
            .in0(N__20493),
            .in1(N__20402),
            .in2(N__20045),
            .in3(N__19446),
            .lcout(\Lab_UT.dictrl.g1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_20_LC_4_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_20_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_20_LC_4_15_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_20_LC_4_15_3  (
            .in0(N__19447),
            .in1(N__18594),
            .in2(N__20409),
            .in3(N__20295),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_16_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_12_LC_4_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_12_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_12_LC_4_15_4 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_12_LC_4_15_4  (
            .in0(N__12840),
            .in1(N__11895),
            .in2(N__11889),
            .in3(N__20576),
            .lcout(\Lab_UT.dictrl.N_2446_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_5_1_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_5_1_0 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_5_1_0  (
            .in0(N__23606),
            .in1(N__12041),
            .in2(N__23692),
            .in3(N__23381),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_5_1_1 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_5_1_1 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_5_1_1  (
            .in0(N__11855),
            .in1(N__23668),
            .in2(_gnd_net_),
            .in3(N__23603),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_5_1_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_5_1_2  (
            .in0(N__23604),
            .in1(N__17551),
            .in2(N__23691),
            .in3(N__23490),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_1_LC_5_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_5_1_3 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_user_1_LC_5_1_3  (
            .in0(N__20959),
            .in1(_gnd_net_),
            .in2(N__12048),
            .in3(N__17555),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__20843));
    defparam \uu2.w_addr_user_2_LC_5_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_5_1_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_2_LC_5_1_4  (
            .in0(N__17556),
            .in1(N__12047),
            .in2(N__17522),
            .in3(N__20960),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__20843));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_1_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_5_1_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_5_1_5  (
            .in0(N__17513),
            .in1(N__23669),
            .in2(N__17376),
            .in3(N__23605),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_0_LC_5_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_5_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_5_1_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_user_0_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__12043),
            .in2(_gnd_net_),
            .in3(N__20958),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__20843));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_5_1_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_5_1_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_5_1_7  (
            .in0(N__12042),
            .in1(N__17514),
            .in2(N__17559),
            .in3(N__13089),
            .lcout(\uu2.un404_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_5_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI1VU6_3_LC_5_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI1VU6_3_LC_5_2_0  (
            .in0(N__21050),
            .in1(N__13077),
            .in2(N__14420),
            .in3(N__12039),
            .lcout(\uu2.un3_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_5_2_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_5_2_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__14415),
            .in2(_gnd_net_),
            .in3(N__20882),
            .lcout(),
            .ltout(\uu2.vbuf_w_addr_user.un448_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_5_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_5_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_5_2_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_5_2_2  (
            .in0(N__23533),
            .in1(N__20921),
            .in2(N__12051),
            .in3(N__20894),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12147),
            .sr(N__20842));
    defparam \uu2.w_addr_user_nesr_3_LC_5_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_5_2_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_5_2_3  (
            .in0(N__12040),
            .in1(N__17518),
            .in2(N__13087),
            .in3(N__17557),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12147),
            .sr(N__20842));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_5_2_4 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_5_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_5_2_4  (
            .in0(N__21051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21014),
            .lcout(\uu2.un426_ci_3 ),
            .ltout(\uu2.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_7_LC_5_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_5_2_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_5_2_5  (
            .in0(N__20920),
            .in1(N__14416),
            .in2(N__12018),
            .in3(N__20883),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12147),
            .sr(N__20842));
    defparam \uu2.r_addr_5_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_5_3_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_5_3_0  (
            .in0(N__12014),
            .in1(N__11982),
            .in2(N__11930),
            .in3(N__11958),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26168),
            .ce(),
            .sr(N__25806));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_5_3_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_5_3_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__12261),
            .in2(_gnd_net_),
            .in3(N__12237),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_5_3_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__12194),
            .in2(_gnd_net_),
            .in3(N__12172),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_1_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_5_3_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_5_3_4 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.l_count_1_LC_5_3_4  (
            .in0(N__12174),
            .in1(_gnd_net_),
            .in2(N__12198),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26168),
            .ce(),
            .sr(N__25806));
    defparam \uu2.l_count_0_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_5_3_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_5_3_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12173),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26168),
            .ce(),
            .sr(N__25806));
    defparam \uu2.w_addr_displaying_nesr_RNO_0_5_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNO_0_5_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNO_0_5_LC_5_3_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNO_0_5_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__16726),
            .in2(_gnd_net_),
            .in3(N__25019),
            .lcout(\uu2.un21_w_addr_displaying_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNID65PE_2_LC_5_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNID65PE_2_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNID65PE_2_LC_5_3_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_user_RNID65PE_2_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__20947),
            .in2(_gnd_net_),
            .in3(N__20823),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_5_4_0 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_5_4_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_5_4_0  (
            .in0(N__14684),
            .in1(N__12138),
            .in2(N__12114),
            .in3(N__25881),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26159),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_5_4_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_5_4_1 .LUT_INIT=16'b0000000111111111;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_5_4_1  (
            .in0(N__13409),
            .in1(N__13542),
            .in2(N__12315),
            .in3(N__12303),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26159),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_5_4_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_5_4_4 .LUT_INIT=16'b1111010111100101;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_5_4_4  (
            .in0(N__13678),
            .in1(N__22069),
            .in2(N__12297),
            .in3(N__13410),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26159),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_5_4_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_5_4_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__12370),
            .in2(_gnd_net_),
            .in3(N__12354),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_5_4_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_5_4_7 .LUT_INIT=16'b1111111001110111;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_5_4_7  (
            .in0(N__13408),
            .in1(N__13679),
            .in2(N__22090),
            .in3(N__12288),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26159),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_5_0 .LUT_INIT=16'b0010011101110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_5_5_0  (
            .in0(N__13672),
            .in1(N__21195),
            .in2(N__22065),
            .in3(N__16287),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_2_tz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_5_5_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_5_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_5_5_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_1_LC_5_5_1  (
            .in0(N__13671),
            .in1(N__12468),
            .in2(_gnd_net_),
            .in3(N__12421),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_5_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_5_2 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_5_5_2  (
            .in0(N__13403),
            .in1(N__13538),
            .in2(N__12306),
            .in3(N__12267),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_5_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_5_5_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_2_LC_5_5_3  (
            .in0(N__13536),
            .in1(N__12467),
            .in2(_gnd_net_),
            .in3(N__12420),
            .lcout(\Lab_UT.dispString.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_5_5 .LUT_INIT=16'b0001010100000101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_5_5_5  (
            .in0(N__13537),
            .in1(N__12469),
            .in2(N__13433),
            .in3(N__12423),
            .lcout(\Lab_UT.dispString.m74_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_5_6 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_5_LC_5_5_6  (
            .in0(N__12422),
            .in1(N__13404),
            .in2(N__12474),
            .in3(N__13539),
            .lcout(\Lab_UT.dispString.m77_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_5_5_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_5_5_7 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_5_5_7  (
            .in0(N__12281),
            .in1(N__13626),
            .in2(N__13688),
            .in3(N__21225),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_5_6_1 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_5_6_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__12510),
            .in2(_gnd_net_),
            .in3(N__14718),
            .lcout(oneSecStrb),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNI7F27_0_LC_5_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNI7F27_0_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNI7F27_0_LC_5_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Lab_UT.dispString.cnt_RNI7F27_0_LC_5_6_3  (
            .in0(N__13535),
            .in1(N__12454),
            .in2(_gnd_net_),
            .in3(N__12408),
            .lcout(\Lab_UT.dispString.N_23_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_5_7_0 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_5_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.sec_clkD_LC_5_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14727),
            .lcout(\uu0.sec_clkDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26137),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m57_LC_5_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m57_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m57_LC_5_7_1 .LUT_INIT=16'b0001000100001100;
    LogicCell40 \Lab_UT.dispString.m57_LC_5_7_1  (
            .in0(N__17865),
            .in1(N__12528),
            .in2(N__12419),
            .in3(N__12452),
            .lcout(\Lab_UT.m57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m60_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m60_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m60_LC_5_7_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dispString.m60_LC_5_7_2  (
            .in0(N__12451),
            .in1(N__16720),
            .in2(_gnd_net_),
            .in3(N__12402),
            .lcout(G_216),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.alarmstate_1_0_i_1_LC_5_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.alarmstate_1_0_i_1_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.alarmstate_1_0_i_1_LC_5_7_3 .LUT_INIT=16'b1111001000100010;
    LogicCell40 \Lab_UT.dispString.alarmstate_1_0_i_1_LC_5_7_3  (
            .in0(N__12407),
            .in1(N__12579),
            .in2(N__12473),
            .in3(N__17864),
            .lcout(),
            .ltout(\Lab_UT.alarmstate_1_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_7_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_1_LC_5_7_4  (
            .in0(N__12418),
            .in1(N__12492),
            .in2(N__12504),
            .in3(N__12498),
            .lcout(G_215),
            .ltout(G_215_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.alarmstate_1_sqmuxa_1_i_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.alarmstate_1_sqmuxa_1_i_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.alarmstate_1_sqmuxa_1_i_LC_5_7_5 .LUT_INIT=16'b1100111111111111;
    LogicCell40 \Lab_UT.dispString.alarmstate_1_sqmuxa_1_i_LC_5_7_5  (
            .in0(_gnd_net_),
            .in1(N__16719),
            .in2(N__12501),
            .in3(N__12450),
            .lcout(G_214),
            .ltout(G_214_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_7_6 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_0_LC_5_7_6  (
            .in0(N__12453),
            .in1(N__12491),
            .in2(N__12483),
            .in3(N__12480),
            .lcout(G_213),
            .ltout(G_213_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_0_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_0_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_0_LC_5_7_7 .LUT_INIT=16'b0000000010101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_0_LC_5_7_7  (
            .in0(N__12406),
            .in1(_gnd_net_),
            .in2(N__12375),
            .in3(N__13555),
            .lcout(\Lab_UT.dispString.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m71_LC_5_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m71_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m71_LC_5_8_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m71_LC_5_8_2  (
            .in0(N__25899),
            .in1(N__26693),
            .in2(N__12624),
            .in3(N__13995),
            .lcout(N_105_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m54_e_LC_5_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m54_e_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m54_e_LC_5_8_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dispString.m54_e_LC_5_8_3  (
            .in0(N__14952),
            .in1(N__14893),
            .in2(_gnd_net_),
            .in3(N__12527),
            .lcout(\Lab_UT.dispString.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI0RBN1_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI0RBN1_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI0RBN1_LC_5_9_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNI0RBN1_LC_5_9_0  (
            .in0(N__19720),
            .in1(N__13773),
            .in2(N__18157),
            .in3(N__22977),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_12_a6_3_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI70I48_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI70I48_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI70I48_LC_5_9_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNI70I48_LC_5_9_1  (
            .in0(N__12573),
            .in1(N__17193),
            .in2(N__12567),
            .in3(N__12564),
            .lcout(\Lab_UT.dictrl.g0_12_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI0UI65_3_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0UI65_3_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0UI65_3_LC_5_9_2 .LUT_INIT=16'b0000100011001000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI0UI65_3_LC_5_9_2  (
            .in0(N__12558),
            .in1(N__12633),
            .in2(N__24547),
            .in3(N__12552),
            .lcout(\Lab_UT.dictrl.N_23_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNINKC83_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNINKC83_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNINKC83_LC_5_10_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_esr_RNINKC83_LC_5_10_0  (
            .in0(N__12642),
            .in1(N__18630),
            .in2(N__15096),
            .in3(N__16833),
            .lcout(\Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_19_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_19_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_19_LC_5_10_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_19_LC_5_10_1  (
            .in0(N__19422),
            .in1(N__15627),
            .in2(N__20375),
            .in3(N__20283),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_11_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_11_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_11_LC_5_10_2 .LUT_INIT=16'b0000000010110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_11_LC_5_10_2  (
            .in0(N__18650),
            .in1(N__26371),
            .in2(N__12546),
            .in3(N__18559),
            .lcout(\Lab_UT.dictrl.m63_d_0_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m107_e_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m107_e_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m107_e_LC_5_10_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dispString.m107_e_LC_5_10_3  (
            .in0(N__19421),
            .in1(N__20282),
            .in2(N__12903),
            .in3(N__18649),
            .lcout(\Lab_UT.dispString.N_112_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI3S8S_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI3S8S_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI3S8S_LC_5_11_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_RNI3S8S_LC_5_11_0  (
            .in0(N__15336),
            .in1(N__15628),
            .in2(N__14834),
            .in3(N__14057),
            .lcout(\Lab_UT.dictrl.g0_12_a6_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_12_o6_1_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_12_o6_1_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_12_o6_1_LC_5_11_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.g0_12_o6_1_LC_5_11_1  (
            .in0(N__25501),
            .in1(N__26667),
            .in2(N__18919),
            .in3(N__13990),
            .lcout(\Lab_UT.dictrl.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_1_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_1_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_1_LC_5_11_2 .LUT_INIT=16'b0011000101110011;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_1_LC_5_11_2  (
            .in0(N__26668),
            .in1(N__26372),
            .in2(N__22820),
            .in3(N__25502),
            .lcout(\Lab_UT.dictrl.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFP8P_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFP8P_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFP8P_LC_5_11_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFP8P_LC_5_11_3  (
            .in0(N__15629),
            .in1(N__14824),
            .in2(_gnd_net_),
            .in3(N__17093),
            .lcout(\Lab_UT.dictrl.m27_d_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_5_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_5_11_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_7_LC_5_11_4  (
            .in0(N__19445),
            .in1(N__15630),
            .in2(N__15342),
            .in3(N__18232),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_a7_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_LC_5_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_LC_5_12_0 .LUT_INIT=16'b0000110100000101;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_LC_5_12_0  (
            .in0(N__16832),
            .in1(N__18346),
            .in2(N__24053),
            .in3(N__14828),
            .lcout(\Lab_UT.dictrl.N_1110_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0H5_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0H5_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0H5_LC_5_12_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0H5_LC_5_12_1  (
            .in0(N__14825),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24003),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDC4_LC_5_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDC4_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDC4_LC_5_12_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDC4_LC_5_12_2  (
            .in0(N__15528),
            .in1(N__18347),
            .in2(N__12636),
            .in3(N__14481),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_1_LC_5_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_1_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_1_LC_5_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_1_LC_5_12_3  (
            .in0(N__14826),
            .in1(N__24004),
            .in2(N__18348),
            .in3(N__16830),
            .lcout(\Lab_UT.dictrl.G_17_i_a5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_0_LC_5_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_0_LC_5_12_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_0_LC_5_12_4  (
            .in0(N__16831),
            .in1(N__18345),
            .in2(N__24054),
            .in3(N__14827),
            .lcout(),
            .ltout(G_17_i_a5_2_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep2_RNI1CHAB_LC_5_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep2_RNI1CHAB_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep2_RNI1CHAB_LC_5_12_5 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \buart.Z_rx.shifter_1_rep2_RNI1CHAB_LC_5_12_5  (
            .in0(N__12804),
            .in1(N__12798),
            .in2(N__12786),
            .in3(N__12849),
            .lcout(G_17_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_e_LC_5_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_e_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_e_LC_5_12_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m22_e_LC_5_12_6  (
            .in0(_gnd_net_),
            .in1(N__12779),
            .in2(_gnd_net_),
            .in3(N__12752),
            .lcout(\Lab_UT.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_9_LC_5_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_9_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_9_LC_5_13_0 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_9_LC_5_13_0  (
            .in0(N__12710),
            .in1(N__12670),
            .in2(_gnd_net_),
            .in3(N__15411),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_7_LC_5_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_7_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_7_LC_5_13_1 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_7_LC_5_13_1  (
            .in0(N__14333),
            .in1(N__18337),
            .in2(N__12735),
            .in3(N__12732),
            .lcout(\Lab_UT.dictrl.m53_d_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_10_LC_5_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_10_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_10_LC_5_13_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_10_LC_5_13_2  (
            .in0(N__14149),
            .in1(N__13002),
            .in2(N__14107),
            .in3(N__14282),
            .lcout(\Lab_UT.dictrl.g2_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_9_LC_5_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_9_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_9_LC_5_13_3 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_9_LC_5_13_3  (
            .in0(N__15412),
            .in1(_gnd_net_),
            .in2(N__12682),
            .in3(N__12711),
            .lcout(\Lab_UT.dictrl.g2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_9_LC_5_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_9_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_9_LC_5_13_4 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_9_LC_5_13_4  (
            .in0(N__12709),
            .in1(N__12669),
            .in2(_gnd_net_),
            .in3(N__15410),
            .lcout(\Lab_UT.dictrl.g2_0_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_9_LC_5_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_9_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_9_LC_5_13_5 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_9_LC_5_13_5  (
            .in0(N__15413),
            .in1(_gnd_net_),
            .in2(N__12683),
            .in3(N__12712),
            .lcout(\Lab_UT.dictrl.g2_0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIMUEI_LC_5_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIMUEI_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIMUEI_LC_5_13_6 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIMUEI_LC_5_13_6  (
            .in0(N__12708),
            .in1(N__12668),
            .in2(_gnd_net_),
            .in3(N__15606),
            .lcout(\Lab_UT.dictrl.g2_0_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m107_e_3_LC_5_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m107_e_3_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m107_e_3_LC_5_13_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dispString.m107_e_3_LC_5_13_7  (
            .in0(N__14150),
            .in1(N__14056),
            .in2(N__12888),
            .in3(N__14276),
            .lcout(\Lab_UT.dispString.m107_eZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m18_LC_5_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m18_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m18_LC_5_14_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \Lab_UT.dictrl.m18_LC_5_14_0  (
            .in0(N__12827),
            .in1(N__12889),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m12_1_LC_5_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m12_1_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m12_1_LC_5_14_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.m12_1_LC_5_14_1  (
            .in0(N__12891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12828),
            .lcout(\Lab_UT.dictrl.m12Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_0_LC_5_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_0_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_i_m2_1_o6_0_LC_5_14_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.g0_i_m2_1_o6_0_LC_5_14_2  (
            .in0(N__14094),
            .in1(N__12890),
            .in2(N__12833),
            .in3(N__14277),
            .lcout(\Lab_UT.dictrl.N_10_1 ),
            .ltout(\Lab_UT.dictrl.N_10_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI5GLB2_LC_5_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI5GLB2_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI5GLB2_LC_5_14_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNI5GLB2_LC_5_14_3  (
            .in0(N__15631),
            .in1(N__18759),
            .in2(N__12867),
            .in3(N__24002),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI60US8_0_LC_5_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI60US8_0_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI60US8_0_LC_5_14_4 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI60US8_0_LC_5_14_4  (
            .in0(N__12864),
            .in1(N__13014),
            .in2(N__12852),
            .in3(N__12957),
            .lcout(N_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_21_LC_5_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_21_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_21_LC_5_14_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_21_LC_5_14_7  (
            .in0(N__15632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18341),
            .lcout(\Lab_UT.dictrl.N_1105_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI12QU_3_LC_5_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI12QU_3_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI12QU_3_LC_5_15_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI12QU_3_LC_5_15_0  (
            .in0(N__20394),
            .in1(N__12834),
            .in2(N__18603),
            .in3(N__15421),
            .lcout(\Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIB5Q7_0_LC_5_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIB5Q7_0_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIB5Q7_0_LC_5_15_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIB5Q7_0_LC_5_15_1  (
            .in0(N__24000),
            .in1(_gnd_net_),
            .in2(N__15422),
            .in3(N__16601),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF3PO3_0_LC_5_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF3PO3_0_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIF3PO3_0_LC_5_15_2 .LUT_INIT=16'b1011000110100000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIF3PO3_0_LC_5_15_2  (
            .in0(N__13023),
            .in1(N__12968),
            .in2(N__13017),
            .in3(N__13008),
            .lcout(\Lab_UT.dictrl.g0_i_m2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNITRQM_2_LC_5_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNITRQM_2_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNITRQM_2_LC_5_15_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNITRQM_2_LC_5_15_3  (
            .in0(N__23999),
            .in1(N__13001),
            .in2(N__15423),
            .in3(N__15366),
            .lcout(\Lab_UT.dictrl.g0_i_m2_1_a6_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIO0FK_3_LC_5_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIO0FK_3_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIO0FK_3_LC_5_15_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIO0FK_3_LC_5_15_4  (
            .in0(N__13000),
            .in1(N__15414),
            .in2(_gnd_net_),
            .in3(N__24001),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTO82_0_LC_5_15_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTO82_0_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTO82_0_LC_5_15_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIQTO82_0_LC_5_15_5  (
            .in0(N__12969),
            .in1(N__16602),
            .in2(N__12960),
            .in3(N__14487),
            .lcout(\Lab_UT.dictrl.G_17_i_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_1_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_6_1_0 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_6_1_0  (
            .in0(N__13238),
            .in1(N__15775),
            .in2(N__12930),
            .in3(N__14522),
            .lcout(\uu2.mem0.N_66_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_1_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_6_1_1 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_6_1_1  (
            .in0(N__15773),
            .in1(N__12929),
            .in2(_gnd_net_),
            .in3(N__13200),
            .lcout(\uu2.mem0.N_56_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI1R353_0_LC_6_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI1R353_0_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI1R353_0_LC_6_1_2 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI1R353_0_LC_6_1_2  (
            .in0(N__23488),
            .in1(N__23362),
            .in2(N__14568),
            .in3(N__23403),
            .lcout(\uu2.N_95_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI1R353_0_0_LC_6_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI1R353_0_0_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI1R353_0_0_LC_6_1_3 .LUT_INIT=16'b0000100010000000;
    LogicCell40 \uu2.w_addr_displaying_RNI1R353_0_0_LC_6_1_3  (
            .in0(N__23402),
            .in1(N__14563),
            .in2(N__23373),
            .in3(N__23489),
            .lcout(\uu2.N_96_mux ),
            .ltout(\uu2.N_96_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_6_1_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_6_1_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_6_1_4  (
            .in0(N__13161),
            .in1(_gnd_net_),
            .in2(N__12918),
            .in3(N__15774),
            .lcout(\uu2.mem0.N_63_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_6_1_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_6_1_5 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_6_1_5  (
            .in0(N__15776),
            .in1(N__13128),
            .in2(N__14526),
            .in3(N__13179),
            .lcout(\uu2.mem0.N_69_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_1_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_6_1_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_6_1_6  (
            .in0(N__13127),
            .in1(N__13287),
            .in2(_gnd_net_),
            .in3(N__15777),
            .lcout(\uu2.mem0.N_71_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_1_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_6_1_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_6_1_7  (
            .in0(N__23404),
            .in1(N__14567),
            .in2(_gnd_net_),
            .in3(N__23487),
            .lcout(\uu2.mem0.N_91_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_2_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_6_2_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_6_2_0  (
            .in0(N__23592),
            .in1(N__13110),
            .in2(N__23706),
            .in3(N__13266),
            .lcout(\uu2.mem0.N_50_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_6_2_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_6_2_1 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_6_2_1  (
            .in0(N__20762),
            .in1(N__23697),
            .in2(N__13088),
            .in3(N__23590),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_2_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_6_2_2 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_6_2_2  (
            .in0(N__23591),
            .in1(N__21013),
            .in2(N__23705),
            .in3(N__17413),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIB6L01_4_LC_6_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIB6L01_4_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIB6L01_4_LC_6_2_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIB6L01_4_LC_6_2_3  (
            .in0(N__20761),
            .in1(_gnd_net_),
            .in2(N__17420),
            .in3(N__17374),
            .lcout(\uu2.N_75_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNO_0_4_LC_6_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNO_0_4_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNO_0_4_LC_6_2_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.w_addr_displaying_RNO_0_4_LC_6_2_4  (
            .in0(N__23473),
            .in1(N__20763),
            .in2(N__23380),
            .in3(N__25028),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_6_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_6_2_5 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu2.w_addr_displaying_4_LC_6_2_5  (
            .in0(N__17414),
            .in1(_gnd_net_),
            .in2(N__13026),
            .in3(N__17375),
            .lcout(\uu2.w_addr_displayingZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__25767));
    defparam \uu2.w_addr_displaying_RNI2HHB1_4_LC_6_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI2HHB1_4_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI2HHB1_4_LC_6_2_6 .LUT_INIT=16'b0100100011100000;
    LogicCell40 \uu2.w_addr_displaying_RNI2HHB1_4_LC_6_2_6  (
            .in0(N__23472),
            .in1(N__17409),
            .in2(N__17381),
            .in3(N__20760),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_LC_6_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_6_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_6_2_7 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \uu2.w_addr_displaying_2_LC_6_2_7  (
            .in0(N__25029),
            .in1(N__23474),
            .in2(N__17377),
            .in3(N__23372),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__25767));
    defparam \uu2.un1_w_user_lf_LC_6_3_0 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_LC_6_3_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.un1_w_user_lf_LC_6_3_0  (
            .in0(N__13193),
            .in1(N__13212),
            .in2(N__13239),
            .in3(N__13175),
            .lcout(\uu2.un1_w_user_lf_0 ),
            .ltout(\uu2.un1_w_user_lf_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_6_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI93NG7_2_LC_6_3_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uu2.w_addr_user_RNI93NG7_2_LC_6_3_1  (
            .in0(N__23642),
            .in1(N__17468),
            .in2(N__13215),
            .in3(N__23578),
            .lcout(\uu2.un28_w_addr_user_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_6_3_2 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_6_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_6_3_2  (
            .in0(N__13261),
            .in1(N__13157),
            .in2(N__13286),
            .in3(N__13298),
            .lcout(\uu2.un1_w_user_lfZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI43E87_2_LC_6_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI43E87_2_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI43E87_2_LC_6_3_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uu2.w_addr_user_RNI43E87_2_LC_6_3_3  (
            .in0(N__25872),
            .in1(N__13206),
            .in2(N__17472),
            .in3(N__23579),
            .lcout(\uu2.w_addr_user_RNI43E87Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.m35_4_LC_6_3_4 .C_ON=1'b0;
    defparam \uu2.m35_4_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.m35_4_LC_6_3_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.m35_4_LC_6_3_4  (
            .in0(N__13192),
            .in1(N__13297),
            .in2(N__13265),
            .in3(N__13174),
            .lcout(),
            .ltout(\uu2.m35Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.m35_LC_6_3_5 .C_ON=1'b0;
    defparam \uu2.m35_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.m35_LC_6_3_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.m35_LC_6_3_5  (
            .in0(N__13156),
            .in1(N__13234),
            .in2(N__13143),
            .in3(N__13279),
            .lcout(\uu2.un1_w_user_cr_0 ),
            .ltout(\uu2.un1_w_user_cr_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_0_LC_6_3_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.un4_w_user_data_rdy_0_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13140),
            .in3(N__23641),
            .lcout(\uu2.un4_w_user_data_rdyZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_6_3_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_6_3_7  (
            .in0(N__13299),
            .in1(N__23662),
            .in2(_gnd_net_),
            .in3(N__23580),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_6_4_1 .LUT_INIT=16'b1100101011001111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_6_4_1  (
            .in0(N__13569),
            .in1(N__13308),
            .in2(N__13454),
            .in3(N__17832),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_6_4_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_6_4_2 .LUT_INIT=16'b0011111100001100;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__13701),
            .in2(N__13302),
            .in3(N__13617),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_6_4_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_6_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dispString.rdy_LC_6_4_3  (
            .in0(N__13570),
            .in1(N__22089),
            .in2(N__13455),
            .in3(N__13704),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_6_4_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_6_4_5 .LUT_INIT=16'b0001000111011101;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_6_4_5  (
            .in0(N__13584),
            .in1(N__13703),
            .in2(_gnd_net_),
            .in3(N__13338),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_6_4_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_6_4_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_6_4_6  (
            .in0(N__13702),
            .in1(N__13447),
            .in2(_gnd_net_),
            .in3(N__13608),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26149),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_5_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_5_2 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_6_5_2  (
            .in0(N__13545),
            .in1(N__21852),
            .in2(N__16347),
            .in3(N__13415),
            .lcout(),
            .ltout(\Lab_UT.dispString.m82_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_6_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_6_5_3 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_6_5_3  (
            .in0(N__14757),
            .in1(N__13546),
            .in2(N__13245),
            .in3(N__22052),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_156_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_6_5_4 .LUT_INIT=16'b0011000011111100;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__13687),
            .in2(N__13242),
            .in3(N__13593),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26141),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_4_1_LC_6_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_4_1_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_4_1_LC_6_5_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_4_1_LC_6_5_5  (
            .in0(N__13414),
            .in1(N__13544),
            .in2(N__13700),
            .in3(N__21624),
            .lcout(\Lab_UT.dispString.b1_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_6_6_1 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_6_6_1  (
            .in0(N__13574),
            .in1(N__17850),
            .in2(N__13451),
            .in3(N__21650),
            .lcout(),
            .ltout(\Lab_UT.dispString.m67_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_6_6_2 .LUT_INIT=16'b0100101000001010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_6_6_2  (
            .in0(N__13573),
            .in1(N__22035),
            .in2(N__13620),
            .in3(N__16307),
            .lcout(\Lab_UT.dispString.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_6_3 .LUT_INIT=16'b1100101011001111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_6_6_3  (
            .in0(N__13575),
            .in1(N__13604),
            .in2(N__13452),
            .in3(N__15996),
            .lcout(\Lab_UT.dispString.N_158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_6_6 .LUT_INIT=16'b0010001001011111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_6_6_6  (
            .in0(N__13571),
            .in1(N__21375),
            .in2(N__16500),
            .in3(N__13434),
            .lcout(),
            .ltout(\Lab_UT.dispString.m90_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_6_7 .LUT_INIT=16'b1101001111110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_6_6_7  (
            .in0(N__22034),
            .in1(N__13572),
            .in2(N__13587),
            .in3(N__16471),
            .lcout(\Lab_UT.dispString.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_7_1 .LUT_INIT=16'b1111101100001011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_6_7_1  (
            .in0(N__13568),
            .in1(N__18003),
            .in2(N__13453),
            .in3(N__13344),
            .lcout(\Lab_UT.dispString.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_rep1_LC_6_8_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_LC_6_8_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep1_LC_6_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18151),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26127),
            .ce(N__14243),
            .sr(N__25826));
    defparam \Lab_UT.dictrl.g1_0_3_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_3_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_3_LC_6_9_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \Lab_UT.dictrl.g1_0_3_LC_6_9_0  (
            .in0(N__20487),
            .in1(N__17111),
            .in2(N__13885),
            .in3(N__19439),
            .lcout(Lab_UT_dictrl_g1_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_8_0_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_8_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_8_0_LC_6_9_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_8_0_LC_6_9_1  (
            .in0(N__14006),
            .in1(N__17631),
            .in2(_gnd_net_),
            .in3(N__14369),
            .lcout(\Lab_UT.dictrl.next_state_RNO_8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI6DFS_0_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI6DFS_0_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI6DFS_0_LC_6_9_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI6DFS_0_LC_6_9_2  (
            .in0(N__13954),
            .in1(N__17112),
            .in2(N__13884),
            .in3(N__16600),
            .lcout(\Lab_UT.dictrl.g0_12_a6_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIGV0QF_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIGV0QF_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIGV0QF_LC_6_9_3 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep2_esr_RNIGV0QF_LC_6_9_3  (
            .in0(N__16449),
            .in1(N__13764),
            .in2(N__14844),
            .in3(N__13755),
            .lcout(\Lab_UT.dictrl.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m15_1_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m15_1_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m15_1_LC_6_9_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \Lab_UT.dictrl.m15_1_LC_6_9_4  (
            .in0(N__13955),
            .in1(_gnd_net_),
            .in2(N__13886),
            .in3(N__17113),
            .lcout(\Lab_UT.dictrl.m15Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.m15Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNIMOKF2_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNIMOKF2_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_10_esr_RNIMOKF2_LC_6_9_5 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_esr_RNIMOKF2_LC_6_9_5  (
            .in0(N__15086),
            .in1(N__17630),
            .in2(N__13749),
            .in3(N__14368),
            .lcout(\Lab_UT.dictrl.m27_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_6_10_0 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_1_LC_6_10_0  (
            .in0(N__13746),
            .in1(N__18960),
            .in2(N__13734),
            .in3(N__13710),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_1_LC_6_10_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__23083),
            .in2(N__13737),
            .in3(N__15002),
            .lcout(\Lab_UT.dictrl.next_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26121),
            .ce(N__16884),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_3_1_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_3_1_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_3_1_LC_6_10_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_3_1_LC_6_10_2  (
            .in0(N__24484),
            .in1(N__22750),
            .in2(_gnd_net_),
            .in3(N__24278),
            .lcout(\Lab_UT.dictrl.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_1_1_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_1_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_1_LC_6_10_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_1_LC_6_10_4  (
            .in0(N__18909),
            .in1(N__18150),
            .in2(N__13725),
            .in3(N__24279),
            .lcout(\Lab_UT.dictrl.g0_i_a4_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNISOI03_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNISOI03_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNISOI03_LC_6_11_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep2_esr_RNISOI03_LC_6_11_0  (
            .in0(N__19331),
            .in1(N__24458),
            .in2(N__14013),
            .in3(N__13991),
            .lcout(\Lab_UT.dictrl.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m12_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m12_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m12_LC_6_11_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m12_LC_6_11_1  (
            .in0(N__20498),
            .in1(N__20075),
            .in2(N__18763),
            .in3(N__14350),
            .lcout(\Lab_UT.dictrl.N_88_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_11_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_11_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_11_LC_6_11_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_11_LC_6_11_2  (
            .in0(N__18740),
            .in1(N__20497),
            .in2(N__20091),
            .in3(N__20310),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_9_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_9_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_9_LC_6_11_3 .LUT_INIT=16'b0000000011111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_9_LC_6_11_3  (
            .in0(N__13893),
            .in1(N__14351),
            .in2(N__13974),
            .in3(N__19332),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m53_d_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_6_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_6_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_6_LC_6_11_4 .LUT_INIT=16'b0111001001110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_6_LC_6_11_4  (
            .in0(N__22818),
            .in1(N__24459),
            .in2(N__13971),
            .in3(N__24345),
            .lcout(\Lab_UT.dictrl.N_1102_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_10_0_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_10_0_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_10_0_LC_6_12_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_10_0_LC_6_12_0  (
            .in0(N__18626),
            .in1(N__18920),
            .in2(_gnd_net_),
            .in3(N__24521),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_6_12_1 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_5_0_LC_6_12_1  (
            .in0(N__24522),
            .in1(N__24292),
            .in2(N__13968),
            .in3(N__19366),
            .lcout(\Lab_UT.dictrl.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_10_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_10_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_10_LC_6_12_2 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_10_LC_6_12_2  (
            .in0(N__13875),
            .in1(N__13965),
            .in2(_gnd_net_),
            .in3(N__15624),
            .lcout(\Lab_UT.dictrl.g2_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_9_0_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_9_0_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_9_0_LC_6_12_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_9_0_LC_6_12_3  (
            .in0(N__13876),
            .in1(N__20502),
            .in2(N__13797),
            .in3(N__20297),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m59_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_6_12_4 .LUT_INIT=16'b0101010100111111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_3_0_LC_6_12_4  (
            .in0(N__19367),
            .in1(N__19380),
            .in2(N__14184),
            .in3(N__24524),
            .lcout(\Lab_UT.dictrl.next_state_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_7_0_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_7_0_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_7_0_LC_6_12_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_7_0_LC_6_12_5  (
            .in0(N__24523),
            .in1(_gnd_net_),
            .in2(N__18937),
            .in3(N__18625),
            .lcout(\Lab_UT.dictrl.m63_d_0_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_0_10_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_0_10_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_0_10_LC_6_13_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.g2_0_10_LC_6_13_0  (
            .in0(N__14278),
            .in1(N__14153),
            .in2(N__14121),
            .in3(N__14060),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_4_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2LLA3_LC_6_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2LLA3_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2LLA3_LC_6_13_1 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2LLA3_LC_6_13_1  (
            .in0(N__14181),
            .in1(N__18321),
            .in2(N__14175),
            .in3(N__14329),
            .lcout(\Lab_UT.dictrl.m53_d_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_10_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_10_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_10_LC_6_13_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_10_LC_6_13_2  (
            .in0(N__14279),
            .in1(N__14152),
            .in2(N__14122),
            .in3(N__14059),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_7_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_7_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_7_LC_6_13_3 .LUT_INIT=16'b0101010001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_7_LC_6_13_3  (
            .in0(N__18322),
            .in1(N__14172),
            .in2(N__14166),
            .in3(N__14330),
            .lcout(\Lab_UT.dictrl.m53_d_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_10_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_10_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_10_LC_6_13_4 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_10_LC_6_13_4  (
            .in0(N__14280),
            .in1(N__14151),
            .in2(N__14123),
            .in3(N__14058),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_7_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_7_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_7_LC_6_13_5 .LUT_INIT=16'b0101010001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_7_LC_6_13_5  (
            .in0(N__18323),
            .in1(N__14163),
            .in2(N__14157),
            .in3(N__14331),
            .lcout(\Lab_UT.dictrl.m53_d_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_10_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_10_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_10_LC_6_13_6 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_10_LC_6_13_6  (
            .in0(N__14281),
            .in1(N__14154),
            .in2(N__14124),
            .in3(N__14061),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_7_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_7_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_7_LC_6_13_7 .LUT_INIT=16'b0101010001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_7_LC_6_13_7  (
            .in0(N__18324),
            .in1(N__14382),
            .in2(N__14376),
            .in3(N__14332),
            .lcout(\Lab_UT.dictrl.m53_d_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIMGCH_0_LC_6_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIMGCH_0_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIMGCH_0_LC_6_14_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIMGCH_0_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__16599),
            .in2(_gnd_net_),
            .in3(N__14283),
            .lcout(\Lab_UT.dictrl.N_11_1 ),
            .ltout(\Lab_UT.dictrl.N_11_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_6_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_6_14_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_12_LC_6_14_2  (
            .in0(N__14835),
            .in1(N__15625),
            .in2(N__14295),
            .in3(N__24048),
            .lcout(\Lab_UT.dictrl.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_14_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_14_3  (
            .in0(N__19368),
            .in1(_gnd_net_),
            .in2(N__15700),
            .in3(N__14292),
            .lcout(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOF_LC_6_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOF_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOF_LC_6_14_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOF_LC_6_14_4  (
            .in0(N__18338),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15626),
            .lcout(\Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0 ),
            .ltout(\Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI4DA69_LC_6_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI4DA69_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI4DA69_LC_6_14_5 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNI4DA69_LC_6_14_5  (
            .in0(N__15692),
            .in1(N__24588),
            .in2(N__14286),
            .in3(N__22978),
            .lcout(\Lab_UT.dictrl.N_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_6_LC_6_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_6_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18156),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26117),
            .ce(N__14237),
            .sr(N__25841));
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_6_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_6_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_0_LC_6_15_1  (
            .in0(N__14457),
            .in1(N__22821),
            .in2(_gnd_net_),
            .in3(N__14214),
            .lcout(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_6_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_6_15_2 .LUT_INIT=16'b0011101100011001;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_0_LC_6_15_2  (
            .in0(N__22822),
            .in1(N__24324),
            .in2(N__14205),
            .in3(N__14193),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m67_am_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_6_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_6_15_3 .LUT_INIT=16'b1111000000110101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_0_LC_6_15_3  (
            .in0(N__14514),
            .in1(N__14508),
            .in2(N__14499),
            .in3(N__22823),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_6_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_0_LC_6_15_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_6_15_4  (
            .in0(N__23138),
            .in1(_gnd_net_),
            .in2(N__14496),
            .in3(N__14493),
            .lcout(\Lab_UT.dictrl.next_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26115),
            .ce(N__16899),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_1_2_LC_6_16_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_2_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_2_LC_6_16_3 .LUT_INIT=16'b0011001110100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_2_LC_6_16_3  (
            .in0(N__24321),
            .in1(N__24552),
            .in2(N__14480),
            .in3(N__22824),
            .lcout(\Lab_UT.dictrl.next_state_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI2USJ_1_LC_6_16_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI2USJ_1_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI2USJ_1_LC_6_16_4 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI2USJ_1_LC_6_16_4  (
            .in0(N__15452),
            .in1(N__24040),
            .in2(_gnd_net_),
            .in3(N__15060),
            .lcout(\Lab_UT.dictrl.G_17_i_a5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIVHI53_LC_6_16_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIVHI53_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIVHI53_LC_6_16_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIVHI53_LC_6_16_5  (
            .in0(N__15623),
            .in1(N__19951),
            .in2(N__18604),
            .in3(N__20143),
            .lcout(\Lab_UT.dictrl.N_65 ),
            .ltout(\Lab_UT.dictrl.N_65_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_6_0_LC_6_16_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_6_0_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_6_0_LC_6_16_6 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_6_0_LC_6_16_6  (
            .in0(N__24551),
            .in1(N__15701),
            .in2(N__14460),
            .in3(N__24320),
            .lcout(\Lab_UT.dictrl.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_0  (
            .in0(N__23680),
            .in1(N__23607),
            .in2(N__21049),
            .in3(N__23291),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_1  (
            .in0(N__23608),
            .in1(N__23676),
            .in2(N__20881),
            .in3(N__24957),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_2 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_2  (
            .in0(N__25101),
            .in1(N__14424),
            .in2(N__23693),
            .in3(N__23609),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI90ME1_0_6_LC_7_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI90ME1_0_6_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI90ME1_0_6_LC_7_1_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI90ME1_0_6_LC_7_1_3  (
            .in0(N__23290),
            .in1(N__25100),
            .in2(N__25173),
            .in3(N__24955),
            .lcout(\uu2.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI90ME1_6_LC_7_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI90ME1_6_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI90ME1_6_LC_7_1_4 .LUT_INIT=16'b1101010111111111;
    LogicCell40 \uu2.w_addr_displaying_RNI90ME1_6_LC_7_1_4  (
            .in0(N__24956),
            .in1(N__25167),
            .in2(N__25104),
            .in3(N__23289),
            .lcout(),
            .ltout(\uu2.N_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNIASN45_LC_7_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNIASN45_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNIASN45_LC_7_1_5 .LUT_INIT=16'b0100110100001001;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNIASN45_LC_7_1_5  (
            .in0(N__17322),
            .in1(N__17433),
            .in2(N__14553),
            .in3(N__15732),
            .lcout(\uu2.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIQBDM1_111_LC_7_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIQBDM1_111_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIQBDM1_111_LC_7_2_0 .LUT_INIT=16'b0000000001111011;
    LogicCell40 \uu2.bitmap_RNIQBDM1_111_LC_7_2_0  (
            .in0(N__14696),
            .in1(N__25076),
            .in2(N__14595),
            .in3(N__15720),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_26_i_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI3JIM3_111_LC_7_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI3JIM3_111_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI3JIM3_111_LC_7_2_1 .LUT_INIT=16'b0111110000101100;
    LogicCell40 \uu2.bitmap_RNI3JIM3_111_LC_7_2_1  (
            .in0(N__25077),
            .in1(N__14697),
            .in2(N__14550),
            .in3(N__14607),
            .lcout(),
            .ltout(\uu2.N_55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIE0KH9_111_LC_7_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIE0KH9_111_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIE0KH9_111_LC_7_2_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.bitmap_RNIE0KH9_111_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(N__14547),
            .in2(N__14538),
            .in3(N__20799),
            .lcout(),
            .ltout(\uu2.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIPFVGP_0_LC_7_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIPFVGP_0_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIPFVGP_0_LC_7_2_3 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \uu2.w_addr_displaying_RNIPFVGP_0_LC_7_2_3  (
            .in0(N__14535),
            .in1(N__17664),
            .in2(N__14529),
            .in3(N__15726),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_7_2_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_7_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_7_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_7_3_0 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_296_LC_7_3_0  (
            .in0(N__16533),
            .in1(N__15504),
            .in2(N__16422),
            .in3(N__16376),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_200_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_7_3_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_200_LC_7_3_1  (
            .in0(N__16375),
            .in1(N__16408),
            .in2(N__15514),
            .in3(N__16532),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_72_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_7_3_2 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_72_LC_7_3_2  (
            .in0(N__16535),
            .in1(N__15506),
            .in2(N__16424),
            .in3(N__16378),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_168_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_7_3_3 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_168_LC_7_3_3  (
            .in0(N__16374),
            .in1(N__16407),
            .in2(N__15513),
            .in3(N__16531),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_40_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_7_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_7_3_4 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_40_LC_7_3_4  (
            .in0(N__16534),
            .in1(N__15505),
            .in2(N__16423),
            .in3(N__16377),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_RNIQS1B1_40_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIQS1B1_40_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIQS1B1_40_LC_7_3_5 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.bitmap_RNIQS1B1_40_LC_7_3_5  (
            .in0(N__20673),
            .in1(N__14622),
            .in2(N__14616),
            .in3(N__14733),
            .lcout(\uu2.N_207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNISSSN_162_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNISSSN_162_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNISSSN_162_LC_7_3_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNISSSN_162_LC_7_3_6  (
            .in0(N__14577),
            .in1(N__20672),
            .in2(_gnd_net_),
            .in3(N__14601),
            .lcout(\uu2.N_195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_7_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_7_3_7 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.bitmap_75_LC_7_3_7  (
            .in0(N__16379),
            .in1(N__16418),
            .in2(N__15515),
            .in3(N__16536),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__25768));
    defparam \uu2.bitmap_66_LC_7_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_7_4_2 .LUT_INIT=16'b0000010000111101;
    LogicCell40 \uu2.bitmap_66_LC_7_4_2  (
            .in0(N__15826),
            .in1(N__15964),
            .in2(N__15881),
            .in3(N__15924),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_66C_net ),
            .ce(),
            .sr(N__25766));
    defparam \uu2.bitmap_RNIIGUI_66_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIIGUI_66_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIIGUI_66_LC_7_4_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNIIGUI_66_LC_7_4_3  (
            .in0(N__14583),
            .in1(N__21126),
            .in2(_gnd_net_),
            .in3(N__14646),
            .lcout(\uu2.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_7_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_7_4_4 .LUT_INIT=16'b0000011100111100;
    LogicCell40 \uu2.bitmap_162_LC_7_4_4  (
            .in0(N__15825),
            .in1(N__15963),
            .in2(N__15880),
            .in3(N__15923),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_66C_net ),
            .ce(),
            .sr(N__25766));
    defparam \uu2.bitmap_RNIHL2N_34_LC_7_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIHL2N_34_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIHL2N_34_LC_7_4_6 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \uu2.bitmap_RNIHL2N_34_LC_7_4_6  (
            .in0(N__24889),
            .in1(N__20676),
            .in2(N__14640),
            .in3(N__14628),
            .lcout(\uu2.bitmap_pmux_15_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_69_LC_7_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_7_4_7 .LUT_INIT=16'b0110011100011111;
    LogicCell40 \uu2.bitmap_69_LC_7_4_7  (
            .in0(N__15925),
            .in1(N__15874),
            .in2(N__15971),
            .in3(N__15827),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_66C_net ),
            .ce(),
            .sr(N__25766));
    defparam \uu2.bitmap_111_LC_7_5_0 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_7_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_7_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14726),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \uu2.vram_rd_clk_det_0_LC_7_5_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_7_5_1 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_7_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14685),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \uu2.vram_rd_clk_det_1_LC_7_5_2 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_7_5_2 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_7_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16023),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \uu2.bitmap_194_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_7_5_4 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_194_LC_7_5_4  (
            .in0(N__15960),
            .in1(N__15918),
            .in2(N__15878),
            .in3(N__15822),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \uu2.bitmap_34_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_7_5_6 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_34_LC_7_5_6  (
            .in0(N__15962),
            .in1(N__15922),
            .in2(N__15879),
            .in3(N__15824),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \uu2.bitmap_290_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_7_5_7 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_290_LC_7_5_7  (
            .in0(N__15823),
            .in1(N__15864),
            .in2(N__15929),
            .in3(N__15961),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_111C_net ),
            .ce(),
            .sr(N__25765));
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_7_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_0_LC_7_6_0  (
            .in0(N__21774),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26146),
            .ce(N__14775),
            .sr(N__25804));
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_1_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25521),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26146),
            .ce(N__14775),
            .sr(N__25804));
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_7_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_2_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26723),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26146),
            .ce(N__14775),
            .sr(N__25804));
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_7_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_3_LC_7_6_3  (
            .in0(N__26421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26146),
            .ce(N__14775),
            .sr(N__25804));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_7_0 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_7_0  (
            .in0(N__18411),
            .in1(N__26420),
            .in2(N__14742),
            .in3(N__22213),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_7_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_7_7_1  (
            .in0(N__22178),
            .in1(N__22209),
            .in2(N__14760),
            .in3(N__18372),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26138),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_1_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_1_LC_7_7_2 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.dispString.m49_1_LC_7_7_2  (
            .in0(N__26231),
            .in1(N__21847),
            .in2(N__22214),
            .in3(N__14755),
            .lcout(\Lab_UT.dispString.m49Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNITK144_3_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNITK144_3_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNITK144_3_LC_7_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNITK144_3_LC_7_7_3  (
            .in0(N__14756),
            .in1(N__22208),
            .in2(_gnd_net_),
            .in3(N__21344),
            .lcout(\Lab_UT.min1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNIR6J44_3_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIR6J44_3_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIR6J44_3_LC_7_7_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNIR6J44_3_LC_7_7_4  (
            .in0(N__21343),
            .in1(_gnd_net_),
            .in2(N__26235),
            .in3(N__21848),
            .lcout(\Lab_UT.min2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_7_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_7_5  (
            .in0(N__21914),
            .in1(N__22281),
            .in2(_gnd_net_),
            .in3(N__21971),
            .lcout(\Lab_UT.didp.countrce4.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_LC_7_8_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_LC_7_8_0  (
            .in0(N__22425),
            .in1(N__22380),
            .in2(N__22467),
            .in3(N__22968),
            .lcout(\Lab_UT.dictrl.state_1_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26132),
            .ce(N__22487),
            .sr(N__25799));
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNI3AA01_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNI3AA01_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNI3AA01_LC_7_8_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep2_esr_RNI3AA01_LC_7_8_1  (
            .in0(N__19779),
            .in1(_gnd_net_),
            .in2(N__19330),
            .in3(N__23084),
            .lcout(\Lab_UT.dictrl.g0_12_a6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_4_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_4_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_4_LC_7_8_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_4_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__19317),
            .in2(_gnd_net_),
            .in3(N__19778),
            .lcout(\Lab_UT.dictrl.g2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNINE144_0_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNINE144_0_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNINE144_0_LC_7_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNINE144_0_LC_7_8_3  (
            .in0(N__16475),
            .in1(N__21301),
            .in2(_gnd_net_),
            .in3(N__21970),
            .lcout(\Lab_UT.min1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPG144_1_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPG144_1_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPG144_1_LC_7_8_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIPG144_1_LC_7_8_4  (
            .in0(N__21302),
            .in1(N__22279),
            .in2(_gnd_net_),
            .in3(N__16282),
            .lcout(\Lab_UT.min1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRI144_2_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRI144_2_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIRI144_2_LC_7_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIRI144_2_LC_7_8_5  (
            .in0(N__21326),
            .in1(N__21907),
            .in2(_gnd_net_),
            .in3(N__16308),
            .lcout(\Lab_UT.min1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI56JGE_1_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI56JGE_1_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI56JGE_1_LC_7_9_0 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI56JGE_1_LC_7_9_0  (
            .in0(N__15044),
            .in1(N__24032),
            .in2(N__23163),
            .in3(N__15248),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_7_9_1 .LUT_INIT=16'b1110000011110001;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_2_LC_7_9_1  (
            .in0(N__24034),
            .in1(N__23152),
            .in2(N__15258),
            .in3(N__15048),
            .lcout(\Lab_UT.dictrl.state_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_7_9_2 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_LC_7_9_2  (
            .in0(N__15045),
            .in1(N__24037),
            .in2(N__23164),
            .in3(N__15249),
            .lcout(\Lab_UT.dictrl.state_2_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_LC_7_9_3 .LUT_INIT=16'b1110000011110001;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep2_esr_LC_7_9_3  (
            .in0(N__24033),
            .in1(N__23148),
            .in2(N__15257),
            .in3(N__15046),
            .lcout(\Lab_UT.dictrl.state_2_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_7_9_4 .LUT_INIT=16'b1111110100000001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_2_LC_7_9_4  (
            .in0(N__15047),
            .in1(N__24038),
            .in2(N__23165),
            .in3(N__15253),
            .lcout(\Lab_UT.dictrl.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_7_9_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_7_9_5 .LUT_INIT=16'b0000111000011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_LC_7_9_5  (
            .in0(N__24035),
            .in1(N__23153),
            .in2(N__15021),
            .in3(N__15006),
            .lcout(\Lab_UT.dictrl.state_i_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI7ECM_LC_7_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI7ECM_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI7ECM_LC_7_9_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNI7ECM_LC_7_9_6  (
            .in0(N__18199),
            .in1(N__19767),
            .in2(N__14985),
            .in3(N__19617),
            .lcout(\Lab_UT.LdASones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_7_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_7_9_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_7_9_7 .LUT_INIT=16'b0001111100001110;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_LC_7_9_7  (
            .in0(N__24036),
            .in1(N__23154),
            .in2(N__15168),
            .in3(N__14976),
            .lcout(\Lab_UT.state_i_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26129),
            .ce(N__22488),
            .sr(N__25802));
    defparam \Lab_UT.dictrl.state_ret_12_RNIRIHQ6_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNIRIHQ6_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNIRIHQ6_LC_7_10_0 .LUT_INIT=16'b0011101100111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNIRIHQ6_LC_7_10_0  (
            .in0(N__15151),
            .in1(N__16978),
            .in2(N__24049),
            .in3(N__15130),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNI2MD42_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNI2MD42_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNI2MD42_LC_7_10_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNI2MD42_LC_7_10_1  (
            .in0(N__25874),
            .in1(N__14964),
            .in2(N__24052),
            .in3(N__14898),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNIROSR8_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNIROSR8_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNIROSR8_LC_7_10_2 .LUT_INIT=16'b1011000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNIROSR8_LC_7_10_2  (
            .in0(N__15152),
            .in1(N__16979),
            .in2(N__14856),
            .in3(N__15131),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI71KU22_1_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI71KU22_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI71KU22_1_LC_7_10_3 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI71KU22_1_LC_7_10_3  (
            .in0(N__22587),
            .in1(N__14853),
            .in2(N__14847),
            .in3(N__23191),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_10_4 .LUT_INIT=16'b0011101100111000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_10_4  (
            .in0(N__15156),
            .in1(N__16987),
            .in2(N__24051),
            .in3(N__15133),
            .lcout(\Lab_UT.dictrl.state_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26125),
            .ce(N__22490),
            .sr(N__25803));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_10_5 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_10_5  (
            .in0(N__23997),
            .in1(N__15153),
            .in2(N__16988),
            .in3(N__15134),
            .lcout(\Lab_UT.dictrl.state_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26125),
            .ce(N__22490),
            .sr(N__25803));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_10_6 .LUT_INIT=16'b0011101100111000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_10_6  (
            .in0(N__15154),
            .in1(N__16983),
            .in2(N__24050),
            .in3(N__15132),
            .lcout(\Lab_UT.dictrl.state_3_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26125),
            .ce(N__22490),
            .sr(N__25803));
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_7_10_7 .LUT_INIT=16'b0100111101001010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_3_LC_7_10_7  (
            .in0(N__23998),
            .in1(N__15155),
            .in2(N__16989),
            .in3(N__15135),
            .lcout(\Lab_UT.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26125),
            .ce(N__22490),
            .sr(N__25803));
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_11_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_11_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_LC_7_11_0  (
            .in0(N__15068),
            .in1(N__15182),
            .in2(_gnd_net_),
            .in3(N__15665),
            .lcout(\Lab_UT.dictrl.state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26123),
            .ce(N__22491),
            .sr(N__25807));
    defparam \Lab_UT.dictrl.state_0_esr_RNIS4PO5_2_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIS4PO5_2_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIS4PO5_2_LC_7_11_1 .LUT_INIT=16'b1000110111011101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIS4PO5_2_LC_7_11_1  (
            .in0(N__22775),
            .in1(N__15108),
            .in2(N__16440),
            .in3(N__24144),
            .lcout(\Lab_UT.dictrl.N_62 ),
            .ltout(\Lab_UT.dictrl.N_62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_11_2 .LUT_INIT=16'b1011000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_esr_LC_7_11_2  (
            .in0(N__15069),
            .in1(N__15183),
            .in2(N__15099),
            .in3(N__22551),
            .lcout(\Lab_UT.dictrl.N_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26123),
            .ce(N__22491),
            .sr(N__25807));
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_1_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_1_LC_7_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIP2CG_1_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__23082),
            .in2(_gnd_net_),
            .in3(N__23911),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_11_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_1_LC_7_11_4  (
            .in0(N__22420),
            .in1(N__22372),
            .in2(N__22463),
            .in3(N__22945),
            .lcout(\Lab_UT.dictrl.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26123),
            .ce(N__22491),
            .sr(N__25807));
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_11_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_11_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_11_5  (
            .in0(N__22943),
            .in1(N__22421),
            .in2(N__22379),
            .in3(N__22458),
            .lcout(\Lab_UT.dictrl.state_fast_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26123),
            .ce(N__22491),
            .sr(N__25807));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_11_6 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_11_6  (
            .in0(N__22419),
            .in1(N__22371),
            .in2(N__22462),
            .in3(N__22944),
            .lcout(\Lab_UT.dictrl.state_1_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26123),
            .ce(N__22491),
            .sr(N__25807));
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ2M68_3_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ2M68_3_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ2M68_3_LC_7_12_0 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIQ2M68_3_LC_7_12_0  (
            .in0(N__15267),
            .in1(N__15231),
            .in2(N__24533),
            .in3(N__15200),
            .lcout(\Lab_UT.dictrl.N_1459_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_71_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_71_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_71_LC_7_12_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.g0_71_LC_7_12_1  (
            .in0(N__18935),
            .in1(N__20597),
            .in2(N__19193),
            .in3(N__20196),
            .lcout(\Lab_UT.dictrl.N_40_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.g0_35_LC_7_12_2  (
            .in0(N__20197),
            .in1(N__19164),
            .in2(N__20601),
            .in3(N__18936),
            .lcout(\Lab_UT.dictrl.N_40_3 ),
            .ltout(\Lab_UT.dictrl.N_40_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_7_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_7_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_7_LC_7_12_3 .LUT_INIT=16'b1000100010001101;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_7_LC_7_12_3  (
            .in0(N__24030),
            .in1(N__19532),
            .in2(N__15225),
            .in3(N__24489),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1462_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_2_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_2_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_2_LC_7_12_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_2_LC_7_12_4  (
            .in0(N__15222),
            .in1(N__15216),
            .in2(N__15207),
            .in3(N__24031),
            .lcout(\Lab_UT.dictrl.N_1460_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI78VA1_1_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI78VA1_1_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI78VA1_1_LC_7_13_0 .LUT_INIT=16'b0000100000001111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI78VA1_1_LC_7_13_0  (
            .in0(N__24304),
            .in1(N__22777),
            .in2(N__24058),
            .in3(N__23119),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNITVS29_3_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNITVS29_3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNITVS29_3_LC_7_13_1 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNITVS29_3_LC_7_13_1  (
            .in0(N__15204),
            .in1(N__15693),
            .in2(N__15186),
            .in3(N__24491),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_7_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_7_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_7_LC_7_13_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_7_LC_7_13_2  (
            .in0(N__24303),
            .in1(N__19959),
            .in2(N__24057),
            .in3(N__22776),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_1_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_1_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_1_LC_7_13_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_1_LC_7_13_3  (
            .in0(N__15441),
            .in1(N__17250),
            .in2(N__15171),
            .in3(N__17292),
            .lcout(\Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_5_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_5_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_5_LC_7_13_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_5_LC_7_13_4  (
            .in0(N__24490),
            .in1(N__15456),
            .in2(_gnd_net_),
            .in3(N__24017),
            .lcout(\Lab_UT.dictrl.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m23_0_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m23_0_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m23_0_LC_7_14_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.m23_0_LC_7_14_0  (
            .in0(N__20159),
            .in1(N__20580),
            .in2(N__20094),
            .in3(N__20325),
            .lcout(\Lab_UT.dictrl.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_7_14_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_15_LC_7_14_1  (
            .in0(N__15399),
            .in1(N__15364),
            .in2(N__15340),
            .in3(N__23963),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_7_14_2 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_11_LC_7_14_2  (
            .in0(N__20157),
            .in1(N__20578),
            .in2(N__15435),
            .in3(N__20323),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_18_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_7_14_3 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_4_LC_7_14_3  (
            .in0(N__15543),
            .in1(N__15432),
            .in2(N__15426),
            .in3(N__23964),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_18_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_18_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_18_LC_7_14_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.g0_18_LC_7_14_4  (
            .in0(N__20158),
            .in1(N__20579),
            .in2(N__18605),
            .in3(N__20324),
            .lcout(\Lab_UT.dictrl.N_40_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_7_14_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_14_LC_7_14_5  (
            .in0(N__15400),
            .in1(N__15365),
            .in2(N__15341),
            .in3(N__23962),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_a7_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_15_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_15_0  (
            .in0(N__15309),
            .in1(N__20215),
            .in2(N__15303),
            .in3(N__19952),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_22_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_7_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_7_15_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_3_LC_7_15_1  (
            .in0(N__20232),
            .in1(N__15294),
            .in2(N__15282),
            .in3(N__15279),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_8_LC_7_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_8_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_8_LC_7_15_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_8_LC_7_15_2  (
            .in0(N__20031),
            .in1(N__20214),
            .in2(_gnd_net_),
            .in3(N__19953),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_97_mux_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_5_LC_7_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_5_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_5_LC_7_15_3 .LUT_INIT=16'b0010001011101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_5_LC_7_15_3  (
            .in0(N__15714),
            .in1(N__19844),
            .in2(N__15705),
            .in3(N__19725),
            .lcout(\Lab_UT.dictrl.N_1102_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_2_LC_7_16_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_2_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_2_LC_7_16_0 .LUT_INIT=16'b0001000000011111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_2_LC_7_16_0  (
            .in0(N__24534),
            .in1(N__15702),
            .in2(N__23166),
            .in3(N__15666),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_2_LC_7_16_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_2_LC_7_16_1 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_7_16_1  (
            .in0(N__15642),
            .in1(N__23159),
            .in2(N__15651),
            .in3(N__15648),
            .lcout(\Lab_UT.dictrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26116),
            .ce(N__16895),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_7_16_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_7_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_2_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__22801),
            .in2(_gnd_net_),
            .in3(N__24322),
            .lcout(\Lab_UT.dictrl.next_state_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNINV3P_2_LC_7_16_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNINV3P_2_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNINV3P_2_LC_7_16_5 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNINV3P_2_LC_7_16_5  (
            .in0(N__15607),
            .in1(N__15539),
            .in2(_gnd_net_),
            .in3(N__24041),
            .lcout(\Lab_UT.dictrl.next_state_RNINV3PZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_203_LC_8_1_0 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_8_1_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_203_LC_8_1_0  (
            .in0(N__16383),
            .in1(N__16425),
            .in2(N__15516),
            .in3(N__16530),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__25774));
    defparam \uu2.bitmap_RNIPJHV_200_LC_8_1_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPJHV_200_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPJHV_200_LC_8_1_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNIPJHV_200_LC_8_1_1  (
            .in0(N__15471),
            .in1(N__17797),
            .in2(_gnd_net_),
            .in3(N__15465),
            .lcout(\uu2.N_199 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_8_1_2 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_8_1_2  (
            .in0(N__17800),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25020),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_203C_net ),
            .ce(),
            .sr(N__25774));
    defparam \uu2.w_addr_displaying_0_rep1_RNIDASJ_LC_8_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNIDASJ_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNIDASJ_LC_8_1_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNIDASJ_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__20742),
            .in2(_gnd_net_),
            .in3(N__17798),
            .lcout(\uu2.w_addr_displaying_0_rep1_RNIDASJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_rep1_RNI8NUT1_LC_8_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNI8NUT1_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNI8NUT1_LC_8_1_4 .LUT_INIT=16'b1000000000000100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNI8NUT1_LC_8_1_4  (
            .in0(N__17799),
            .in1(N__17565),
            .in2(N__17382),
            .in3(N__20754),
            .lcout(\uu2.bitmap_pmux_sn_N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIBTRT7_0_LC_8_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIBTRT7_0_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIBTRT7_0_LC_8_2_0 .LUT_INIT=16'b0110000011111001;
    LogicCell40 \uu2.w_addr_displaying_RNIBTRT7_0_LC_8_2_0  (
            .in0(N__23328),
            .in1(N__23462),
            .in2(N__17751),
            .in3(N__17586),
            .lcout(\uu2.N_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIBP86_2_LC_8_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIBP86_2_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIBP86_2_LC_8_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIBP86_2_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__20628),
            .in2(_gnd_net_),
            .in3(N__20661),
            .lcout(\uu2.N_24_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_LC_8_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_8_2_2 .LUT_INIT=16'b1100110001100110;
    LogicCell40 \uu2.w_addr_displaying_1_LC_8_2_2  (
            .in0(N__23330),
            .in1(N__23464),
            .in2(_gnd_net_),
            .in3(N__24999),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__25771));
    defparam \uu2.w_addr_displaying_fast_2_LC_8_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_8_2_3 .LUT_INIT=16'b1011111101000000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_8_2_3  (
            .in0(N__25001),
            .in1(N__23334),
            .in2(N__23485),
            .in3(N__20629),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__25771));
    defparam \uu2.w_addr_displaying_fast_1_LC_8_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_1_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_1_LC_8_2_4 .LUT_INIT=16'b1010101001011010;
    LogicCell40 \uu2.w_addr_displaying_fast_1_LC_8_2_4  (
            .in0(N__20784),
            .in1(_gnd_net_),
            .in2(N__23343),
            .in3(N__25000),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__25771));
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_8_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_8_2_5 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_8_2_5  (
            .in0(N__20633),
            .in1(N__20662),
            .in2(_gnd_net_),
            .in3(N__20783),
            .lcout(\uu2.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIU1AF7_0_LC_8_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIU1AF7_0_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIU1AF7_0_LC_8_2_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.w_addr_displaying_RNIU1AF7_0_LC_8_2_6  (
            .in0(N__23329),
            .in1(N__23463),
            .in2(_gnd_net_),
            .in3(N__24998),
            .lcout(\uu2.w_addr_displaying_RNIU1AF7Z0Z_0 ),
            .ltout(\uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_3_LC_8_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_3_LC_8_2_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.w_addr_displaying_fast_3_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__17654),
            .in2(N__15975),
            .in3(N__20663),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1C_net ),
            .ce(),
            .sr(N__25771));
    defparam \uu2.bitmap_197_LC_8_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_8_3_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_197_LC_8_3_0  (
            .in0(N__15972),
            .in1(N__15930),
            .in2(N__15885),
            .in3(N__15831),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__25769));
    defparam \uu2.bitmap_RNIOMUI_69_LC_8_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIOMUI_69_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIOMUI_69_LC_8_3_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNIOMUI_69_LC_8_3_1  (
            .in0(N__15789),
            .in1(N__21127),
            .in2(_gnd_net_),
            .in3(N__15783),
            .lcout(\uu2.N_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_7_LC_8_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_3_2 .LUT_INIT=16'b0100110001100110;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_8_3_2  (
            .in0(N__23252),
            .in1(N__21132),
            .in2(N__25162),
            .in3(N__15772),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__25769));
    defparam \uu2.w_addr_displaying_7_LC_8_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_8_3_3 .LUT_INIT=16'b0010101001100110;
    LogicCell40 \uu2.w_addr_displaying_7_LC_8_3_3  (
            .in0(N__25088),
            .in1(N__23250),
            .in2(N__25169),
            .in3(N__15769),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__25769));
    defparam \uu2.w_addr_displaying_8_LC_8_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_8_3_4 .LUT_INIT=16'b0101001011110000;
    LogicCell40 \uu2.w_addr_displaying_8_LC_8_3_4  (
            .in0(N__23251),
            .in1(N__15770),
            .in2(N__25163),
            .in3(N__25089),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__25769));
    defparam \uu2.w_addr_displaying_RNIHDHP6_8_LC_8_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIHDHP6_8_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIHDHP6_8_LC_8_3_5 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \uu2.w_addr_displaying_RNIHDHP6_8_LC_8_3_5  (
            .in0(N__25087),
            .in1(N__23249),
            .in2(N__25168),
            .in3(N__15768),
            .lcout(\uu2.w_addr_displaying_RNIHDHP6Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_8_LC_8_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_8_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_8_LC_8_3_6 .LUT_INIT=16'b0101111100100000;
    LogicCell40 \uu2.w_addr_displaying_fast_8_LC_8_3_6  (
            .in0(N__25079),
            .in1(N__15771),
            .in2(N__23256),
            .in3(N__24890),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__25769));
    defparam \uu2.w_addr_displaying_RNIR2PL_8_LC_8_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIR2PL_8_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIR2PL_8_LC_8_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_RNIR2PL_8_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__25078),
            .in2(_gnd_net_),
            .in3(N__25136),
            .lcout(\uu2.w_addr_displaying_RNIR2PLZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_2_LC_8_4_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_8_4_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_8_4_0 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_8_4_0  (
            .in0(N__16254),
            .in1(N__16191),
            .in2(N__16152),
            .in3(N__16103),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26170),
            .ce(N__16089),
            .sr(N__25842));
    defparam \uu2.bitmap_RNI71NJ_72_LC_8_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI71NJ_72_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI71NJ_72_LC_8_4_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNI71NJ_72_LC_8_4_1  (
            .in0(N__17801),
            .in1(N__16044),
            .in2(_gnd_net_),
            .in3(N__16038),
            .lcout(\uu2.N_196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_8_4_2 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_8_4_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_8_4_2  (
            .in0(N__16032),
            .in1(N__16022),
            .in2(_gnd_net_),
            .in3(N__25873),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_0_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_0_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_0_LC_8_5_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.dispString.m49_0_LC_8_5_0  (
            .in0(N__25222),
            .in1(N__16336),
            .in2(N__17715),
            .in3(N__15988),
            .lcout(\Lab_UT.dispString.m49Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNINAM54_3_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNINAM54_3_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNINAM54_3_LC_8_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNINAM54_3_LC_8_5_1  (
            .in0(N__15989),
            .in1(N__21340),
            .in2(_gnd_net_),
            .in3(N__17711),
            .lcout(\Lab_UT.sec2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNIPO4L3_3_LC_8_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIPO4L3_3_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIPO4L3_3_LC_8_5_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNIPO4L3_3_LC_8_5_2  (
            .in0(N__21341),
            .in1(_gnd_net_),
            .in2(N__25227),
            .in3(N__16337),
            .lcout(\Lab_UT.sec1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_8_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_8_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_3_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26413),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26161),
            .ce(N__18021),
            .sr(N__25813));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJ6M54_1_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJ6M54_1_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJ6M54_1_LC_8_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIJ6M54_1_LC_8_5_4  (
            .in0(N__21336),
            .in1(N__21255),
            .in2(_gnd_net_),
            .in3(N__21190),
            .lcout(\Lab_UT.sec2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_8_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_1_LC_8_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25523),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26161),
            .ce(N__18021),
            .sr(N__25813));
    defparam \Lab_UT.didp.regrce3.q_esr_RNIN2J44_1_LC_8_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIN2J44_1_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIN2J44_1_LC_8_5_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNIN2J44_1_LC_8_5_6  (
            .in0(N__21620),
            .in1(_gnd_net_),
            .in2(N__21348),
            .in3(N__26577),
            .lcout(\Lab_UT.min2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNIP4J44_2_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIP4J44_2_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIP4J44_2_LC_8_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNIP4J44_2_LC_8_5_7  (
            .in0(N__21342),
            .in1(N__26499),
            .in2(_gnd_net_),
            .in3(N__21651),
            .lcout(\Lab_UT.min2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_8_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_1_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25522),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26153),
            .ce(N__16323),
            .sr(N__25809));
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_8_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_2_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26724),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26153),
            .ce(N__16323),
            .sr(N__25809));
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_8_6_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_3_LC_8_6_2  (
            .in0(N__26422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26153),
            .ce(N__16323),
            .sr(N__25809));
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_8_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_0_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21775),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26153),
            .ce(N__16323),
            .sr(N__25809));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_8_7_0 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_8_7_0  (
            .in0(N__18407),
            .in1(N__26715),
            .in2(N__16677),
            .in3(N__21905),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_7_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_8_7_1  (
            .in0(N__21906),
            .in1(N__22177),
            .in2(N__16311),
            .in3(N__18371),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26147),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_3_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_3_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_3_LC_8_7_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dispString.m49_3_LC_8_7_2  (
            .in0(N__16303),
            .in1(N__22269),
            .in2(N__16286),
            .in3(N__21904),
            .lcout(),
            .ltout(\Lab_UT.dispString.m49Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_12_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_12_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_12_LC_8_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dispString.m49_12_LC_8_7_3  (
            .in0(N__16557),
            .in1(N__16548),
            .in2(N__16542),
            .in3(N__21588),
            .lcout(\Lab_UT.dispString.m49Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_8_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_0_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21805),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26139),
            .ce(N__21821),
            .sr(N__25801));
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_8_8_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_8_8_1  (
            .in0(N__16644),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25878),
            .lcout(\Lab_UT.didp.regrce3.LdAMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNILRDD3_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNILRDD3_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNILRDD3_LC_8_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNILRDD3_LC_8_8_2  (
            .in0(N__18032),
            .in1(N__16655),
            .in2(N__16628),
            .in3(N__16643),
            .lcout(\Lab_UT.loadalarm_0 ),
            .ltout(\Lab_UT.loadalarm_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNIL0J44_0_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIL0J44_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNIL0J44_0_LC_8_8_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNIL0J44_0_LC_8_8_3  (
            .in0(N__26538),
            .in1(N__16490),
            .in2(N__16539),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.min2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_7_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_7_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_7_LC_8_8_4 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.dispString.m49_7_LC_8_8_4  (
            .in0(N__16489),
            .in1(N__26537),
            .in2(N__16476),
            .in3(N__21948),
            .lcout(\Lab_UT.dispString.m49Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIAOPO_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIAOPO_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIAOPO_LC_8_9_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNIAOPO_LC_8_9_0  (
            .in0(N__22948),
            .in1(N__18287),
            .in2(N__19048),
            .in3(N__16797),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_12_a6_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIK3DC4_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIK3DC4_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIK3DC4_LC_8_9_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNIK3DC4_LC_8_9_1  (
            .in0(N__18155),
            .in1(N__19198),
            .in2(N__16452),
            .in3(N__18780),
            .lcout(\Lab_UT.dictrl.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_14_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_14_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_14_LC_8_9_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_14_LC_8_9_2  (
            .in0(N__19040),
            .in1(_gnd_net_),
            .in2(N__19210),
            .in3(N__18153),
            .lcout(\Lab_UT.dictrl.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIG5AU_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIG5AU_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIG5AU_LC_8_9_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNIG5AU_LC_8_9_3  (
            .in0(N__18154),
            .in1(N__19041),
            .in2(N__18224),
            .in3(N__19197),
            .lcout(\Lab_UT.dictrl.m35_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__22266),
            .in2(_gnd_net_),
            .in3(N__21952),
            .lcout(\Lab_UT.didp.countrce4.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNI9E421_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNI9E421_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNI9E421_LC_8_9_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNI9E421_LC_8_9_5  (
            .in0(N__19615),
            .in1(N__18170),
            .in2(_gnd_net_),
            .in3(N__19271),
            .lcout(\Lab_UT.LdAMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI79EL_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI79EL_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI79EL_LC_8_9_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNI79EL_LC_8_9_6  (
            .in0(N__22947),
            .in1(N__19616),
            .in2(N__18217),
            .in3(N__16795),
            .lcout(\Lab_UT.LdAMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIULEV_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIULEV_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIULEV_LC_8_9_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNIULEV_LC_8_9_7  (
            .in0(N__16796),
            .in1(N__22946),
            .in2(N__19310),
            .in3(N__19618),
            .lcout(\Lab_UT.LdAStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_LC_8_10_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_ess_LC_8_10_0 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_LC_8_10_0  (
            .in0(N__16611),
            .in1(N__22878),
            .in2(N__17229),
            .in3(N__22588),
            .lcout(\Lab_UT.dicRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_10_1 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_10_1  (
            .in0(N__17016),
            .in1(N__16860),
            .in2(N__17046),
            .in3(N__17148),
            .lcout(\Lab_UT.dictrl.state_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_10_2 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_10_2  (
            .in0(N__17145),
            .in1(N__17037),
            .in2(N__16862),
            .in3(N__17013),
            .lcout(\Lab_UT.dictrl.state_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_LC_8_10_3 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep2_esr_LC_8_10_3  (
            .in0(N__17014),
            .in1(N__16856),
            .in2(N__17045),
            .in3(N__17146),
            .lcout(\Lab_UT.dictrl.state_0_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_10_4 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_0_LC_8_10_4  (
            .in0(N__17147),
            .in1(N__17041),
            .in2(N__16863),
            .in3(N__17015),
            .lcout(\Lab_UT.dictrl.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIN23OR_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIN23OR_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNIN23OR_LC_8_10_6 .LUT_INIT=16'b0000000000010011;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNIN23OR_LC_8_10_6  (
            .in0(N__17144),
            .in1(N__17036),
            .in2(N__16861),
            .in3(N__17012),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_0 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_10_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_10_7 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_LC_8_10_7  (
            .in0(N__22589),
            .in1(N__22552),
            .in2(N__16992),
            .in3(N__17214),
            .lcout(\Lab_UT.LdStens_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26130),
            .ce(N__22489),
            .sr(N__25808));
    defparam \Lab_UT.dictrl.next_state_RNICLDV_3_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNICLDV_3_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNICLDV_3_LC_8_11_0 .LUT_INIT=16'b0001101100001010;
    LogicCell40 \Lab_UT.dictrl.next_state_RNICLDV_3_LC_8_11_0  (
            .in0(N__23905),
            .in1(N__19305),
            .in2(N__16908),
            .in3(N__16834),
            .lcout(\Lab_UT.dictrl.next_state_latmux_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_8_11_1  (
            .in0(N__16955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26126),
            .ce(N__16894),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI4JJN_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI4JJN_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_RNI4JJN_LC_8_11_2 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_RNI4JJN_LC_8_11_2  (
            .in0(N__19850),
            .in1(N__19306),
            .in2(N__24012),
            .in3(N__16836),
            .lcout(\Lab_UT.dictrl.G_17_i_a5_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_8_11_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_5_LC_8_11_3  (
            .in0(N__16835),
            .in1(N__19851),
            .in2(N__19329),
            .in3(N__23909),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_8_11_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_2_LC_8_11_4  (
            .in0(N__16770),
            .in1(N__16761),
            .in2(N__16749),
            .in3(N__16746),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_8_11_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_1_LC_8_11_5  (
            .in0(N__25926),
            .in1(N__16733),
            .in2(N__16737),
            .in3(N__22550),
            .lcout(\Lab_UT.dictrl.state_ret_12and_0_ns_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_8_11_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_0_LC_8_11_6  (
            .in0(N__23910),
            .in1(N__25925),
            .in2(N__22560),
            .in3(N__16734),
            .lcout(\Lab_UT.dictrl.state_ret_12and_0_ns_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI6TSE1_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI6TSE1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNI6TSE1_LC_8_12_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_RNI6TSE1_LC_8_12_0  (
            .in0(N__25494),
            .in1(N__26687),
            .in2(_gnd_net_),
            .in3(N__17205),
            .lcout(\Lab_UT.dictrl.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_7_1_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_7_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_7_1_LC_8_12_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_7_1_LC_8_12_1  (
            .in0(N__26688),
            .in1(N__18927),
            .in2(N__26391),
            .in3(N__25497),
            .lcout(\Lab_UT.dictrl.g0_i_a4_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_16_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_16_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_16_LC_8_12_2 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_16_LC_8_12_2  (
            .in0(N__25496),
            .in1(N__26370),
            .in2(N__18938),
            .in3(N__26689),
            .lcout(\Lab_UT.dictrl.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_i_m2_5_N_3L3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_i_m2_5_N_3L3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_i_m2_5_N_3L3_LC_8_12_3 .LUT_INIT=16'b0001111100000000;
    LogicCell40 \Lab_UT.dictrl.g0_i_m2_5_N_3L3_LC_8_12_3  (
            .in0(N__26686),
            .in1(N__25495),
            .in2(N__26390),
            .in3(N__17107),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3_3_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3_3_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3_3_LC_8_12_4 .LUT_INIT=16'b0100011101110111;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3_3_LC_8_12_4  (
            .in0(N__18243),
            .in1(N__17165),
            .in2(N__17181),
            .in3(N__17178),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNII5BFA_2_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNII5BFA_2_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNII5BFA_2_LC_8_12_5 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNII5BFA_2_LC_8_12_5  (
            .in0(N__17166),
            .in1(N__17244),
            .in2(N__17151),
            .in3(N__17052),
            .lcout(\Lab_UT.dictrl.N_1792_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIQV2R6_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIQV2R6_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNIQV2R6_LC_8_13_0 .LUT_INIT=16'b0100010011101111;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep2_esr_RNIQV2R6_LC_8_13_0  (
            .in0(N__19830),
            .in1(N__17127),
            .in2(N__18432),
            .in3(N__19700),
            .lcout(\Lab_UT.dictrl.N_1102_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_16_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_16_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_16_LC_8_13_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_16_LC_8_13_1  (
            .in0(N__20595),
            .in1(N__17118),
            .in2(N__18606),
            .in3(N__20217),
            .lcout(\Lab_UT.dictrl.N_40_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_13_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_13_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_13_LC_8_13_3 .LUT_INIT=16'b0011000100010001;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_13_LC_8_13_3  (
            .in0(N__19315),
            .in1(N__24016),
            .in2(N__18939),
            .in3(N__19831),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_4_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_4_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_4_LC_8_13_4 .LUT_INIT=16'b0001000010100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_4_LC_8_13_4  (
            .in0(N__17262),
            .in1(N__20596),
            .in2(N__17253),
            .in3(N__19316),
            .lcout(\Lab_UT.dictrl.g0_i_m2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_17_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_LC_8_13_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_17_LC_8_13_5  (
            .in0(N__18602),
            .in1(N__20218),
            .in2(_gnd_net_),
            .in3(N__19958),
            .lcout(\Lab_UT.dictrl.N_97_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_8_14_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_8_14_0  (
            .in0(N__24271),
            .in1(N__20205),
            .in2(N__19211),
            .in3(N__23981),
            .lcout(\Lab_UT.dictrl.g0_i_a5_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_36_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_36_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_36_LC_8_14_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dictrl.g0_36_LC_8_14_1  (
            .in0(N__19956),
            .in1(_gnd_net_),
            .in2(N__20221),
            .in3(N__19199),
            .lcout(\Lab_UT.dictrl.N_97_mux_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_65_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_65_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_65_LC_8_14_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_65_LC_8_14_2  (
            .in0(N__20077),
            .in1(N__20198),
            .in2(_gnd_net_),
            .in3(N__19954),
            .lcout(\Lab_UT.dictrl.N_97_mux_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m40_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m40_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m40_LC_8_14_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \Lab_UT.dictrl.m40_LC_8_14_3  (
            .in0(N__19955),
            .in1(_gnd_net_),
            .in2(N__20220),
            .in3(N__20078),
            .lcout(\Lab_UT.dictrl.N_97_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_0_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_0_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_0_LC_8_14_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_0_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__23123),
            .in2(_gnd_net_),
            .in3(N__23983),
            .lcout(\Lab_UT.dictrl.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_2_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_2_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_2_LC_8_14_5 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_2_LC_8_14_5  (
            .in0(N__23982),
            .in1(_gnd_net_),
            .in2(N__23155),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_0_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_0_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_0_LC_8_14_6 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_0_LC_8_14_6  (
            .in0(N__17268),
            .in1(N__17310),
            .in2(N__17217),
            .in3(N__22979),
            .lcout(\Lab_UT.dictrl.next_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_1_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_1_LC_8_14_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_1_LC_8_14_7  (
            .in0(N__24294),
            .in1(N__19227),
            .in2(N__24555),
            .in3(N__24578),
            .lcout(\Lab_UT.dictrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_4_LC_8_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_4_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_4_LC_8_15_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_4_LC_8_15_0  (
            .in0(N__19822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19314),
            .lcout(\Lab_UT.dictrl.g2_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_8_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_8_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__19311),
            .in2(_gnd_net_),
            .in3(N__19819),
            .lcout(\Lab_UT.dictrl.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_15_LC_8_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_15_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_15_LC_8_15_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_15_LC_8_15_2  (
            .in0(N__19823),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24013),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_6_LC_8_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_6_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_6_LC_8_15_3 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_6_LC_8_15_3  (
            .in0(N__19357),
            .in1(N__17304),
            .in2(N__17295),
            .in3(N__24293),
            .lcout(\Lab_UT.dictrl.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_4_LC_8_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_4_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_4_LC_8_15_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_4_LC_8_15_4  (
            .in0(N__19821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19313),
            .lcout(\Lab_UT.dictrl.g2_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_4_LC_8_15_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_4_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_4_LC_8_15_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_4_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__19312),
            .in2(_gnd_net_),
            .in3(N__19820),
            .lcout(\Lab_UT.dictrl.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_6_LC_8_15_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_6_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_6_LC_8_15_6 .LUT_INIT=16'b1100110100000001;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_6_LC_8_15_6  (
            .in0(N__19226),
            .in1(N__24014),
            .in2(N__19736),
            .in3(N__19538),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1462_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_3_LC_8_15_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_3_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNO_3_LC_8_15_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNO_3_LC_8_15_7  (
            .in0(N__24015),
            .in1(N__17283),
            .in2(N__17277),
            .in3(N__17274),
            .lcout(\Lab_UT.dictrl.N_1460_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_8_LC_8_16_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_8_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_8_LC_8_16_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_8_LC_8_16_1  (
            .in0(N__20090),
            .in1(N__20216),
            .in2(_gnd_net_),
            .in3(N__19957),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_97_mux_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_5_LC_8_16_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_5_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_5_LC_8_16_2 .LUT_INIT=16'b0010001011101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_5_LC_8_16_2  (
            .in0(N__17580),
            .in1(N__19824),
            .in2(N__17568),
            .in3(N__19724),
            .lcout(\Lab_UT.dictrl.N_1102_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI316V_8_LC_9_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI316V_8_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI316V_8_LC_9_1_0 .LUT_INIT=16'b0001010000001010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI316V_8_LC_9_1_0  (
            .in0(N__24894),
            .in1(N__23277),
            .in2(N__24954),
            .in3(N__21135),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_9_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI9006_8_LC_9_1_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.w_addr_user_nesr_RNI9006_8_LC_9_1_1  (
            .in0(N__23543),
            .in1(N__20872),
            .in2(_gnd_net_),
            .in3(N__17558),
            .lcout(),
            .ltout(\uu2.un3_w_addr_user_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIINVH_2_LC_9_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIINVH_2_LC_9_1_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu2.w_addr_user_RNIINVH_2_LC_9_1_2  (
            .in0(N__21015),
            .in1(N__17523),
            .in2(N__17487),
            .in3(N__17484),
            .lcout(\uu2.un3_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_5_LC_9_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_5_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_5_LC_9_1_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_5_LC_9_1_3  (
            .in0(N__23278),
            .in1(N__23418),
            .in2(N__23385),
            .in3(N__23471),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_5C_net ),
            .ce(N__17448),
            .sr(N__25778));
    defparam \uu2.w_addr_displaying_fast_RNI3FPC1_1_LC_9_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI3FPC1_1_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI3FPC1_1_LC_9_2_0 .LUT_INIT=16'b0101101001000010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI3FPC1_1_LC_9_2_0  (
            .in0(N__20789),
            .in1(N__17367),
            .in2(N__17421),
            .in3(N__17687),
            .lcout(\uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIUO0E_1_LC_9_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIUO0E_1_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIUO0E_1_LC_9_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIUO0E_1_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__17415),
            .in2(_gnd_net_),
            .in3(N__20788),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(\uu2.bitmap_pmux_sn_N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIRB2A1_4_LC_9_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIRB2A1_4_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIRB2A1_4_LC_9_2_2 .LUT_INIT=16'b1010001101010011;
    LogicCell40 \uu2.w_addr_displaying_RNIRB2A1_4_LC_9_2_2  (
            .in0(N__17419),
            .in1(N__17653),
            .in2(N__17385),
            .in3(N__17366),
            .lcout(\uu2.bitmap_pmux_sn_m15_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIMLNS2_1_LC_9_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIMLNS2_1_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIMLNS2_1_LC_9_2_3 .LUT_INIT=16'b0101000010000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIMLNS2_1_LC_9_2_3  (
            .in0(N__17688),
            .in1(N__20610),
            .in2(N__17679),
            .in3(N__17670),
            .lcout(\uu2.bitmap_pmux_29_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_LC_9_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_LC_9_2_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.w_addr_displaying_3_LC_9_2_4  (
            .in0(N__17655),
            .in1(N__20755),
            .in2(_gnd_net_),
            .in3(N__17637),
            .lcout(\uu2.w_addr_displayingZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3C_net ),
            .ce(),
            .sr(N__25775));
    defparam \Lab_UT.dictrl.m12_2_LC_9_2_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m12_2_LC_9_2_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m12_2_LC_9_2_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.m12_2_LC_9_2_5  (
            .in0(N__18764),
            .in1(N__20508),
            .in2(_gnd_net_),
            .in3(N__18587),
            .lcout(\Lab_UT.dictrl.m12Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_9_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_9_3_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_215_LC_9_3_0  (
            .in0(N__24768),
            .in1(N__24741),
            .in2(N__24693),
            .in3(N__24636),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__25772));
    defparam \uu2.bitmap_RNIE8OP_212_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIE8OP_212_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIE8OP_212_LC_9_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNIE8OP_212_LC_9_3_1  (
            .in0(N__24909),
            .in1(N__24828),
            .in2(_gnd_net_),
            .in3(N__17613),
            .lcout(),
            .ltout(\uu2.N_198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0SET1_3_LC_9_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0SET1_3_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0SET1_3_LC_9_3_2 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \uu2.w_addr_displaying_RNI0SET1_3_LC_9_3_2  (
            .in0(N__25090),
            .in1(N__20743),
            .in2(N__17607),
            .in3(N__24804),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIPTJR3_3_LC_9_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIPTJR3_3_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIPTJR3_3_LC_9_3_3 .LUT_INIT=16'b0111000001111010;
    LogicCell40 \uu2.w_addr_displaying_RNIPTJR3_3_LC_9_3_3  (
            .in0(N__20744),
            .in1(N__17604),
            .in2(N__17595),
            .in3(N__17592),
            .lcout(\uu2.bitmap_pmux_27_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_9_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_9_4_1 .LUT_INIT=16'b0010011110011111;
    LogicCell40 \uu2.bitmap_93_LC_9_4_1  (
            .in0(N__21409),
            .in1(N__21504),
            .in2(N__21457),
            .in3(N__21550),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__25770));
    defparam \uu2.bitmap_221_LC_9_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_9_4_2 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_221_LC_9_4_2  (
            .in0(N__21549),
            .in1(N__21447),
            .in2(N__21513),
            .in3(N__21408),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__25770));
    defparam \uu2.w_addr_displaying_0_rep1_RNINHPP1_LC_9_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_RNINHPP1_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_0_rep1_RNINHPP1_LC_9_4_3 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_RNINHPP1_LC_9_4_3  (
            .in0(N__20756),
            .in1(N__17805),
            .in2(N__17772),
            .in3(N__17760),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_25_i_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI5BFC3_3_LC_9_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI5BFC3_3_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI5BFC3_3_LC_9_4_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.w_addr_displaying_RNI5BFC3_3_LC_9_4_4  (
            .in0(N__20757),
            .in1(N__21147),
            .in2(N__17754),
            .in3(N__17727),
            .lcout(\uu2.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI95TJ_93_LC_9_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI95TJ_93_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI95TJ_93_LC_9_4_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.bitmap_RNI95TJ_93_LC_9_4_5  (
            .in0(N__17739),
            .in1(N__17733),
            .in2(_gnd_net_),
            .in3(N__21131),
            .lcout(\uu2.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m43_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m43_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m43_LC_9_5_0 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \Lab_UT.dispString.m43_LC_9_5_0  (
            .in0(N__21361),
            .in1(N__25560),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dispString.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIL8M54_2_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIL8M54_2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIL8M54_2_LC_9_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIL8M54_2_LC_9_5_6  (
            .in0(N__21347),
            .in1(N__17900),
            .in2(_gnd_net_),
            .in3(N__17828),
            .lcout(\Lab_UT.sec2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_9_6_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNI28771_3_LC_9_6_0  (
            .in0(N__21256),
            .in1(N__17901),
            .in2(N__17954),
            .in3(N__17712),
            .lcout(\Lab_UT.didp.un18_ce ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_9_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_9_6_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_9_6_1  (
            .in0(N__17902),
            .in1(N__17953),
            .in2(_gnd_net_),
            .in3(N__21258),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_9_6_2 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_9_6_2  (
            .in0(N__22523),
            .in1(N__26412),
            .in2(N__17721),
            .in3(N__17713),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_9_6_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_9_6_3  (
            .in0(N__21998),
            .in1(N__22643),
            .in2(N__17718),
            .in3(N__17714),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26162),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_6_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_6_4  (
            .in0(N__21257),
            .in1(_gnd_net_),
            .in2(N__17955),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_6_5 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_6_5  (
            .in0(N__17903),
            .in1(N__22522),
            .in2(N__17910),
            .in3(N__26730),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_9_6_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_9_6_6  (
            .in0(N__17904),
            .in1(N__22642),
            .in2(N__17907),
            .in3(N__21997),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26162),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_9_6_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_9_6_7  (
            .in0(N__22641),
            .in1(N__18048),
            .in2(N__21999),
            .in3(N__21259),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26162),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_4_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_4_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_4_LC_9_7_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dispString.m49_4_LC_9_7_1  (
            .in0(N__17899),
            .in1(N__17845),
            .in2(N__25599),
            .in3(N__17821),
            .lcout(),
            .ltout(\Lab_UT.dispString.m49Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_LC_9_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dispString.m49_LC_9_7_2  (
            .in0(N__17874),
            .in1(N__21171),
            .in2(N__17868),
            .in3(N__17964),
            .lcout(\Lab_UT.dispString.N_128_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNINM4L3_2_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNINM4L3_2_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNINM4L3_2_LC_9_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNINM4L3_2_LC_9_7_3  (
            .in0(N__25598),
            .in1(N__21327),
            .in2(_gnd_net_),
            .in3(N__17846),
            .lcout(\Lab_UT.sec1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_2_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26722),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26154),
            .ce(N__18014),
            .sr(N__25810));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH4M54_0_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH4M54_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH4M54_0_LC_9_7_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIH4M54_0_LC_9_7_5  (
            .in0(N__21303),
            .in1(N__17939),
            .in2(_gnd_net_),
            .in3(N__17999),
            .lcout(\Lab_UT.sec2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_9_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_0_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21802),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26154),
            .ce(N__18014),
            .sr(N__25810));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_0 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_0  (
            .in0(N__21263),
            .in1(N__25520),
            .in2(N__22524),
            .in3(N__17936),
            .lcout(\Lab_UT.didp.countrce1.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_8_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__25879),
            .in2(_gnd_net_),
            .in3(N__18039),
            .lcout(\Lab_UT.didp.regrce1.LdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_11_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_11_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_11_LC_9_8_3 .LUT_INIT=16'b0000100100000000;
    LogicCell40 \Lab_UT.dispString.m49_11_LC_9_8_3  (
            .in0(N__17935),
            .in1(N__17998),
            .in2(N__17982),
            .in3(N__17970),
            .lcout(\Lab_UT.dispString.m49Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_8_5 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_8_5  (
            .in0(N__17937),
            .in1(N__22521),
            .in2(_gnd_net_),
            .in3(N__21804),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_9_8_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_9_8_6  (
            .in0(N__21986),
            .in1(N__22644),
            .in2(N__17958),
            .in3(N__17938),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26148),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_9_9_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_9_9_0  (
            .in0(N__24536),
            .in1(N__22766),
            .in2(N__23162),
            .in3(N__18225),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(\Lab_UT.LdMtens_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_9_9_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.didp.ce_RNIDJKH1_3_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17913),
            .in3(N__22334),
            .lcout(\Lab_UT.didp.un1_dicLdMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_9_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_9_2  (
            .in0(N__18395),
            .in1(N__21803),
            .in2(_gnd_net_),
            .in3(N__21959),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_9_3 .LUT_INIT=16'b0101000001000001;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_9_9_3  (
            .in0(N__22184),
            .in1(N__18399),
            .in2(N__18414),
            .in3(N__22335),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26140),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_9_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_9_4  (
            .in0(N__25519),
            .in1(N__22267),
            .in2(N__18406),
            .in3(N__21960),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_9_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_9_9_5  (
            .in0(N__22185),
            .in1(N__22268),
            .in2(N__18375),
            .in3(N__18359),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26140),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_6_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_6_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_6_LC_9_10_0 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_6_LC_9_10_0  (
            .in0(N__24368),
            .in1(N__23984),
            .in2(N__19527),
            .in3(N__19666),
            .lcout(\Lab_UT.dictrl.N_1462_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJ_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJ_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJ_LC_9_10_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJ_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__18271),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_0_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_9_10_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_9_10_4  (
            .in0(N__18233),
            .in1(N__24485),
            .in2(N__22113),
            .in3(N__18171),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26133),
            .ce(),
            .sr(N__25814));
    defparam \Lab_UT.didp.ce_1_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_9_10_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_9_10_5  (
            .in0(N__22143),
            .in1(N__22108),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26133),
            .ce(),
            .sr(N__25814));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_8_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_8_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_8_LC_9_11_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_8_LC_9_11_0  (
            .in0(N__19203),
            .in1(N__18158),
            .in2(_gnd_net_),
            .in3(N__19049),
            .lcout(\Lab_UT.dictrl.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_6_1_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_6_1_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_6_1_LC_9_11_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_6_1_LC_9_11_1  (
            .in0(N__18159),
            .in1(N__21786),
            .in2(_gnd_net_),
            .in3(N__19712),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_i_a4_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_4_1_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_4_1_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_4_1_LC_9_11_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_4_1_LC_9_11_2  (
            .in0(N__19204),
            .in1(N__19059),
            .in2(N__19053),
            .in3(N__19050),
            .lcout(\Lab_UT.dictrl.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITVU03_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITVU03_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITVU03_LC_9_11_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNITVU03_LC_9_11_3  (
            .in0(N__18948),
            .in1(N__19961),
            .in2(N__18934),
            .in3(N__19711),
            .lcout(\Lab_UT.dictrl.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_LC_9_12_0 .LUT_INIT=16'b0100010000000100;
    LogicCell40 \Lab_UT.dictrl.m22_LC_9_12_0  (
            .in0(N__18569),
            .in1(N__20191),
            .in2(N__18771),
            .in3(N__18651),
            .lcout(\Lab_UT.dictrl.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_8_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_8_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_8_LC_9_12_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_8_LC_9_12_2  (
            .in0(N__18570),
            .in1(N__20192),
            .in2(_gnd_net_),
            .in3(N__19960),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_97_mux_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_5_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_5_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_5_LC_9_12_3 .LUT_INIT=16'b0010001011101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_5_LC_9_12_3  (
            .in0(N__18471),
            .in1(N__19833),
            .in2(N__18459),
            .in3(N__19716),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1102_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_3_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_3_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_3_LC_9_12_4 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_3_LC_9_12_4  (
            .in0(N__18456),
            .in1(N__18444),
            .in2(N__18435),
            .in3(N__24039),
            .lcout(\Lab_UT.dictrl.N_1460_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_LC_9_13_0 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_LC_9_13_0  (
            .in0(N__18431),
            .in1(N__24146),
            .in2(N__19458),
            .in3(N__19328),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1106_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIDHBB9_0_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDHBB9_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDHBB9_0_LC_9_13_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIDHBB9_0_LC_9_13_1  (
            .in0(N__24544),
            .in1(N__20532),
            .in2(N__18417),
            .in3(N__24277),
            .lcout(\Lab_UT.dictrl.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_1_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_0_LC_9_13_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.g1_1_0_LC_9_13_2  (
            .in0(N__20070),
            .in1(N__20395),
            .in2(_gnd_net_),
            .in3(N__19448),
            .lcout(\Lab_UT.dictrl.g1_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m28_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m28_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m28_LC_9_13_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Lab_UT.dictrl.m28_LC_9_13_3  (
            .in0(N__19449),
            .in1(_gnd_net_),
            .in2(N__20407),
            .in3(N__20071),
            .lcout(\Lab_UT.dictrl.N_59 ),
            .ltout(\Lab_UT.dictrl.N_59_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_0_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_0_LC_9_13_4 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_0_LC_9_13_4  (
            .in0(N__19351),
            .in1(N__24145),
            .in2(N__19335),
            .in3(N__19326),
            .lcout(\Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNICN0J_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNICN0J_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep2_esr_RNICN0J_LC_9_13_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep2_esr_RNICN0J_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__19327),
            .in2(_gnd_net_),
            .in3(N__19832),
            .lcout(\Lab_UT.dictrl.g2_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_50_LC_9_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_50_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_50_LC_9_14_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.g0_50_LC_9_14_0  (
            .in0(N__20322),
            .in1(N__20086),
            .in2(N__20223),
            .in3(N__20594),
            .lcout(\Lab_UT.dictrl.N_40_5 ),
            .ltout(\Lab_UT.dictrl.N_40_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_6_LC_9_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_6_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_6_LC_9_14_1 .LUT_INIT=16'b1000100010001101;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_6_LC_9_14_1  (
            .in0(N__23966),
            .in1(N__19528),
            .in2(N__19230),
            .in3(N__19714),
            .lcout(\Lab_UT.dictrl.N_1462_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_43_LC_9_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_43_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_43_LC_9_14_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.g0_43_LC_9_14_2  (
            .in0(N__20321),
            .in1(N__20082),
            .in2(N__20222),
            .in3(N__20592),
            .lcout(\Lab_UT.dictrl.N_40_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_26_LC_9_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_26_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_26_LC_9_14_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_26_LC_9_14_3  (
            .in0(N__20593),
            .in1(N__20207),
            .in2(N__20093),
            .in3(N__20320),
            .lcout(\Lab_UT.dictrl.N_40_2 ),
            .ltout(\Lab_UT.dictrl.N_40_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_6_LC_9_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_6_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_6_LC_9_14_4 .LUT_INIT=16'b1100110000000101;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_6_LC_9_14_4  (
            .in0(N__19713),
            .in1(N__19534),
            .in2(N__19215),
            .in3(N__23965),
            .lcout(\Lab_UT.dictrl.N_1462_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_64_LC_9_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_64_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_64_LC_9_14_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.g0_64_LC_9_14_5  (
            .in0(N__20591),
            .in1(N__20206),
            .in2(N__20092),
            .in3(N__20319),
            .lcout(\Lab_UT.dictrl.N_40_7 ),
            .ltout(\Lab_UT.dictrl.N_40_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIIKGR3_1_LC_9_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIIKGR3_1_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIIKGR3_1_LC_9_14_6 .LUT_INIT=16'b1100110000000101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIIKGR3_1_LC_9_14_6  (
            .in0(N__19715),
            .in1(N__19533),
            .in2(N__20526),
            .in3(N__23967),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1462_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNIQRMCB_LC_9_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNIQRMCB_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNIQRMCB_LC_9_14_7 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNIQRMCB_LC_9_14_7  (
            .in0(N__23968),
            .in1(N__20523),
            .in2(N__20517),
            .in3(N__20514),
            .lcout(\Lab_UT.dictrl.N_1460_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_9_15_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_9_15_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_9_LC_9_15_0  (
            .in0(N__20504),
            .in1(N__20408),
            .in2(N__20076),
            .in3(N__20318),
            .lcout(\Lab_UT.dictrl.g0_i_m2_0_a7_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_8_LC_9_15_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_8_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_8_LC_9_15_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_8_LC_9_15_1  (
            .in0(N__20219),
            .in1(N__20049),
            .in2(_gnd_net_),
            .in3(N__19962),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_97_mux_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_5_LC_9_15_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_5_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_5_LC_9_15_2 .LUT_INIT=16'b0010001011101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_5_LC_9_15_2  (
            .in0(N__19863),
            .in1(N__19843),
            .in2(N__19740),
            .in3(N__19734),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1102_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_3_LC_9_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_3_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_3_LC_9_15_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_3_LC_9_15_3  (
            .in0(N__19572),
            .in1(N__19557),
            .in2(N__19551),
            .in3(N__24055),
            .lcout(\Lab_UT.dictrl.N_1460_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_16_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_16_4 .LUT_INIT=16'b0000111110001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_16_4  (
            .in0(N__19548),
            .in1(N__24546),
            .in2(N__19542),
            .in3(N__24063),
            .lcout(\Lab_UT.dictrl.g0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_5_LC_11_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_11_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_11_1_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_5_LC_11_1_0  (
            .in0(N__20972),
            .in1(N__20930),
            .in2(N__21012),
            .in3(N__21037),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__20844));
    defparam \uu2.w_addr_user_4_LC_11_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_11_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_11_1_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.w_addr_user_4_LC_11_1_1  (
            .in0(N__20929),
            .in1(N__20999),
            .in2(_gnd_net_),
            .in3(N__20971),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__20844));
    defparam \uu2.w_addr_user_6_LC_11_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_11_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_11_1_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_11_1_2  (
            .in0(N__20973),
            .in1(N__20931),
            .in2(N__20907),
            .in3(N__20871),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_5C_net ),
            .ce(),
            .sr(N__20844));
    defparam \uu2.w_addr_displaying_RNIMNI42_3_LC_11_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIMNI42_3_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIMNI42_3_LC_11_2_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.w_addr_displaying_RNIMNI42_3_LC_11_2_0  (
            .in0(N__25102),
            .in1(N__20759),
            .in2(N__20685),
            .in3(N__24843),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI9SFF4_1_LC_11_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI9SFF4_1_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI9SFF4_1_LC_11_2_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI9SFF4_1_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__20691),
            .in2(N__20802),
            .in3(N__21087),
            .lcout(\uu2.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIR9TO_1_LC_11_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIR9TO_1_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIR9TO_1_LC_11_2_2 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIR9TO_1_LC_11_2_2  (
            .in0(N__20790),
            .in1(N__25170),
            .in2(_gnd_net_),
            .in3(N__20758),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNILMVP_180_LC_11_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNILMVP_180_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNILMVP_180_LC_11_2_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNILMVP_180_LC_11_2_3  (
            .in0(N__20674),
            .in1(N__21081),
            .in2(_gnd_net_),
            .in3(N__24900),
            .lcout(\uu2.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIBP86_0_2_LC_11_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIBP86_0_2_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIBP86_0_2_LC_11_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIBP86_0_2_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__20675),
            .in2(_gnd_net_),
            .in3(N__20634),
            .lcout(\uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_314_LC_11_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_11_3_0 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_314_LC_11_3_0  (
            .in0(N__21421),
            .in1(N__21529),
            .in2(N__21578),
            .in3(N__21475),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__25776));
    defparam \uu2.bitmap_218_LC_11_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_11_3_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_218_LC_11_3_1  (
            .in0(N__21474),
            .in1(N__21571),
            .in2(N__21531),
            .in3(N__21420),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__25776));
    defparam \uu2.bitmap_90_LC_11_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_11_3_2 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_90_LC_11_3_2  (
            .in0(N__21422),
            .in1(N__21530),
            .in2(N__21579),
            .in3(N__21476),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__25776));
    defparam \uu2.bitmap_RNIC7SJ_90_LC_11_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIC7SJ_90_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIC7SJ_90_LC_11_3_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.bitmap_RNIC7SJ_90_LC_11_3_3  (
            .in0(N__21159),
            .in1(N__21153),
            .in2(_gnd_net_),
            .in3(N__21133),
            .lcout(\uu2.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIE7RK_58_LC_11_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIE7RK_58_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIE7RK_58_LC_11_3_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNIE7RK_58_LC_11_3_5  (
            .in0(N__21080),
            .in1(N__24892),
            .in2(_gnd_net_),
            .in3(N__21384),
            .lcout(),
            .ltout(\uu2.bitmap_RNIE7RKZ0Z_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIOQVH1_7_LC_11_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIOQVH1_7_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIOQVH1_7_LC_11_3_6 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIOQVH1_7_LC_11_3_6  (
            .in0(N__21134),
            .in1(_gnd_net_),
            .in2(N__21090),
            .in3(N__21063),
            .lcout(\uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI020Q_186_LC_11_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI020Q_186_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI020Q_186_LC_11_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNI020Q_186_LC_11_3_7  (
            .in0(N__21057),
            .in1(N__24891),
            .in2(_gnd_net_),
            .in3(N__21079),
            .lcout(\uu2.bitmap_RNI020QZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_11_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_11_4_0 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_87_LC_11_4_0  (
            .in0(N__24621),
            .in1(N__24687),
            .in2(N__24730),
            .in3(N__24786),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__25773));
    defparam \uu2.bitmap_308_LC_11_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_11_4_1 .LUT_INIT=16'b0000011000011101;
    LogicCell40 \uu2.bitmap_308_LC_11_4_1  (
            .in0(N__24784),
            .in1(N__24718),
            .in2(N__24694),
            .in3(N__24619),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__25773));
    defparam \uu2.bitmap_186_LC_11_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_11_4_4 .LUT_INIT=16'b0000011100111100;
    LogicCell40 \uu2.bitmap_186_LC_11_4_4  (
            .in0(N__21428),
            .in1(N__21470),
            .in2(N__21525),
            .in3(N__21569),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__25773));
    defparam \uu2.bitmap_58_LC_11_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_11_4_5 .LUT_INIT=16'b1011011011101111;
    LogicCell40 \uu2.bitmap_58_LC_11_4_5  (
            .in0(N__21570),
            .in1(N__21517),
            .in2(N__21477),
            .in3(N__21429),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__25773));
    defparam \uu2.bitmap_52_LC_11_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_11_4_7 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_52_LC_11_4_7  (
            .in0(N__24785),
            .in1(N__24719),
            .in2(N__24695),
            .in3(N__24620),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_87C_net ),
            .ce(),
            .sr(N__25773));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_11_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_11_5_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_11_5_0  (
            .in0(N__25554),
            .in1(N__25588),
            .in2(N__25226),
            .in3(N__25297),
            .lcout(\Lab_UT.didp.un24_ce_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_11_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_11_5_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_0_LC_11_5_1  (
            .in0(N__25260),
            .in1(N__21806),
            .in2(_gnd_net_),
            .in3(N__25555),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_11_5_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_11_5_2  (
            .in0(N__25556),
            .in1(N__25330),
            .in2(N__21378),
            .in3(N__25362),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26179),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNIJI4L3_0_LC_11_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIJI4L3_0_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIJI4L3_0_LC_11_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNIJI4L3_0_LC_11_5_3  (
            .in0(N__21345),
            .in1(N__25553),
            .in2(_gnd_net_),
            .in3(N__21374),
            .lcout(\Lab_UT.sec1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNILK4L3_1_LC_11_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNILK4L3_1_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNILK4L3_1_LC_11_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNILK4L3_1_LC_11_5_4  (
            .in0(N__21221),
            .in1(N__21346),
            .in2(_gnd_net_),
            .in3(N__25296),
            .lcout(\Lab_UT.sec1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_5_LC_11_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_5_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_5_LC_11_5_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dispString.m49_5_LC_11_5_5  (
            .in0(N__21264),
            .in1(N__21220),
            .in2(N__25302),
            .in3(N__21194),
            .lcout(\Lab_UT.dispString.m49Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_11_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_11_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_1_LC_11_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25524),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26171),
            .ce(N__21828),
            .sr(N__25816));
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_11_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_11_6_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_2_LC_11_6_1  (
            .in0(_gnd_net_),
            .in1(N__26739),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26171),
            .ce(N__21828),
            .sr(N__25816));
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_11_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_3_LC_11_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26424),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26171),
            .ce(N__21828),
            .sr(N__25816));
    defparam \Lab_UT.didp.countrce3.q_0_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_11_7_0 .LUT_INIT=16'b0000110000001001;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_11_7_0  (
            .in0(N__22320),
            .in1(N__21666),
            .in2(N__26259),
            .in3(N__26458),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26164),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_11_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_11_7_1 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_11_7_1  (
            .in0(N__26457),
            .in1(N__21807),
            .in2(_gnd_net_),
            .in3(N__26531),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_11_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_11_7_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNI4EIS1_2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__22319),
            .in2(_gnd_net_),
            .in3(N__26455),
            .lcout(\Lab_UT.didp.un1_dicLdMones_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_11_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_11_7_3 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_11_7_3  (
            .in0(N__21657),
            .in1(N__26256),
            .in2(N__21660),
            .in3(N__26566),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26164),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_11_7_4 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_1_LC_11_7_4  (
            .in0(N__26530),
            .in1(N__26456),
            .in2(N__26573),
            .in3(N__25481),
            .lcout(\Lab_UT.didp.countrce3.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m49_2_LC_11_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m49_2_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m49_2_LC_11_7_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dispString.m49_2_LC_11_7_5  (
            .in0(N__21640),
            .in1(N__26562),
            .in2(N__21613),
            .in3(N__26482),
            .lcout(\Lab_UT.dispString.m49Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_1_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_11_8_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_11_8_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_11_8_0  (
            .in0(N__22147),
            .in1(_gnd_net_),
            .in2(N__22111),
            .in3(N__22302),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.ce_3_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_11_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_11_8_1  (
            .in0(N__25184),
            .in1(N__22095),
            .in2(N__22305),
            .in3(N__22148),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.reset_2_LC_11_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_11_8_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_11_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_11_8_2  (
            .in0(N__22149),
            .in1(N__25185),
            .in2(N__22112),
            .in3(N__22304),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.ce_2_LC_11_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_11_8_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_11_8_3  (
            .in0(N__22303),
            .in1(N__22094),
            .in2(_gnd_net_),
            .in3(N__22145),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_11_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_11_8_4  (
            .in0(N__22144),
            .in1(N__25183),
            .in2(N__22109),
            .in3(N__22298),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_11_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_11_8_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_11_8_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_11_8_5  (
            .in0(N__21882),
            .in1(N__22280),
            .in2(N__22221),
            .in3(N__22218),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.reset_0_LC_11_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_11_8_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_11_8_6 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_11_8_6  (
            .in0(N__22146),
            .in1(_gnd_net_),
            .in2(N__22110),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26155),
            .ce(),
            .sr(N__25811));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_11_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_11_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_11_8_7  (
            .in0(N__21972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21918),
            .lcout(\Lab_UT.didp.reset_12_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_11_9_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI5U3I_1_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__21876),
            .in2(_gnd_net_),
            .in3(N__21864),
            .lcout(\Lab_UT.didp.un1_dicLdStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_2_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_2_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_2_LC_11_9_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_2_LC_11_9_4  (
            .in0(N__23132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23958),
            .lcout(\Lab_UT.dictrl.g2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_11_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_11_9_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_11_9_6  (
            .in0(N__24535),
            .in1(N__22765),
            .in2(N__23160),
            .in3(N__24308),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_0_LC_11_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_0_LC_11_10_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_0_LC_11_10_0  (
            .in0(N__22854),
            .in1(N__22689),
            .in2(N__22674),
            .in3(N__22980),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_11_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_11_10_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_11_10_1 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_LC_11_10_1  (
            .in0(N__23204),
            .in1(N__22567),
            .in2(N__22662),
            .in3(N__22605),
            .lcout(\Lab_UT.LdSones_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26143),
            .ce(N__22486),
            .sr(N__25815));
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_11_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_11_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_11_10_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_LC_11_10_2  (
            .in0(N__23001),
            .in1(N__22604),
            .in2(N__22569),
            .in3(N__23203),
            .lcout(\Lab_UT.LdStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26143),
            .ce(N__22486),
            .sr(N__25815));
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_11_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_11_10_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI51AM_0_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__22659),
            .in2(_gnd_net_),
            .in3(N__22650),
            .lcout(\Lab_UT.didp.un1_dicLdSones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_11_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_11_10_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_LC_11_10_4  (
            .in0(N__23172),
            .in1(N__22603),
            .in2(N__22568),
            .in3(N__23202),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26143),
            .ce(N__22486),
            .sr(N__25815));
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_0_1_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_0_1_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIP2CG_0_1_LC_11_11_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIP2CG_0_1_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__23133),
            .in2(_gnd_net_),
            .in3(N__23827),
            .lcout(\Lab_UT.dictrl.g2_5 ),
            .ltout(\Lab_UT.dictrl.g2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIRP7EL_LC_11_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIRP7EL_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIRP7EL_LC_11_11_1 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIRP7EL_LC_11_11_1  (
            .in0(N__22418),
            .in1(N__22967),
            .in2(N__22383),
            .in3(N__22370),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_11_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_LC_11_11_2  (
            .in0(N__23229),
            .in1(N__23220),
            .in2(N__23211),
            .in3(N__23208),
            .lcout(\Lab_UT.dictrl.un1_next_state66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26134),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_2_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_2_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_2_LC_11_11_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_2_LC_11_11_3  (
            .in0(N__23828),
            .in1(_gnd_net_),
            .in2(N__23161),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_0_LC_11_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_0_LC_11_11_4 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_0_LC_11_11_4  (
            .in0(N__23715),
            .in1(N__22966),
            .in2(N__23175),
            .in3(N__22833),
            .lcout(\Lab_UT.dictrl.next_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_2_LC_11_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_2_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_2_LC_11_12_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_2_LC_11_12_4  (
            .in0(N__23137),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23829),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_0_LC_11_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_0_LC_11_12_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_0_LC_11_12_5  (
            .in0(N__23013),
            .in1(N__24351),
            .in2(N__23004),
            .in3(N__22973),
            .lcout(\Lab_UT.dictrl.next_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_3_LC_11_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_3_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_3_LC_11_12_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_3_LC_11_12_6  (
            .in0(N__24306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24545),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1105_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_1_LC_11_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_1_LC_11_12_7 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_1_LC_11_12_7  (
            .in0(N__22992),
            .in1(N__24108),
            .in2(N__22983),
            .in3(N__22972),
            .lcout(\Lab_UT.dictrl.N_79_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_1_LC_11_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_1_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_8_ess_RNO_1_LC_11_13_1 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_RNO_1_LC_11_13_1  (
            .in0(N__24584),
            .in1(N__22866),
            .in2(N__24323),
            .in3(N__24543),
            .lcout(\Lab_UT.dictrl.g1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_1_LC_11_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_1_LC_11_13_4 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_1_LC_11_13_4  (
            .in0(N__22845),
            .in1(N__24309),
            .in2(N__24554),
            .in3(N__24582),
            .lcout(\Lab_UT.dictrl.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_1_LC_11_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_1_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNO_1_LC_11_13_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNO_1_LC_11_13_5  (
            .in0(N__24583),
            .in1(N__24307),
            .in2(N__24553),
            .in3(N__24372),
            .lcout(\Lab_UT.dictrl.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_4_LC_11_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_4_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_ess_RNO_4_LC_11_14_7 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_ess_RNO_4_LC_11_14_7  (
            .in0(N__24341),
            .in1(N__24305),
            .in2(N__24162),
            .in3(N__24147),
            .lcout(\Lab_UT.dictrl.N_1106_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_3_LC_11_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_3_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_RNO_3_LC_11_15_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_RNO_3_LC_11_15_4  (
            .in0(N__24099),
            .in1(N__24087),
            .in2(N__24075),
            .in3(N__24056),
            .lcout(\Lab_UT.dictrl.N_1460_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_12_2_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_12_2_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_12_2_0  (
            .in0(N__23704),
            .in1(N__23616),
            .in2(N__23544),
            .in3(N__25171),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_12_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_12_2_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uu2.w_addr_displaying_0_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(N__23327),
            .in2(_gnd_net_),
            .in3(N__25030),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__25780));
    defparam \uu2.w_addr_displaying_nesr_RNIA8E42_5_LC_12_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIA8E42_5_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIA8E42_5_LC_12_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIA8E42_5_LC_12_2_2  (
            .in0(N__23486),
            .in1(N__23417),
            .in2(N__23342),
            .in3(N__23295),
            .lcout(\uu2.N_14_i ),
            .ltout(\uu2.N_14_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI6OAF2_6_LC_12_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI6OAF2_6_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI6OAF2_6_LC_12_2_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI6OAF2_6_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23259),
            .in3(N__24936),
            .lcout(\uu2.N_15_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_0_LC_12_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_12_2_4 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_12_2_4  (
            .in0(N__25031),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24824),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__25780));
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_12_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNO_0_6_LC_12_2_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.w_addr_displaying_RNO_0_6_LC_12_2_5  (
            .in0(N__25172),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25103),
            .lcout(),
            .ltout(\uu2.N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_6_LC_12_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_LC_12_2_6 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_LC_12_2_6 .LUT_INIT=16'b1101100111001100;
    LogicCell40 \uu2.w_addr_displaying_6_LC_12_2_6  (
            .in0(N__25032),
            .in1(N__24937),
            .in2(N__24966),
            .in3(N__24963),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_0C_net ),
            .ce(),
            .sr(N__25780));
    defparam \uu2.bitmap_212_LC_12_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_12_3_1 .LUT_INIT=16'b0001000100000101;
    LogicCell40 \uu2.bitmap_212_LC_12_3_1  (
            .in0(N__24632),
            .in1(N__24692),
            .in2(N__24795),
            .in3(N__24740),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_212C_net ),
            .ce(),
            .sr(N__25779));
    defparam \uu2.bitmap_180_LC_12_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_12_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_12_3_3 .LUT_INIT=16'b0001001100111100;
    LogicCell40 \uu2.bitmap_180_LC_12_3_3  (
            .in0(N__24631),
            .in1(N__24691),
            .in2(N__24794),
            .in3(N__24739),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_212C_net ),
            .ce(),
            .sr(N__25779));
    defparam \uu2.bitmap_RNIB3QK_52_LC_12_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIB3QK_52_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIB3QK_52_LC_12_3_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.bitmap_RNIB3QK_52_LC_12_3_5  (
            .in0(N__24893),
            .in1(N__24855),
            .in2(_gnd_net_),
            .in3(N__24849),
            .lcout(\uu2.N_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNISLTD_84_LC_12_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNISLTD_84_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNISLTD_84_LC_12_3_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNISLTD_84_LC_12_3_7  (
            .in0(N__24837),
            .in1(N__24594),
            .in2(_gnd_net_),
            .in3(N__24820),
            .lcout(\uu2.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_84_LC_12_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_12_4_7 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \uu2.bitmap_84_LC_12_4_7  (
            .in0(N__24787),
            .in1(N__24723),
            .in2(N__24696),
            .in3(N__24622),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_84C_net ),
            .ce(),
            .sr(N__25777));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_12_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_12_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_3_LC_12_5_1  (
            .in0(N__25298),
            .in1(N__25586),
            .in2(_gnd_net_),
            .in3(N__25557),
            .lcout(\Lab_UT.didp.countrce2.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_12_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_12_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_2_LC_12_5_2  (
            .in0(N__25558),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25299),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_12_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_12_5_3 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_12_5_3  (
            .in0(N__25589),
            .in1(N__26738),
            .in2(N__25605),
            .in3(N__25264),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_12_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_12_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_12_5_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_12_5_4  (
            .in0(N__25587),
            .in1(N__25331),
            .in2(N__25602),
            .in3(N__25364),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26187),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_12_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_12_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_12_5_5 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_12_5_5  (
            .in0(N__25365),
            .in1(N__25191),
            .in2(N__25335),
            .in3(N__25221),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26187),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_12_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_12_5_6 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_1_LC_12_5_6  (
            .in0(N__25559),
            .in1(N__25493),
            .in2(N__25266),
            .in3(N__25300),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_12_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_12_5_7 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_12_5_7  (
            .in0(N__25301),
            .in1(N__25363),
            .in2(N__25338),
            .in3(N__25329),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26187),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_12_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_12_6_7 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_12_6_7  (
            .in0(N__25272),
            .in1(N__26423),
            .in2(N__25265),
            .in3(N__25220),
            .lcout(\Lab_UT.didp.countrce2.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_12_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_12_7_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_12_7_1  (
            .in0(N__26570),
            .in1(N__26527),
            .in2(N__26497),
            .in3(N__26228),
            .lcout(\Lab_UT.didp.countrce3.ce_12_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_12_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_12_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_12_7_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_2_LC_12_7_2  (
            .in0(N__26528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26572),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_12_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_12_7_3 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_12_7_3  (
            .in0(N__26492),
            .in1(N__26459),
            .in2(N__26742),
            .in3(N__26731),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_12_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_12_7_4 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_12_7_4  (
            .in0(N__26257),
            .in1(N__26267),
            .in2(N__26580),
            .in3(N__26493),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26172),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_12_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_12_7_5 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_3_LC_12_7_5  (
            .in0(N__26571),
            .in1(N__26529),
            .in2(N__26498),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_12_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_12_7_6 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_12_7_6  (
            .in0(N__26229),
            .in1(N__26460),
            .in2(N__26427),
            .in3(N__26388),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_12_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_12_7_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_12_7_7  (
            .in0(N__26268),
            .in1(N__26258),
            .in2(N__26238),
            .in3(N__26230),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__26172),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_ctle_LC_12_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_ctle_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep2_esr_ctle_LC_12_8_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep2_esr_ctle_LC_12_8_7  (
            .in0(_gnd_net_),
            .in1(N__25918),
            .in2(_gnd_net_),
            .in3(N__25875),
            .lcout(bu_rx_data_rdy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
