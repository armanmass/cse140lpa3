-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 19 2019 07:10:59

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19571\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19546\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19536\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19518\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19490\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19436\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19400\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19382\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19179\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19173\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19142\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19133\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19055\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19038\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19029\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18952\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18904\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18902\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18890\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18874\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18707\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18704\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18700\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18688\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18668\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18656\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18653\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18527\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18505\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18439\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18179\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18122\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18017\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17946\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17931\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17877\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17870\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17703\ : std_logic;
signal \N__17702\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17652\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17459\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17411\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17358\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17318\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17258\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17234\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17228\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17150\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17054\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17039\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17031\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17003\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16877\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16811\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16790\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16402\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16295\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16256\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16199\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16187\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16112\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15992\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15914\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15787\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15644\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15332\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15180\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15139\ : std_logic;
signal \N__15136\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15124\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14900\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14731\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14525\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14519\ : std_logic;
signal \N__14516\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14498\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14400\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14246\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14117\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13985\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13862\ : std_logic;
signal \N__13859\ : std_logic;
signal \N__13856\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12940\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8957\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \INVuu2.r_data_reg_4C_net\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \uu0.un88_ci_3_cascade_\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.un4_l_count_13_cascade_\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.un4_l_count_16\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.un404_ci_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \uu0.sec_clkDZ0\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \INVuu2.bitmap_111C_net\ : std_logic;
signal \uu0.un55_ci\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \Lab_UT.alarmchar10_i_2\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_2\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_6\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_7\ : std_logic;
signal \uu2.N_102_cascade_\ : std_logic;
signal \uu2.N_61_i\ : std_logic;
signal \INVuu2.w_addr_user_8C_net\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_4\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_3_6\ : std_logic;
signal \uu2.mem0.g1_3_0_cascade_\ : std_logic;
signal \uu2.mem0.N_63_0_i\ : std_logic;
signal \uu2.mem0.G_17_0_0_0\ : std_logic;
signal \N_72_mux\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_3\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_2_6\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_cascade_\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.N_105\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \INVuu2.w_addr_user_1C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.alarmchar_2_1_1\ : std_logic;
signal \resetGen.reset_count_2_0_4_cascade_\ : std_logic;
signal \Lab_UT.alarmchar10\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_4\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.un241_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu2.un1_l_count_1_2_0_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu2.un1_l_count_2_2_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \uu2.N_155\ : std_logic;
signal \uu2.N_106\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.N_102\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.N_97\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \INVuu2.w_addr_user_nesr_0C_net\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_12\ : std_logic;
signal \uu2.N_41_0_cascade_\ : std_logic;
signal \uu2.N_132_mux\ : std_logic;
signal \uu2.N_132_mux_cascade_\ : std_logic;
signal \uu2.mem0.N_94_i\ : std_logic;
signal \uu2.N_15_i\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_0C_net\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_5\ : std_logic;
signal \uu2.mem0.N_13_1_0_0\ : std_logic;
signal \uu2.mem0.i14_mux_0_0_0_cascade_\ : std_logic;
signal \uu2.mem0.N_8_0_0_1\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_6\ : std_logic;
signal \Lab_UT.bcd2segment1.m68_bmZ0\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_a2Z0Z_4\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \uu2.w_data_i_o2_4Z0Z_0_cascade_\ : std_logic;
signal \N_96_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.m59_bmZ0\ : std_logic;
signal \Lab_UT.bcd2segment1.m52_amZ0\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.m59_amZ0\ : std_logic;
signal \Lab_UT.dictrl.un1_next_alarmstate21_0\ : std_logic;
signal \Lab_UT.cnt_0\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_0_0\ : std_logic;
signal \Lab_UT.dictrl.G_74\ : std_logic;
signal \Lab_UT.bcd2segment1.N_187_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.N_189_cascade_\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.mem0.N_107_0_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_1\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \uu2.mem0.N_130_mux_cascade_\ : std_logic;
signal \uu2.mem0.N_54_0_i\ : std_logic;
signal \uu2.mem0.N_17_0_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_5\ : std_logic;
signal \uu2.mem0.N_107_0_0\ : std_logic;
signal \uu2.mem0.N_74_0_0_1\ : std_logic;
signal \uu2.mem0.g0_7_0_0_2_cascade_\ : std_logic;
signal \uu2.mem0.N_3_0_cascade_\ : std_logic;
signal \uu2.mem0.N_98_0_0_0\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \uu2.N_1585_0_0\ : std_logic;
signal \Lab_UT.bcd2segment1.i6_mux_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.m68_amZ0\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal rst : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_0\ : std_logic;
signal clk : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_\ : std_logic;
signal \uu2.mem0.g1_2_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0\ : std_logic;
signal \uu2.mem0.g0_7_0_0_1\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_3C_net\ : std_logic;
signal \Lab_UT.alarmchar9_cascade_\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment1.N_160\ : std_logic;
signal \Lab_UT.bcd2segment1.i5_mux_cascade_\ : std_logic;
signal \Lab_UT.cnt_2\ : std_logic;
signal \Lab_UT.bcd2segment1.m42_amZ0_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.m52_bmZ0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_42_i\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.idle_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_222_cascade_\ : std_logic;
signal \Lab_UT.dictrl.alarmstateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_i_3_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \Lab_UT.q_5_1_cascade_\ : std_logic;
signal \buart.Z_rx.ser_clk_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z4\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_194_cascade_\ : std_logic;
signal \uu2.mem0.N_92_0_cascade_\ : std_logic;
signal \uu2.mem0.m73_ns_1_0\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_1_4\ : std_logic;
signal \INVuu2.bitmap_90C_net\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.mem0.N_92_0_0_cascade_\ : std_logic;
signal \uu2.mem0.m73_ns_1_0_0_1\ : std_logic;
signal \uu2.mem0.N_74_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_34\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \uu2.mem0.N_93_i\ : std_logic;
signal \uu2.mem0.N_57_0_0\ : std_logic;
signal \uu2.mem0.N_67_0\ : std_logic;
signal \uu2.mem0.g0_1_cascade_\ : std_logic;
signal \uu2.mem0.g0_2\ : std_logic;
signal \uu2.mem0.i14_mux\ : std_logic;
signal \uu2.mem0.N_126_0\ : std_logic;
signal \uu2.mem0.g0_1_3_cascade_\ : std_logic;
signal \uu2.mem0.G_13_0_a2_0_1\ : std_logic;
signal \uu2.mem0.N_22_cascade_\ : std_logic;
signal \uu2.mem0.N_66_0_i\ : std_logic;
signal \uu2.mem0.g0_i_m2_1\ : std_logic;
signal \uu2.mem0.g2_0_0_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1\ : std_logic;
signal \uu2.N_67_1_0\ : std_logic;
signal \uu2.N_67_1_0_cascade_\ : std_logic;
signal \uu2.mem0.N_55_0_0_0\ : std_logic;
signal \uu2.mem0.g2_1\ : std_logic;
signal \INVuu2.w_addr_displaying_1C_net\ : std_logic;
signal \Lab_UT.bcd2segment1.N_250_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.i2_mux_cascade_\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.m95_i_m2_i_m2_1_cascade_\ : std_logic;
signal \uu2.N_16_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_displaying_3_rep1_nesrC_net\ : std_logic;
signal \Lab_UT.N_27_i\ : std_logic;
signal \resetGen.escKeyZ0Z_4\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \Lab_UT.didp.did_alarmMatch_1_cascade_\ : std_logic;
signal \Lab_UT.zero\ : std_logic;
signal \Lab_UT.alarmMatch\ : std_logic;
signal \Lab_UT.didp.countrce3.did_alarmMatch_0\ : std_logic;
signal \Lab_UT.q_5_3\ : std_logic;
signal \Lab_UT.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.q_5_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_1\ : std_logic;
signal \Lab_UT.dictrl.N_97_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_\ : std_logic;
signal \resetGen.escKeyZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_0_1\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5\ : std_logic;
signal \Lab_UT.dictrl.un1_state_16_cascade_\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_1 : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.bcd2segment1.N_127_mux_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.N_235_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.N_237_cascade_\ : std_logic;
signal \INVuu2.bitmap_162C_net\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.N_101_0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_242_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_\ : std_logic;
signal \uu2.N_1580_0_cascade_\ : std_logic;
signal \uu2.N_77_0\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.N_1581_0\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \INVuu2.bitmap_75C_net\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \uu2.mem0.N_134_mux_cascade_\ : std_logic;
signal \uu2.w_data_i_0_tzZ0Z_0\ : std_logic;
signal \uu2.mem0.N_60_0_i\ : std_logic;
signal \uu2.mem0.N_55_0\ : std_logic;
signal \uu2.N_126_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_67\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_66\ : std_logic;
signal \uu2.N_126\ : std_logic;
signal \uu2.mem0.g0_7_0_0\ : std_logic;
signal \uu2.mem0.N_57_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_5_1\ : std_logic;
signal \uu2.mem0.g0_7_0_3\ : std_logic;
signal \uu2.N_16\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_57\ : std_logic;
signal \uu2.mem0.N_13_0\ : std_logic;
signal \uu2.N_8\ : std_logic;
signal \uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_4\ : std_logic;
signal \INVuu2.w_addr_displaying_4_rep1C_net\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \uu2.N_9_i\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \uu2.mem0.N_9_cascade_\ : std_logic;
signal \uu2.mem0.N_15\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.mem0.N_7\ : std_logic;
signal \uu2.mem0.m317_0_a6_0_cascade_\ : std_logic;
signal \uu2.mem0.N_6_0\ : std_logic;
signal \uu2.mem0.m317_0_0\ : std_logic;
signal \uu2.mem0.N_11_0_0_cascade_\ : std_logic;
signal \uu2.mem0.N_6_0_0_0\ : std_logic;
signal \uu2.w_addr_displaying_4_repZ0Z1\ : std_logic;
signal \uu2.mem0.N_5_0\ : std_logic;
signal \uu2.mem0.N_14\ : std_logic;
signal \uu2.mem0.g1_2_2_2_1\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \Lab_UT.bcd2segment1.N_239\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.N_115\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \INVuu2.bitmap_34C_net\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_0\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \INVuu2.bitmap_180C_net\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.N_9_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment1.N_181\ : std_logic;
signal \Lab_UT.bcd2segment1.N_229\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.bcd2segment1.N_233\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.dicRun_2_reti\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_set\ : std_logic;
signal \buart.Z_rx.bitcount_lm_3_cascade_\ : std_logic;
signal \Lab_UT.m72_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1\ : std_logic;
signal \Lab_UT.un1_state_13\ : std_logic;
signal \Lab_UT.un1_state_13_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.un1_state_11\ : std_logic;
signal \Lab_UT.dictrl.un1_state_11_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1\ : std_logic;
signal \Lab_UT.bcd2segment1.N_264\ : std_logic;
signal \Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state16Z0Z_5\ : std_logic;
signal \Lab_UT.m68_0_ns_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state16Z0Z_4\ : std_logic;
signal \Lab_UT.state_3\ : std_logic;
signal \Lab_UT.state_1\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.state_2\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_0Z0Z_1\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.m76_am_1\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \Lab_UT.bcd2segment1.N_244\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \Lab_UT.bcd2segment1.N_246_cascade_\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.bcd2segment1.N_248_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.m76_bm_1_0\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \INVuu2.bitmap_168C_net\ : std_logic;
signal \uu2.mem0.g1_2_2\ : std_logic;
signal \uu2.mem0.g2_0_0_0_0\ : std_logic;
signal \uu2.mem0.g2_2\ : std_logic;
signal \uu2.w_addr_displaying_2_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_4_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_69\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_displaying_ness_6C_net\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_0\ : std_logic;
signal \uu2.mem0.G_13_0_a2_1_cascade_\ : std_logic;
signal \uu2.mem0.G_13_0_a3_1_2\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \uu2.mem0.G_13_0_a2_2_cascade_\ : std_logic;
signal \N_96\ : std_logic;
signal \uu2.mem0.G_13_0_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0\ : std_logic;
signal \uu2.N_12_i_cascade_\ : std_logic;
signal \uu2.N_67\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.un21_w_addr_displaying_i\ : std_logic;
signal \uu2.N_12_i\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \INVuu2.w_addr_displaying_7_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.N_272_cascade_\ : std_logic;
signal \uu2.mem0.m317_0_a6_1_0\ : std_logic;
signal \uu2.mem0.N_13\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \Lab_UT.Run\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \INVuu2.bitmap_58C_net\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.w_addr_displaying_8_repZ0Z1\ : std_logic;
signal \uu2.N_272\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z2\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_\ : std_logic;
signal \uu2.mem0.N_294\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \uu2.mem0.N_271\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_80\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.w_addr_displaying_7_repZ0Z1\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \uu2.mem0.N_98_0\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_166\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_RNO_0Z0Z_3\ : std_logic;
signal \bfn_9_10_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \buart.Z_rx.bitcount_lm_4\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_1\ : std_logic;
signal \Lab_UT.cnt_3\ : std_logic;
signal \Lab_UT.cnt_1\ : std_logic;
signal \Lab_UT.bcd2segment1.m42_bmZ0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \buart.Z_rx.bitcount_lm_0\ : std_logic;
signal \buart.Z_rx.un1_sample_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_3\ : std_logic;
signal \Lab_UT.m68_0_ns\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_lm_1\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_lm_2\ : std_logic;
signal \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_1\ : std_logic;
signal \Lab_UT.dictrl.un1_state_21_reti_i\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_rx.valid_0_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \bu_rx_data_rdy_cascade_\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_rx.idle_0\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal \buart.Z_rx.ser_clk_2\ : std_logic;
signal \buart.Z_rx.ser_clk_3\ : std_logic;
signal \buart.Z_rx.idle_cascade_\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \buart.Z_rx.bitcountlde_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_2\ : std_logic;
signal \Lab_UT.state_i_3_3\ : std_logic;
signal \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_retZ0Z_4\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_0\ : std_logic;
signal \Lab_UT.state_i_3_1\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_2 : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_0\ : std_logic;
signal \Lab_UT.bcd2segment1.N_192\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_5\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_3\ : std_logic;
signal \Lab_UT.bcd2segment2.segmentUQ_0_4\ : std_logic;
signal \Lab_UT.three_2_cascade_\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.didp.countrce2.un15_ce_2\ : std_logic;
signal \Lab_UT.didp.countrce2.un15_ce_2_cascade_\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.three_2_0\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.dictrl.dicRun_2\ : std_logic;
signal \Lab_UT.state_i_3_2\ : std_logic;
signal \Lab_UT.state_0\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.nine\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.q_RNI84NN1_2\ : std_logic;
signal rst_g : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_g : std_logic;
signal \oneSecStrb_i\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal sd_wire : std_logic;
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    sd <= sd_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__7230\&\N__7599\&\N__7572\&\N__7746\&\N__7689\&\N__7638\&\N__15894\&\N__15764\&\N__15848\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__8394\&\N__8403\&\N__10212\&\N__8478\&\N__8433\&\N__8412\&\N__10128\&\N__10548\&\N__12111\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__10086\&'0'&\N__11808\&'0'&\N__9192\&'0'&\N__8460\&'0'&\N__11028\&'0'&\N__10968\&'0'&\N__9171\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__7023\,
            RESETB => \N__16614\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18496\,
            RE => \N__16607\,
            WCLKE => \N__10508\,
            WCLK => \N__18495\,
            WE => \N__10509\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19573\,
            DIN => \N__19572\,
            DOUT => \N__19571\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__19573\,
            PADOUT => \N__19572\,
            PADIN => \N__19571\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19564\,
            DIN => \N__19563\,
            DOUT => \N__19562\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19564\,
            PADOUT => \N__19563\,
            PADIN => \N__19562\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19555\,
            DIN => \N__19554\,
            DOUT => \N__19553\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__19555\,
            PADOUT => \N__19554\,
            PADIN => \N__19553\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19546\,
            DIN => \N__19545\,
            DOUT => \N__19544\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__19546\,
            PADOUT => \N__19545\,
            PADIN => \N__19544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19537\,
            DIN => \N__19536\,
            DOUT => \N__19535\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19537\,
            PADOUT => \N__19536\,
            PADIN => \N__19535\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__18469\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19528\,
            DIN => \N__19527\,
            DOUT => \N__19526\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__19528\,
            PADOUT => \N__19527\,
            PADIN => \N__19526\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19519\,
            DIN => \N__19518\,
            DOUT => \N__19517\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__19519\,
            PADOUT => \N__19518\,
            PADIN => \N__19517\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19510\,
            DIN => \N__19509\,
            DOUT => \N__19508\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__19510\,
            PADOUT => \N__19509\,
            PADIN => \N__19508\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19501\,
            DIN => \N__19500\,
            DOUT => \N__19499\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19501\,
            PADOUT => \N__19500\,
            PADIN => \N__19499\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19492\,
            DIN => \N__19491\,
            DOUT => \N__19490\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__19492\,
            PADOUT => \N__19491\,
            PADIN => \N__19490\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7038\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4752\ : CascadeMux
    port map (
            O => \N__19473\,
            I => \N__19469\
        );

    \I__4751\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19458\
        );

    \I__4750\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19458\
        );

    \I__4749\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19458\
        );

    \I__4748\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19458\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__19458\,
            I => \N__19455\
        );

    \I__4746\ : Odrv4
    port map (
            O => \N__19455\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__4745\ : InMux
    port map (
            O => \N__19452\,
            I => \N__19446\
        );

    \I__4744\ : InMux
    port map (
            O => \N__19451\,
            I => \N__19446\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__19446\,
            I => \Lab_UT.three_2_0\
        );

    \I__4742\ : InMux
    port map (
            O => \N__19443\,
            I => \N__19440\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N__19437\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__19437\,
            I => \N__19425\
        );

    \I__4739\ : InMux
    port map (
            O => \N__19436\,
            I => \N__19417\
        );

    \I__4738\ : InMux
    port map (
            O => \N__19435\,
            I => \N__19417\
        );

    \I__4737\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19414\
        );

    \I__4736\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19407\
        );

    \I__4735\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19407\
        );

    \I__4734\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19407\
        );

    \I__4733\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19400\
        );

    \I__4732\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19400\
        );

    \I__4731\ : InMux
    port map (
            O => \N__19428\,
            I => \N__19400\
        );

    \I__4730\ : Span4Mux_h
    port map (
            O => \N__19425\,
            I => \N__19397\
        );

    \I__4729\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19390\
        );

    \I__4728\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19390\
        );

    \I__4727\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19390\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__19417\,
            I => \N__19387\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__19414\,
            I => \N__19382\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19382\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__19400\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__4722\ : Odrv4
    port map (
            O => \N__19397\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__19390\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__4720\ : Odrv12
    port map (
            O => \N__19387\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__4719\ : Odrv12
    port map (
            O => \N__19382\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__4718\ : CascadeMux
    port map (
            O => \N__19371\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__4717\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19364\
        );

    \I__4716\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19359\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__19364\,
            I => \N__19356\
        );

    \I__4714\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19351\
        );

    \I__4713\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19351\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__19359\,
            I => \N__19345\
        );

    \I__4711\ : Span4Mux_v
    port map (
            O => \N__19356\,
            I => \N__19340\
        );

    \I__4710\ : LocalMux
    port map (
            O => \N__19351\,
            I => \N__19340\
        );

    \I__4709\ : InMux
    port map (
            O => \N__19350\,
            I => \N__19335\
        );

    \I__4708\ : InMux
    port map (
            O => \N__19349\,
            I => \N__19330\
        );

    \I__4707\ : InMux
    port map (
            O => \N__19348\,
            I => \N__19330\
        );

    \I__4706\ : Span4Mux_v
    port map (
            O => \N__19345\,
            I => \N__19324\
        );

    \I__4705\ : Span4Mux_h
    port map (
            O => \N__19340\,
            I => \N__19324\
        );

    \I__4704\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19319\
        );

    \I__4703\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19319\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__19335\,
            I => \N__19314\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19314\
        );

    \I__4700\ : InMux
    port map (
            O => \N__19329\,
            I => \N__19309\
        );

    \I__4699\ : Span4Mux_v
    port map (
            O => \N__19324\,
            I => \N__19306\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19301\
        );

    \I__4697\ : Span12Mux_s10_h
    port map (
            O => \N__19314\,
            I => \N__19301\
        );

    \I__4696\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19296\
        );

    \I__4695\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19296\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__19309\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__19306\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4692\ : Odrv12
    port map (
            O => \N__19301\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__19296\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__4690\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19278\
        );

    \I__4689\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19275\
        );

    \I__4688\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19270\
        );

    \I__4687\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19270\
        );

    \I__4686\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19265\
        );

    \I__4685\ : InMux
    port map (
            O => \N__19282\,
            I => \N__19265\
        );

    \I__4684\ : InMux
    port map (
            O => \N__19281\,
            I => \N__19261\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__19278\,
            I => \N__19257\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19253\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__19270\,
            I => \N__19250\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19247\
        );

    \I__4679\ : CascadeMux
    port map (
            O => \N__19264\,
            I => \N__19244\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__19261\,
            I => \N__19240\
        );

    \I__4677\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19237\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__19257\,
            I => \N__19234\
        );

    \I__4675\ : InMux
    port map (
            O => \N__19256\,
            I => \N__19231\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__19253\,
            I => \N__19228\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__19250\,
            I => \N__19221\
        );

    \I__4672\ : Span4Mux_s3_v
    port map (
            O => \N__19247\,
            I => \N__19221\
        );

    \I__4671\ : InMux
    port map (
            O => \N__19244\,
            I => \N__19218\
        );

    \I__4670\ : InMux
    port map (
            O => \N__19243\,
            I => \N__19215\
        );

    \I__4669\ : Span4Mux_h
    port map (
            O => \N__19240\,
            I => \N__19212\
        );

    \I__4668\ : LocalMux
    port map (
            O => \N__19237\,
            I => \N__19203\
        );

    \I__4667\ : Span4Mux_h
    port map (
            O => \N__19234\,
            I => \N__19203\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__19231\,
            I => \N__19203\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__19228\,
            I => \N__19203\
        );

    \I__4664\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19198\
        );

    \I__4663\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19198\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__19221\,
            I => \N__19195\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__19218\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__19215\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4659\ : Odrv4
    port map (
            O => \N__19212\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__19203\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__19198\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__19195\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4655\ : CascadeMux
    port map (
            O => \N__19182\,
            I => \N__19174\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__19181\,
            I => \N__19170\
        );

    \I__4653\ : CascadeMux
    port map (
            O => \N__19180\,
            I => \N__19167\
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__19179\,
            I => \N__19164\
        );

    \I__4651\ : CascadeMux
    port map (
            O => \N__19178\,
            I => \N__19161\
        );

    \I__4650\ : CascadeMux
    port map (
            O => \N__19177\,
            I => \N__19158\
        );

    \I__4649\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19155\
        );

    \I__4648\ : InMux
    port map (
            O => \N__19173\,
            I => \N__19152\
        );

    \I__4647\ : InMux
    port map (
            O => \N__19170\,
            I => \N__19147\
        );

    \I__4646\ : InMux
    port map (
            O => \N__19167\,
            I => \N__19147\
        );

    \I__4645\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19142\
        );

    \I__4644\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19142\
        );

    \I__4643\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19137\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__19155\,
            I => \N__19133\
        );

    \I__4641\ : LocalMux
    port map (
            O => \N__19152\,
            I => \N__19130\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19125\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__19142\,
            I => \N__19125\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__19141\,
            I => \N__19122\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__19140\,
            I => \N__19119\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__19137\,
            I => \N__19116\
        );

    \I__4635\ : CascadeMux
    port map (
            O => \N__19136\,
            I => \N__19112\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__19133\,
            I => \N__19109\
        );

    \I__4633\ : Span4Mux_v
    port map (
            O => \N__19130\,
            I => \N__19104\
        );

    \I__4632\ : Span4Mux_v
    port map (
            O => \N__19125\,
            I => \N__19104\
        );

    \I__4631\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19099\
        );

    \I__4630\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19099\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__19116\,
            I => \N__19096\
        );

    \I__4628\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19091\
        );

    \I__4627\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19091\
        );

    \I__4626\ : Span4Mux_v
    port map (
            O => \N__19109\,
            I => \N__19088\
        );

    \I__4625\ : Span4Mux_h
    port map (
            O => \N__19104\,
            I => \N__19083\
        );

    \I__4624\ : LocalMux
    port map (
            O => \N__19099\,
            I => \N__19083\
        );

    \I__4623\ : Odrv4
    port map (
            O => \N__19096\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__19091\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__4621\ : Odrv4
    port map (
            O => \N__19088\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__4620\ : Odrv4
    port map (
            O => \N__19083\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__4619\ : InMux
    port map (
            O => \N__19074\,
            I => \N__19065\
        );

    \I__4618\ : InMux
    port map (
            O => \N__19073\,
            I => \N__19060\
        );

    \I__4617\ : InMux
    port map (
            O => \N__19072\,
            I => \N__19060\
        );

    \I__4616\ : InMux
    port map (
            O => \N__19071\,
            I => \N__19055\
        );

    \I__4615\ : InMux
    port map (
            O => \N__19070\,
            I => \N__19055\
        );

    \I__4614\ : InMux
    port map (
            O => \N__19069\,
            I => \N__19048\
        );

    \I__4613\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19048\
        );

    \I__4612\ : LocalMux
    port map (
            O => \N__19065\,
            I => \N__19045\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__19060\,
            I => \N__19040\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__19055\,
            I => \N__19040\
        );

    \I__4609\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19032\
        );

    \I__4608\ : InMux
    port map (
            O => \N__19053\,
            I => \N__19032\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__19029\
        );

    \I__4606\ : Span4Mux_s3_v
    port map (
            O => \N__19045\,
            I => \N__19026\
        );

    \I__4605\ : Span4Mux_s3_v
    port map (
            O => \N__19040\,
            I => \N__19021\
        );

    \I__4604\ : InMux
    port map (
            O => \N__19039\,
            I => \N__19014\
        );

    \I__4603\ : InMux
    port map (
            O => \N__19038\,
            I => \N__19014\
        );

    \I__4602\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19014\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__19032\,
            I => \N__19011\
        );

    \I__4600\ : Span4Mux_v
    port map (
            O => \N__19029\,
            I => \N__19006\
        );

    \I__4599\ : Span4Mux_v
    port map (
            O => \N__19026\,
            I => \N__19006\
        );

    \I__4598\ : InMux
    port map (
            O => \N__19025\,
            I => \N__19001\
        );

    \I__4597\ : InMux
    port map (
            O => \N__19024\,
            I => \N__19001\
        );

    \I__4596\ : Span4Mux_h
    port map (
            O => \N__19021\,
            I => \N__18998\
        );

    \I__4595\ : LocalMux
    port map (
            O => \N__19014\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__19011\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__19006\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__19001\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__4591\ : Odrv4
    port map (
            O => \N__18998\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__4590\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18984\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__18984\,
            I => \N__18980\
        );

    \I__4588\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18977\
        );

    \I__4587\ : Span12Mux_s1_h
    port map (
            O => \N__18980\,
            I => \N__18972\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__18977\,
            I => \N__18972\
        );

    \I__4585\ : Odrv12
    port map (
            O => \N__18972\,
            I => \Lab_UT.dictrl.dicRun_2\
        );

    \I__4584\ : InMux
    port map (
            O => \N__18969\,
            I => \N__18964\
        );

    \I__4583\ : InMux
    port map (
            O => \N__18968\,
            I => \N__18961\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__18967\,
            I => \N__18956\
        );

    \I__4581\ : LocalMux
    port map (
            O => \N__18964\,
            I => \N__18949\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18946\
        );

    \I__4579\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18943\
        );

    \I__4578\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18938\
        );

    \I__4577\ : InMux
    port map (
            O => \N__18956\,
            I => \N__18938\
        );

    \I__4576\ : InMux
    port map (
            O => \N__18955\,
            I => \N__18933\
        );

    \I__4575\ : InMux
    port map (
            O => \N__18954\,
            I => \N__18933\
        );

    \I__4574\ : InMux
    port map (
            O => \N__18953\,
            I => \N__18928\
        );

    \I__4573\ : InMux
    port map (
            O => \N__18952\,
            I => \N__18928\
        );

    \I__4572\ : Span4Mux_h
    port map (
            O => \N__18949\,
            I => \N__18925\
        );

    \I__4571\ : Span4Mux_h
    port map (
            O => \N__18946\,
            I => \N__18918\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__18943\,
            I => \N__18918\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__18938\,
            I => \N__18918\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__18933\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__18928\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__18925\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4565\ : Odrv4
    port map (
            O => \N__18918\,
            I => \Lab_UT.state_i_3_2\
        );

    \I__4564\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18905\
        );

    \I__4563\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18897\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__18905\,
            I => \N__18890\
        );

    \I__4561\ : InMux
    port map (
            O => \N__18904\,
            I => \N__18887\
        );

    \I__4560\ : InMux
    port map (
            O => \N__18903\,
            I => \N__18878\
        );

    \I__4559\ : InMux
    port map (
            O => \N__18902\,
            I => \N__18878\
        );

    \I__4558\ : InMux
    port map (
            O => \N__18901\,
            I => \N__18878\
        );

    \I__4557\ : InMux
    port map (
            O => \N__18900\,
            I => \N__18878\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__18897\,
            I => \N__18874\
        );

    \I__4555\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18865\
        );

    \I__4554\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18865\
        );

    \I__4553\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18865\
        );

    \I__4552\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18865\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__18890\,
            I => \N__18858\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__18887\,
            I => \N__18858\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__18878\,
            I => \N__18858\
        );

    \I__4548\ : InMux
    port map (
            O => \N__18877\,
            I => \N__18855\
        );

    \I__4547\ : Odrv4
    port map (
            O => \N__18874\,
            I => \Lab_UT.state_0\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__18865\,
            I => \Lab_UT.state_0\
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__18858\,
            I => \Lab_UT.state_0\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__18855\,
            I => \Lab_UT.state_0\
        );

    \I__4543\ : InMux
    port map (
            O => \N__18846\,
            I => \N__18836\
        );

    \I__4542\ : InMux
    port map (
            O => \N__18845\,
            I => \N__18836\
        );

    \I__4541\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18836\
        );

    \I__4540\ : InMux
    port map (
            O => \N__18843\,
            I => \N__18833\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__18836\,
            I => \N__18830\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__18833\,
            I => \N__18827\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__18830\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__4536\ : Odrv4
    port map (
            O => \N__18827\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__4535\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18819\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__18819\,
            I => \N__18816\
        );

    \I__4533\ : Span4Mux_h
    port map (
            O => \N__18816\,
            I => \N__18811\
        );

    \I__4532\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18808\
        );

    \I__4531\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18805\
        );

    \I__4530\ : Odrv4
    port map (
            O => \N__18811\,
            I => \Lab_UT.nine\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__18808\,
            I => \Lab_UT.nine\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__18805\,
            I => \Lab_UT.nine\
        );

    \I__4527\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18788\
        );

    \I__4526\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18788\
        );

    \I__4525\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18788\
        );

    \I__4524\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18785\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__18788\,
            I => \N__18782\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__18785\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__18782\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__4520\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18772\
        );

    \I__4519\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18767\
        );

    \I__4518\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18767\
        );

    \I__4517\ : LocalMux
    port map (
            O => \N__18772\,
            I => \N__18761\
        );

    \I__4516\ : LocalMux
    port map (
            O => \N__18767\,
            I => \N__18761\
        );

    \I__4515\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18758\
        );

    \I__4514\ : Span4Mux_h
    port map (
            O => \N__18761\,
            I => \N__18755\
        );

    \I__4513\ : LocalMux
    port map (
            O => \N__18758\,
            I => \Lab_UT.q_RNI84NN1_2\
        );

    \I__4512\ : Odrv4
    port map (
            O => \N__18755\,
            I => \Lab_UT.q_RNI84NN1_2\
        );

    \I__4511\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18738\
        );

    \I__4510\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18735\
        );

    \I__4509\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18732\
        );

    \I__4508\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18729\
        );

    \I__4507\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18726\
        );

    \I__4506\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18719\
        );

    \I__4505\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18719\
        );

    \I__4504\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18719\
        );

    \I__4503\ : SRMux
    port map (
            O => \N__18742\,
            I => \N__18714\
        );

    \I__4502\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18714\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__18738\,
            I => \N__18684\
        );

    \I__4500\ : LocalMux
    port map (
            O => \N__18735\,
            I => \N__18681\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__18732\,
            I => \N__18678\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__18729\,
            I => \N__18675\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18672\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18669\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__18714\,
            I => \N__18645\
        );

    \I__4494\ : SRMux
    port map (
            O => \N__18713\,
            I => \N__18534\
        );

    \I__4493\ : SRMux
    port map (
            O => \N__18712\,
            I => \N__18534\
        );

    \I__4492\ : SRMux
    port map (
            O => \N__18711\,
            I => \N__18534\
        );

    \I__4491\ : SRMux
    port map (
            O => \N__18710\,
            I => \N__18534\
        );

    \I__4490\ : SRMux
    port map (
            O => \N__18709\,
            I => \N__18534\
        );

    \I__4489\ : SRMux
    port map (
            O => \N__18708\,
            I => \N__18534\
        );

    \I__4488\ : SRMux
    port map (
            O => \N__18707\,
            I => \N__18534\
        );

    \I__4487\ : SRMux
    port map (
            O => \N__18706\,
            I => \N__18534\
        );

    \I__4486\ : SRMux
    port map (
            O => \N__18705\,
            I => \N__18534\
        );

    \I__4485\ : SRMux
    port map (
            O => \N__18704\,
            I => \N__18534\
        );

    \I__4484\ : SRMux
    port map (
            O => \N__18703\,
            I => \N__18534\
        );

    \I__4483\ : SRMux
    port map (
            O => \N__18702\,
            I => \N__18534\
        );

    \I__4482\ : SRMux
    port map (
            O => \N__18701\,
            I => \N__18534\
        );

    \I__4481\ : SRMux
    port map (
            O => \N__18700\,
            I => \N__18534\
        );

    \I__4480\ : SRMux
    port map (
            O => \N__18699\,
            I => \N__18534\
        );

    \I__4479\ : SRMux
    port map (
            O => \N__18698\,
            I => \N__18534\
        );

    \I__4478\ : SRMux
    port map (
            O => \N__18697\,
            I => \N__18534\
        );

    \I__4477\ : SRMux
    port map (
            O => \N__18696\,
            I => \N__18534\
        );

    \I__4476\ : SRMux
    port map (
            O => \N__18695\,
            I => \N__18534\
        );

    \I__4475\ : SRMux
    port map (
            O => \N__18694\,
            I => \N__18534\
        );

    \I__4474\ : SRMux
    port map (
            O => \N__18693\,
            I => \N__18534\
        );

    \I__4473\ : SRMux
    port map (
            O => \N__18692\,
            I => \N__18534\
        );

    \I__4472\ : SRMux
    port map (
            O => \N__18691\,
            I => \N__18534\
        );

    \I__4471\ : SRMux
    port map (
            O => \N__18690\,
            I => \N__18534\
        );

    \I__4470\ : SRMux
    port map (
            O => \N__18689\,
            I => \N__18534\
        );

    \I__4469\ : SRMux
    port map (
            O => \N__18688\,
            I => \N__18534\
        );

    \I__4468\ : SRMux
    port map (
            O => \N__18687\,
            I => \N__18534\
        );

    \I__4467\ : Glb2LocalMux
    port map (
            O => \N__18684\,
            I => \N__18534\
        );

    \I__4466\ : Glb2LocalMux
    port map (
            O => \N__18681\,
            I => \N__18534\
        );

    \I__4465\ : Glb2LocalMux
    port map (
            O => \N__18678\,
            I => \N__18534\
        );

    \I__4464\ : Glb2LocalMux
    port map (
            O => \N__18675\,
            I => \N__18534\
        );

    \I__4463\ : Glb2LocalMux
    port map (
            O => \N__18672\,
            I => \N__18534\
        );

    \I__4462\ : Glb2LocalMux
    port map (
            O => \N__18669\,
            I => \N__18534\
        );

    \I__4461\ : SRMux
    port map (
            O => \N__18668\,
            I => \N__18534\
        );

    \I__4460\ : SRMux
    port map (
            O => \N__18667\,
            I => \N__18534\
        );

    \I__4459\ : SRMux
    port map (
            O => \N__18666\,
            I => \N__18534\
        );

    \I__4458\ : SRMux
    port map (
            O => \N__18665\,
            I => \N__18534\
        );

    \I__4457\ : SRMux
    port map (
            O => \N__18664\,
            I => \N__18534\
        );

    \I__4456\ : SRMux
    port map (
            O => \N__18663\,
            I => \N__18534\
        );

    \I__4455\ : SRMux
    port map (
            O => \N__18662\,
            I => \N__18534\
        );

    \I__4454\ : SRMux
    port map (
            O => \N__18661\,
            I => \N__18534\
        );

    \I__4453\ : SRMux
    port map (
            O => \N__18660\,
            I => \N__18534\
        );

    \I__4452\ : SRMux
    port map (
            O => \N__18659\,
            I => \N__18534\
        );

    \I__4451\ : SRMux
    port map (
            O => \N__18658\,
            I => \N__18534\
        );

    \I__4450\ : SRMux
    port map (
            O => \N__18657\,
            I => \N__18534\
        );

    \I__4449\ : SRMux
    port map (
            O => \N__18656\,
            I => \N__18534\
        );

    \I__4448\ : SRMux
    port map (
            O => \N__18655\,
            I => \N__18534\
        );

    \I__4447\ : SRMux
    port map (
            O => \N__18654\,
            I => \N__18534\
        );

    \I__4446\ : SRMux
    port map (
            O => \N__18653\,
            I => \N__18534\
        );

    \I__4445\ : SRMux
    port map (
            O => \N__18652\,
            I => \N__18534\
        );

    \I__4444\ : SRMux
    port map (
            O => \N__18651\,
            I => \N__18534\
        );

    \I__4443\ : SRMux
    port map (
            O => \N__18650\,
            I => \N__18534\
        );

    \I__4442\ : SRMux
    port map (
            O => \N__18649\,
            I => \N__18534\
        );

    \I__4441\ : SRMux
    port map (
            O => \N__18648\,
            I => \N__18534\
        );

    \I__4440\ : Glb2LocalMux
    port map (
            O => \N__18645\,
            I => \N__18534\
        );

    \I__4439\ : GlobalMux
    port map (
            O => \N__18534\,
            I => \N__18531\
        );

    \I__4438\ : gio2CtrlBuf
    port map (
            O => \N__18531\,
            I => rst_g
        );

    \I__4437\ : CascadeMux
    port map (
            O => \N__18528\,
            I => \N__18523\
        );

    \I__4436\ : InMux
    port map (
            O => \N__18527\,
            I => \N__18517\
        );

    \I__4435\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18517\
        );

    \I__4434\ : InMux
    port map (
            O => \N__18523\,
            I => \N__18512\
        );

    \I__4433\ : InMux
    port map (
            O => \N__18522\,
            I => \N__18512\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__18517\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__18512\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__4430\ : ClkMux
    port map (
            O => \N__18507\,
            I => \N__18252\
        );

    \I__4429\ : ClkMux
    port map (
            O => \N__18506\,
            I => \N__18252\
        );

    \I__4428\ : ClkMux
    port map (
            O => \N__18505\,
            I => \N__18252\
        );

    \I__4427\ : ClkMux
    port map (
            O => \N__18504\,
            I => \N__18252\
        );

    \I__4426\ : ClkMux
    port map (
            O => \N__18503\,
            I => \N__18252\
        );

    \I__4425\ : ClkMux
    port map (
            O => \N__18502\,
            I => \N__18252\
        );

    \I__4424\ : ClkMux
    port map (
            O => \N__18501\,
            I => \N__18252\
        );

    \I__4423\ : ClkMux
    port map (
            O => \N__18500\,
            I => \N__18252\
        );

    \I__4422\ : ClkMux
    port map (
            O => \N__18499\,
            I => \N__18252\
        );

    \I__4421\ : ClkMux
    port map (
            O => \N__18498\,
            I => \N__18252\
        );

    \I__4420\ : ClkMux
    port map (
            O => \N__18497\,
            I => \N__18252\
        );

    \I__4419\ : ClkMux
    port map (
            O => \N__18496\,
            I => \N__18252\
        );

    \I__4418\ : ClkMux
    port map (
            O => \N__18495\,
            I => \N__18252\
        );

    \I__4417\ : ClkMux
    port map (
            O => \N__18494\,
            I => \N__18252\
        );

    \I__4416\ : ClkMux
    port map (
            O => \N__18493\,
            I => \N__18252\
        );

    \I__4415\ : ClkMux
    port map (
            O => \N__18492\,
            I => \N__18252\
        );

    \I__4414\ : ClkMux
    port map (
            O => \N__18491\,
            I => \N__18252\
        );

    \I__4413\ : ClkMux
    port map (
            O => \N__18490\,
            I => \N__18252\
        );

    \I__4412\ : ClkMux
    port map (
            O => \N__18489\,
            I => \N__18252\
        );

    \I__4411\ : ClkMux
    port map (
            O => \N__18488\,
            I => \N__18252\
        );

    \I__4410\ : ClkMux
    port map (
            O => \N__18487\,
            I => \N__18252\
        );

    \I__4409\ : ClkMux
    port map (
            O => \N__18486\,
            I => \N__18252\
        );

    \I__4408\ : ClkMux
    port map (
            O => \N__18485\,
            I => \N__18252\
        );

    \I__4407\ : ClkMux
    port map (
            O => \N__18484\,
            I => \N__18252\
        );

    \I__4406\ : ClkMux
    port map (
            O => \N__18483\,
            I => \N__18252\
        );

    \I__4405\ : ClkMux
    port map (
            O => \N__18482\,
            I => \N__18252\
        );

    \I__4404\ : ClkMux
    port map (
            O => \N__18481\,
            I => \N__18252\
        );

    \I__4403\ : ClkMux
    port map (
            O => \N__18480\,
            I => \N__18252\
        );

    \I__4402\ : ClkMux
    port map (
            O => \N__18479\,
            I => \N__18252\
        );

    \I__4401\ : ClkMux
    port map (
            O => \N__18478\,
            I => \N__18252\
        );

    \I__4400\ : ClkMux
    port map (
            O => \N__18477\,
            I => \N__18252\
        );

    \I__4399\ : ClkMux
    port map (
            O => \N__18476\,
            I => \N__18252\
        );

    \I__4398\ : ClkMux
    port map (
            O => \N__18475\,
            I => \N__18252\
        );

    \I__4397\ : ClkMux
    port map (
            O => \N__18474\,
            I => \N__18252\
        );

    \I__4396\ : ClkMux
    port map (
            O => \N__18473\,
            I => \N__18252\
        );

    \I__4395\ : ClkMux
    port map (
            O => \N__18472\,
            I => \N__18252\
        );

    \I__4394\ : ClkMux
    port map (
            O => \N__18471\,
            I => \N__18252\
        );

    \I__4393\ : ClkMux
    port map (
            O => \N__18470\,
            I => \N__18252\
        );

    \I__4392\ : ClkMux
    port map (
            O => \N__18469\,
            I => \N__18252\
        );

    \I__4391\ : ClkMux
    port map (
            O => \N__18468\,
            I => \N__18252\
        );

    \I__4390\ : ClkMux
    port map (
            O => \N__18467\,
            I => \N__18252\
        );

    \I__4389\ : ClkMux
    port map (
            O => \N__18466\,
            I => \N__18252\
        );

    \I__4388\ : ClkMux
    port map (
            O => \N__18465\,
            I => \N__18252\
        );

    \I__4387\ : ClkMux
    port map (
            O => \N__18464\,
            I => \N__18252\
        );

    \I__4386\ : ClkMux
    port map (
            O => \N__18463\,
            I => \N__18252\
        );

    \I__4385\ : ClkMux
    port map (
            O => \N__18462\,
            I => \N__18252\
        );

    \I__4384\ : ClkMux
    port map (
            O => \N__18461\,
            I => \N__18252\
        );

    \I__4383\ : ClkMux
    port map (
            O => \N__18460\,
            I => \N__18252\
        );

    \I__4382\ : ClkMux
    port map (
            O => \N__18459\,
            I => \N__18252\
        );

    \I__4381\ : ClkMux
    port map (
            O => \N__18458\,
            I => \N__18252\
        );

    \I__4380\ : ClkMux
    port map (
            O => \N__18457\,
            I => \N__18252\
        );

    \I__4379\ : ClkMux
    port map (
            O => \N__18456\,
            I => \N__18252\
        );

    \I__4378\ : ClkMux
    port map (
            O => \N__18455\,
            I => \N__18252\
        );

    \I__4377\ : ClkMux
    port map (
            O => \N__18454\,
            I => \N__18252\
        );

    \I__4376\ : ClkMux
    port map (
            O => \N__18453\,
            I => \N__18252\
        );

    \I__4375\ : ClkMux
    port map (
            O => \N__18452\,
            I => \N__18252\
        );

    \I__4374\ : ClkMux
    port map (
            O => \N__18451\,
            I => \N__18252\
        );

    \I__4373\ : ClkMux
    port map (
            O => \N__18450\,
            I => \N__18252\
        );

    \I__4372\ : ClkMux
    port map (
            O => \N__18449\,
            I => \N__18252\
        );

    \I__4371\ : ClkMux
    port map (
            O => \N__18448\,
            I => \N__18252\
        );

    \I__4370\ : ClkMux
    port map (
            O => \N__18447\,
            I => \N__18252\
        );

    \I__4369\ : ClkMux
    port map (
            O => \N__18446\,
            I => \N__18252\
        );

    \I__4368\ : ClkMux
    port map (
            O => \N__18445\,
            I => \N__18252\
        );

    \I__4367\ : ClkMux
    port map (
            O => \N__18444\,
            I => \N__18252\
        );

    \I__4366\ : ClkMux
    port map (
            O => \N__18443\,
            I => \N__18252\
        );

    \I__4365\ : ClkMux
    port map (
            O => \N__18442\,
            I => \N__18252\
        );

    \I__4364\ : ClkMux
    port map (
            O => \N__18441\,
            I => \N__18252\
        );

    \I__4363\ : ClkMux
    port map (
            O => \N__18440\,
            I => \N__18252\
        );

    \I__4362\ : ClkMux
    port map (
            O => \N__18439\,
            I => \N__18252\
        );

    \I__4361\ : ClkMux
    port map (
            O => \N__18438\,
            I => \N__18252\
        );

    \I__4360\ : ClkMux
    port map (
            O => \N__18437\,
            I => \N__18252\
        );

    \I__4359\ : ClkMux
    port map (
            O => \N__18436\,
            I => \N__18252\
        );

    \I__4358\ : ClkMux
    port map (
            O => \N__18435\,
            I => \N__18252\
        );

    \I__4357\ : ClkMux
    port map (
            O => \N__18434\,
            I => \N__18252\
        );

    \I__4356\ : ClkMux
    port map (
            O => \N__18433\,
            I => \N__18252\
        );

    \I__4355\ : ClkMux
    port map (
            O => \N__18432\,
            I => \N__18252\
        );

    \I__4354\ : ClkMux
    port map (
            O => \N__18431\,
            I => \N__18252\
        );

    \I__4353\ : ClkMux
    port map (
            O => \N__18430\,
            I => \N__18252\
        );

    \I__4352\ : ClkMux
    port map (
            O => \N__18429\,
            I => \N__18252\
        );

    \I__4351\ : ClkMux
    port map (
            O => \N__18428\,
            I => \N__18252\
        );

    \I__4350\ : ClkMux
    port map (
            O => \N__18427\,
            I => \N__18252\
        );

    \I__4349\ : ClkMux
    port map (
            O => \N__18426\,
            I => \N__18252\
        );

    \I__4348\ : ClkMux
    port map (
            O => \N__18425\,
            I => \N__18252\
        );

    \I__4347\ : ClkMux
    port map (
            O => \N__18424\,
            I => \N__18252\
        );

    \I__4346\ : ClkMux
    port map (
            O => \N__18423\,
            I => \N__18252\
        );

    \I__4345\ : GlobalMux
    port map (
            O => \N__18252\,
            I => \N__18249\
        );

    \I__4344\ : gio2CtrlBuf
    port map (
            O => \N__18249\,
            I => clk_g
        );

    \I__4343\ : SRMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18239\
        );

    \I__4341\ : SRMux
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__4340\ : Span4Mux_v
    port map (
            O => \N__18239\,
            I => \N__18230\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__18236\,
            I => \N__18230\
        );

    \I__4338\ : SRMux
    port map (
            O => \N__18235\,
            I => \N__18227\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__18230\,
            I => \N__18224\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__18227\,
            I => \N__18220\
        );

    \I__4335\ : IoSpan4Mux
    port map (
            O => \N__18224\,
            I => \N__18217\
        );

    \I__4334\ : SRMux
    port map (
            O => \N__18223\,
            I => \N__18214\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__18220\,
            I => \N__18211\
        );

    \I__4332\ : Span4Mux_s2_h
    port map (
            O => \N__18217\,
            I => \N__18206\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__18214\,
            I => \N__18206\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__18211\,
            I => \N__18201\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__18206\,
            I => \N__18201\
        );

    \I__4328\ : Span4Mux_h
    port map (
            O => \N__18201\,
            I => \N__18198\
        );

    \I__4327\ : Odrv4
    port map (
            O => \N__18198\,
            I => \oneSecStrb_i\
        );

    \I__4326\ : InMux
    port map (
            O => \N__18195\,
            I => \N__18192\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__18192\,
            I => \N__18189\
        );

    \I__4324\ : Span4Mux_h
    port map (
            O => \N__18189\,
            I => \N__18186\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__18186\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_4\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__18183\,
            I => \Lab_UT.three_2_cascade_\
        );

    \I__4321\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18175\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__18179\,
            I => \N__18172\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__18178\,
            I => \N__18167\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__18175\,
            I => \N__18163\
        );

    \I__4317\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18150\
        );

    \I__4316\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18150\
        );

    \I__4315\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18150\
        );

    \I__4314\ : InMux
    port map (
            O => \N__18167\,
            I => \N__18145\
        );

    \I__4313\ : InMux
    port map (
            O => \N__18166\,
            I => \N__18145\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__18163\,
            I => \N__18142\
        );

    \I__4311\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18137\
        );

    \I__4310\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18137\
        );

    \I__4309\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18130\
        );

    \I__4308\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18130\
        );

    \I__4307\ : InMux
    port map (
            O => \N__18158\,
            I => \N__18130\
        );

    \I__4306\ : InMux
    port map (
            O => \N__18157\,
            I => \N__18127\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__18150\,
            I => \N__18122\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__18145\,
            I => \N__18122\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__18142\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__18137\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__18130\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__18127\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__4299\ : Odrv12
    port map (
            O => \N__18122\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__4298\ : CascadeMux
    port map (
            O => \N__18111\,
            I => \N__18108\
        );

    \I__4297\ : InMux
    port map (
            O => \N__18108\,
            I => \N__18105\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18102\
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__18102\,
            I => \Lab_UT.didp.countrce2.un15_ce_2\
        );

    \I__4294\ : CascadeMux
    port map (
            O => \N__18099\,
            I => \Lab_UT.didp.countrce2.un15_ce_2_cascade_\
        );

    \I__4293\ : InMux
    port map (
            O => \N__18096\,
            I => \N__18092\
        );

    \I__4292\ : InMux
    port map (
            O => \N__18095\,
            I => \N__18077\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__18092\,
            I => \N__18074\
        );

    \I__4290\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18069\
        );

    \I__4289\ : InMux
    port map (
            O => \N__18090\,
            I => \N__18069\
        );

    \I__4288\ : InMux
    port map (
            O => \N__18089\,
            I => \N__18062\
        );

    \I__4287\ : InMux
    port map (
            O => \N__18088\,
            I => \N__18062\
        );

    \I__4286\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18062\
        );

    \I__4285\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18055\
        );

    \I__4284\ : InMux
    port map (
            O => \N__18085\,
            I => \N__18055\
        );

    \I__4283\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18055\
        );

    \I__4282\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18046\
        );

    \I__4281\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18046\
        );

    \I__4280\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18046\
        );

    \I__4279\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18046\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__18077\,
            I => \N__18037\
        );

    \I__4277\ : Span12Mux_s6_h
    port map (
            O => \N__18074\,
            I => \N__18037\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__18069\,
            I => \N__18037\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__18062\,
            I => \N__18037\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__18055\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__18046\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__4272\ : Odrv12
    port map (
            O => \N__18037\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__4271\ : CascadeMux
    port map (
            O => \N__18030\,
            I => \Lab_UT.didp.countrce2.un20_qPone_cascade_\
        );

    \I__4270\ : CascadeMux
    port map (
            O => \N__18027\,
            I => \N__18022\
        );

    \I__4269\ : InMux
    port map (
            O => \N__18026\,
            I => \N__18012\
        );

    \I__4268\ : InMux
    port map (
            O => \N__18025\,
            I => \N__18007\
        );

    \I__4267\ : InMux
    port map (
            O => \N__18022\,
            I => \N__18007\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__18021\,
            I => \N__18004\
        );

    \I__4265\ : CascadeMux
    port map (
            O => \N__18020\,
            I => \N__18000\
        );

    \I__4264\ : CascadeMux
    port map (
            O => \N__18019\,
            I => \N__17997\
        );

    \I__4263\ : CascadeMux
    port map (
            O => \N__18018\,
            I => \N__17994\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__18017\,
            I => \N__17991\
        );

    \I__4261\ : InMux
    port map (
            O => \N__18016\,
            I => \N__17986\
        );

    \I__4260\ : InMux
    port map (
            O => \N__18015\,
            I => \N__17986\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__18012\,
            I => \N__17981\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__18007\,
            I => \N__17981\
        );

    \I__4257\ : InMux
    port map (
            O => \N__18004\,
            I => \N__17974\
        );

    \I__4256\ : InMux
    port map (
            O => \N__18003\,
            I => \N__17974\
        );

    \I__4255\ : InMux
    port map (
            O => \N__18000\,
            I => \N__17974\
        );

    \I__4254\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17971\
        );

    \I__4253\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17966\
        );

    \I__4252\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17966\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__17986\,
            I => \N__17961\
        );

    \I__4250\ : Span4Mux_h
    port map (
            O => \N__17981\,
            I => \N__17961\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__17974\,
            I => \N__17958\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__17971\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__17966\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__17961\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4245\ : Odrv12
    port map (
            O => \N__17958\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4244\ : InMux
    port map (
            O => \N__17949\,
            I => \N__17940\
        );

    \I__4243\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17940\
        );

    \I__4242\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17937\
        );

    \I__4241\ : InMux
    port map (
            O => \N__17946\,
            I => \N__17934\
        );

    \I__4240\ : InMux
    port map (
            O => \N__17945\,
            I => \N__17931\
        );

    \I__4239\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17928\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__17937\,
            I => \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__17934\,
            I => \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__17931\,
            I => \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\
        );

    \I__4235\ : Odrv4
    port map (
            O => \N__17928\,
            I => \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\
        );

    \I__4234\ : InMux
    port map (
            O => \N__17919\,
            I => \N__17916\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17913\
        );

    \I__4232\ : Span4Mux_h
    port map (
            O => \N__17913\,
            I => \N__17908\
        );

    \I__4231\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17905\
        );

    \I__4230\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17902\
        );

    \I__4229\ : Odrv4
    port map (
            O => \N__17908\,
            I => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__17905\,
            I => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__17902\,
            I => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1\
        );

    \I__4226\ : CascadeMux
    port map (
            O => \N__17895\,
            I => \N__17891\
        );

    \I__4225\ : CascadeMux
    port map (
            O => \N__17894\,
            I => \N__17888\
        );

    \I__4224\ : InMux
    port map (
            O => \N__17891\,
            I => \N__17881\
        );

    \I__4223\ : InMux
    port map (
            O => \N__17888\,
            I => \N__17881\
        );

    \I__4222\ : InMux
    port map (
            O => \N__17887\,
            I => \N__17878\
        );

    \I__4221\ : CascadeMux
    port map (
            O => \N__17886\,
            I => \N__17871\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__17881\,
            I => \N__17865\
        );

    \I__4219\ : LocalMux
    port map (
            O => \N__17878\,
            I => \N__17865\
        );

    \I__4218\ : InMux
    port map (
            O => \N__17877\,
            I => \N__17862\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__17876\,
            I => \N__17856\
        );

    \I__4216\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17849\
        );

    \I__4215\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17849\
        );

    \I__4214\ : InMux
    port map (
            O => \N__17871\,
            I => \N__17849\
        );

    \I__4213\ : CascadeMux
    port map (
            O => \N__17870\,
            I => \N__17846\
        );

    \I__4212\ : Span4Mux_v
    port map (
            O => \N__17865\,
            I => \N__17841\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__17862\,
            I => \N__17841\
        );

    \I__4210\ : InMux
    port map (
            O => \N__17861\,
            I => \N__17832\
        );

    \I__4209\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17832\
        );

    \I__4208\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17832\
        );

    \I__4207\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17832\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__17849\,
            I => \N__17829\
        );

    \I__4205\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17826\
        );

    \I__4204\ : Span4Mux_h
    port map (
            O => \N__17841\,
            I => \N__17823\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__17832\,
            I => \N__17816\
        );

    \I__4202\ : Span4Mux_v
    port map (
            O => \N__17829\,
            I => \N__17816\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__17826\,
            I => \N__17816\
        );

    \I__4200\ : Sp12to4
    port map (
            O => \N__17823\,
            I => \N__17813\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__17816\,
            I => \N__17810\
        );

    \I__4198\ : Odrv12
    port map (
            O => \N__17813\,
            I => \Lab_UT.dictrl.state_retZ0Z_4\
        );

    \I__4197\ : Odrv4
    port map (
            O => \N__17810\,
            I => \Lab_UT.dictrl.state_retZ0Z_4\
        );

    \I__4196\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17800\
        );

    \I__4195\ : InMux
    port map (
            O => \N__17804\,
            I => \N__17797\
        );

    \I__4194\ : InMux
    port map (
            O => \N__17803\,
            I => \N__17793\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17790\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__17797\,
            I => \N__17787\
        );

    \I__4191\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17784\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__17793\,
            I => \Lab_UT.dictrl.next_state_set_0\
        );

    \I__4189\ : Odrv4
    port map (
            O => \N__17790\,
            I => \Lab_UT.dictrl.next_state_set_0\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__17787\,
            I => \Lab_UT.dictrl.next_state_set_0\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__17784\,
            I => \Lab_UT.dictrl.next_state_set_0\
        );

    \I__4186\ : InMux
    port map (
            O => \N__17775\,
            I => \N__17770\
        );

    \I__4185\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17765\
        );

    \I__4184\ : InMux
    port map (
            O => \N__17773\,
            I => \N__17765\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__17770\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4182\ : LocalMux
    port map (
            O => \N__17765\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__4181\ : CascadeMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__4180\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17753\
        );

    \I__4179\ : InMux
    port map (
            O => \N__17756\,
            I => \N__17749\
        );

    \I__4178\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17746\
        );

    \I__4177\ : InMux
    port map (
            O => \N__17752\,
            I => \N__17743\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__17749\,
            I => \N__17736\
        );

    \I__4175\ : Span4Mux_v
    port map (
            O => \N__17746\,
            I => \N__17731\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__17743\,
            I => \N__17731\
        );

    \I__4173\ : InMux
    port map (
            O => \N__17742\,
            I => \N__17726\
        );

    \I__4172\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17726\
        );

    \I__4171\ : InMux
    port map (
            O => \N__17740\,
            I => \N__17723\
        );

    \I__4170\ : InMux
    port map (
            O => \N__17739\,
            I => \N__17720\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__17736\,
            I => bu_rx_data_3
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__17731\,
            I => bu_rx_data_3
        );

    \I__4167\ : LocalMux
    port map (
            O => \N__17726\,
            I => bu_rx_data_3
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__17723\,
            I => bu_rx_data_3
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__17720\,
            I => bu_rx_data_3
        );

    \I__4164\ : InMux
    port map (
            O => \N__17709\,
            I => \N__17705\
        );

    \I__4163\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17698\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__17705\,
            I => \N__17695\
        );

    \I__4161\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17692\
        );

    \I__4160\ : InMux
    port map (
            O => \N__17703\,
            I => \N__17687\
        );

    \I__4159\ : InMux
    port map (
            O => \N__17702\,
            I => \N__17687\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__17701\,
            I => \N__17683\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__17698\,
            I => \N__17674\
        );

    \I__4156\ : Span4Mux_h
    port map (
            O => \N__17695\,
            I => \N__17674\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17674\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__17687\,
            I => \N__17674\
        );

    \I__4153\ : InMux
    port map (
            O => \N__17686\,
            I => \N__17669\
        );

    \I__4152\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17669\
        );

    \I__4151\ : Span4Mux_v
    port map (
            O => \N__17674\,
            I => \N__17664\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__17669\,
            I => \N__17664\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__17664\,
            I => bu_rx_data_2
        );

    \I__4148\ : CEMux
    port map (
            O => \N__17661\,
            I => \N__17657\
        );

    \I__4147\ : CEMux
    port map (
            O => \N__17660\,
            I => \N__17654\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17649\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__17654\,
            I => \N__17646\
        );

    \I__4144\ : CEMux
    port map (
            O => \N__17653\,
            I => \N__17643\
        );

    \I__4143\ : CEMux
    port map (
            O => \N__17652\,
            I => \N__17640\
        );

    \I__4142\ : Span4Mux_v
    port map (
            O => \N__17649\,
            I => \N__17637\
        );

    \I__4141\ : Span4Mux_v
    port map (
            O => \N__17646\,
            I => \N__17634\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__17643\,
            I => \N__17631\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__17640\,
            I => \N__17628\
        );

    \I__4138\ : Span4Mux_h
    port map (
            O => \N__17637\,
            I => \N__17625\
        );

    \I__4137\ : Span4Mux_h
    port map (
            O => \N__17634\,
            I => \N__17622\
        );

    \I__4136\ : Span4Mux_h
    port map (
            O => \N__17631\,
            I => \N__17619\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__17628\,
            I => \N__17616\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__17625\,
            I => \buart.Z_rx.sample\
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__17622\,
            I => \buart.Z_rx.sample\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__17619\,
            I => \buart.Z_rx.sample\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__17616\,
            I => \buart.Z_rx.sample\
        );

    \I__4130\ : InMux
    port map (
            O => \N__17607\,
            I => \N__17604\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__17604\,
            I => \N__17601\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__17601\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_0\
        );

    \I__4127\ : InMux
    port map (
            O => \N__17598\,
            I => \N__17595\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__17595\,
            I => \N__17592\
        );

    \I__4125\ : Odrv4
    port map (
            O => \N__17592\,
            I => \Lab_UT.bcd2segment1.N_192\
        );

    \I__4124\ : InMux
    port map (
            O => \N__17589\,
            I => \N__17586\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__17586\,
            I => \N__17583\
        );

    \I__4122\ : Span4Mux_s3_v
    port map (
            O => \N__17583\,
            I => \N__17580\
        );

    \I__4121\ : Span4Mux_v
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__4120\ : Odrv4
    port map (
            O => \N__17577\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_5\
        );

    \I__4119\ : InMux
    port map (
            O => \N__17574\,
            I => \N__17571\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__17571\,
            I => \N__17568\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__17568\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_3\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__17565\,
            I => \N__17562\
        );

    \I__4115\ : InMux
    port map (
            O => \N__17562\,
            I => \N__17558\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__17561\,
            I => \N__17555\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__17558\,
            I => \N__17552\
        );

    \I__4112\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17549\
        );

    \I__4111\ : Span4Mux_v
    port map (
            O => \N__17552\,
            I => \N__17542\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__17549\,
            I => \N__17542\
        );

    \I__4109\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17539\
        );

    \I__4108\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17536\
        );

    \I__4107\ : Odrv4
    port map (
            O => \N__17542\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__17539\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__17536\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__4104\ : InMux
    port map (
            O => \N__17529\,
            I => \N__17526\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__17526\,
            I => \N__17522\
        );

    \I__4102\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17517\
        );

    \I__4101\ : Span4Mux_h
    port map (
            O => \N__17522\,
            I => \N__17514\
        );

    \I__4100\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17511\
        );

    \I__4099\ : InMux
    port map (
            O => \N__17520\,
            I => \N__17508\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__17517\,
            I => \N__17505\
        );

    \I__4097\ : Odrv4
    port map (
            O => \N__17514\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__17511\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__17508\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__4094\ : Odrv4
    port map (
            O => \N__17505\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__4093\ : CEMux
    port map (
            O => \N__17496\,
            I => \N__17490\
        );

    \I__4092\ : CEMux
    port map (
            O => \N__17495\,
            I => \N__17487\
        );

    \I__4091\ : CEMux
    port map (
            O => \N__17494\,
            I => \N__17484\
        );

    \I__4090\ : CEMux
    port map (
            O => \N__17493\,
            I => \N__17481\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__17490\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17487\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__17484\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__17481\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__4085\ : SRMux
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__17469\,
            I => \N__17466\
        );

    \I__4083\ : Span4Mux_h
    port map (
            O => \N__17466\,
            I => \N__17462\
        );

    \I__4082\ : InMux
    port map (
            O => \N__17465\,
            I => \N__17459\
        );

    \I__4081\ : Odrv4
    port map (
            O => \N__17462\,
            I => \Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__17459\,
            I => \Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17454\,
            I => \N__17446\
        );

    \I__4078\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17443\
        );

    \I__4077\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17436\
        );

    \I__4076\ : InMux
    port map (
            O => \N__17451\,
            I => \N__17436\
        );

    \I__4075\ : InMux
    port map (
            O => \N__17450\,
            I => \N__17436\
        );

    \I__4074\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17433\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__17446\,
            I => \N__17430\
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__17443\,
            I => \N__17425\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__17436\,
            I => \N__17425\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__17433\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__4069\ : Odrv12
    port map (
            O => \N__17430\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__17425\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__17418\,
            I => \buart.Z_rx.valid_0_cascade_\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__17415\,
            I => \N__17412\
        );

    \I__4065\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17406\
        );

    \I__4064\ : InMux
    port map (
            O => \N__17411\,
            I => \N__17399\
        );

    \I__4063\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17399\
        );

    \I__4062\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17396\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__17406\,
            I => \N__17393\
        );

    \I__4060\ : InMux
    port map (
            O => \N__17405\,
            I => \N__17390\
        );

    \I__4059\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17387\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__17399\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__17396\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__17393\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__17390\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__17387\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__17376\,
            I => \bu_rx_data_rdy_cascade_\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__17373\,
            I => \N__17369\
        );

    \I__4051\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17361\
        );

    \I__4050\ : InMux
    port map (
            O => \N__17369\,
            I => \N__17361\
        );

    \I__4049\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17358\
        );

    \I__4048\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17353\
        );

    \I__4047\ : InMux
    port map (
            O => \N__17366\,
            I => \N__17353\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__17361\,
            I => \N__17350\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__17358\,
            I => \N__17345\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__17353\,
            I => \N__17345\
        );

    \I__4043\ : Odrv12
    port map (
            O => \N__17350\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__17345\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__4041\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17334\
        );

    \I__4040\ : InMux
    port map (
            O => \N__17339\,
            I => \N__17331\
        );

    \I__4039\ : InMux
    port map (
            O => \N__17338\,
            I => \N__17326\
        );

    \I__4038\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17326\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__17334\,
            I => \N__17323\
        );

    \I__4036\ : LocalMux
    port map (
            O => \N__17331\,
            I => \N__17318\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__17326\,
            I => \N__17318\
        );

    \I__4034\ : Odrv12
    port map (
            O => \N__17323\,
            I => \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1\
        );

    \I__4033\ : Odrv4
    port map (
            O => \N__17318\,
            I => \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1\
        );

    \I__4032\ : InMux
    port map (
            O => \N__17313\,
            I => \N__17310\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17310\,
            I => \Lab_UT.dictrl.next_state_out_2\
        );

    \I__4030\ : InMux
    port map (
            O => \N__17307\,
            I => \N__17302\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__17306\,
            I => \N__17299\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__17305\,
            I => \N__17295\
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__17302\,
            I => \N__17292\
        );

    \I__4026\ : InMux
    port map (
            O => \N__17299\,
            I => \N__17289\
        );

    \I__4025\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17286\
        );

    \I__4024\ : InMux
    port map (
            O => \N__17295\,
            I => \N__17283\
        );

    \I__4023\ : Odrv4
    port map (
            O => \N__17292\,
            I => \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__17289\,
            I => \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__17286\,
            I => \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__17283\,
            I => \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__17274\,
            I => \N__17270\
        );

    \I__4018\ : CascadeMux
    port map (
            O => \N__17273\,
            I => \N__17264\
        );

    \I__4017\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17261\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17269\,
            I => \N__17258\
        );

    \I__4015\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17253\
        );

    \I__4014\ : InMux
    port map (
            O => \N__17267\,
            I => \N__17253\
        );

    \I__4013\ : InMux
    port map (
            O => \N__17264\,
            I => \N__17250\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__17261\,
            I => \N__17247\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__17258\,
            I => \N__17242\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__17253\,
            I => \N__17242\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__17250\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__4008\ : Odrv4
    port map (
            O => \N__17247\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__4007\ : Odrv12
    port map (
            O => \N__17242\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__17235\,
            I => \N__17231\
        );

    \I__4005\ : InMux
    port map (
            O => \N__17234\,
            I => \N__17224\
        );

    \I__4004\ : InMux
    port map (
            O => \N__17231\,
            I => \N__17219\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17219\
        );

    \I__4002\ : InMux
    port map (
            O => \N__17229\,
            I => \N__17214\
        );

    \I__4001\ : InMux
    port map (
            O => \N__17228\,
            I => \N__17214\
        );

    \I__4000\ : InMux
    port map (
            O => \N__17227\,
            I => \N__17211\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__17224\,
            I => \N__17204\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__17219\,
            I => \N__17204\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__17214\,
            I => \N__17204\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__17211\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__3995\ : Odrv12
    port map (
            O => \N__17204\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__17199\,
            I => \N__17193\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__17198\,
            I => \N__17190\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__17197\,
            I => \N__17187\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__17196\,
            I => \N__17183\
        );

    \I__3990\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17179\
        );

    \I__3989\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17176\
        );

    \I__3988\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17173\
        );

    \I__3987\ : InMux
    port map (
            O => \N__17186\,
            I => \N__17168\
        );

    \I__3986\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17168\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__17182\,
            I => \N__17165\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__17179\,
            I => \N__17156\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__17176\,
            I => \N__17156\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__17173\,
            I => \N__17156\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__17168\,
            I => \N__17156\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17153\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__17156\,
            I => \N__17150\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__17153\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__3977\ : Odrv4
    port map (
            O => \N__17150\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17142\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__17142\,
            I => \buart.Z_rx.idle_0\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17135\
        );

    \I__3973\ : InMux
    port map (
            O => \N__17138\,
            I => \N__17132\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__17135\,
            I => \buart.Z_rx.idle\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__17132\,
            I => \buart.Z_rx.idle\
        );

    \I__3970\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17124\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__17124\,
            I => \N__17118\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17123\,
            I => \N__17115\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17110\
        );

    \I__3966\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17110\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__17118\,
            I => \N__17105\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__17115\,
            I => \N__17105\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17110\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__17105\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__17100\,
            I => \N__17095\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17091\
        );

    \I__3959\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17088\
        );

    \I__3958\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17084\
        );

    \I__3957\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17081\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17076\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17088\,
            I => \N__17076\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17087\,
            I => \N__17073\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__17084\,
            I => \N__17066\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__17081\,
            I => \N__17066\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__17076\,
            I => \N__17066\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__17073\,
            I => \buart.Z_rx.ser_clk_3\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__17066\,
            I => \buart.Z_rx.ser_clk_3\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__17061\,
            I => \buart.Z_rx.idle_cascade_\
        );

    \I__3947\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17055\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__17055\,
            I => \N__17051\
        );

    \I__3945\ : InMux
    port map (
            O => \N__17054\,
            I => \N__17048\
        );

    \I__3944\ : Span4Mux_h
    port map (
            O => \N__17051\,
            I => \N__17045\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__17048\,
            I => bu_rx_data_rdy
        );

    \I__3942\ : Odrv4
    port map (
            O => \N__17045\,
            I => bu_rx_data_rdy
        );

    \I__3941\ : CascadeMux
    port map (
            O => \N__17040\,
            I => \N__17034\
        );

    \I__3940\ : CascadeMux
    port map (
            O => \N__17039\,
            I => \N__17031\
        );

    \I__3939\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17022\
        );

    \I__3938\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17022\
        );

    \I__3937\ : InMux
    port map (
            O => \N__17034\,
            I => \N__17022\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17031\,
            I => \N__17022\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__17022\,
            I => \N__17018\
        );

    \I__3934\ : InMux
    port map (
            O => \N__17021\,
            I => \N__17015\
        );

    \I__3933\ : Odrv12
    port map (
            O => \N__17018\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__17015\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17010\,
            I => \N__17007\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17007\,
            I => \N__17003\
        );

    \I__3929\ : InMux
    port map (
            O => \N__17006\,
            I => \N__16999\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__17003\,
            I => \N__16995\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17002\,
            I => \N__16992\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__16999\,
            I => \N__16989\
        );

    \I__3925\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16986\
        );

    \I__3924\ : Odrv4
    port map (
            O => \N__16995\,
            I => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__16992\,
            I => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\
        );

    \I__3922\ : Odrv4
    port map (
            O => \N__16989\,
            I => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__16986\,
            I => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__16977\,
            I => \N__16973\
        );

    \I__3919\ : InMux
    port map (
            O => \N__16976\,
            I => \N__16969\
        );

    \I__3918\ : InMux
    port map (
            O => \N__16973\,
            I => \N__16966\
        );

    \I__3917\ : InMux
    port map (
            O => \N__16972\,
            I => \N__16963\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__16969\,
            I => \N__16960\
        );

    \I__3915\ : LocalMux
    port map (
            O => \N__16966\,
            I => \N__16956\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__16963\,
            I => \N__16953\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__16960\,
            I => \N__16950\
        );

    \I__3912\ : InMux
    port map (
            O => \N__16959\,
            I => \N__16947\
        );

    \I__3911\ : Odrv4
    port map (
            O => \N__16956\,
            I => \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__16953\,
            I => \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\
        );

    \I__3909\ : Odrv4
    port map (
            O => \N__16950\,
            I => \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__16947\,
            I => \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\
        );

    \I__3907\ : InMux
    port map (
            O => \N__16938\,
            I => \N__16932\
        );

    \I__3906\ : InMux
    port map (
            O => \N__16937\,
            I => \N__16929\
        );

    \I__3905\ : InMux
    port map (
            O => \N__16936\,
            I => \N__16926\
        );

    \I__3904\ : InMux
    port map (
            O => \N__16935\,
            I => \N__16923\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16920\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16915\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__16926\,
            I => \N__16915\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__16923\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3899\ : Odrv4
    port map (
            O => \N__16920\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3898\ : Odrv4
    port map (
            O => \N__16915\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3897\ : InMux
    port map (
            O => \N__16908\,
            I => \N__16900\
        );

    \I__3896\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16900\
        );

    \I__3895\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16897\
        );

    \I__3894\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16894\
        );

    \I__3893\ : LocalMux
    port map (
            O => \N__16900\,
            I => \N__16890\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16885\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__16894\,
            I => \N__16885\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__16893\,
            I => \N__16879\
        );

    \I__3889\ : Span4Mux_h
    port map (
            O => \N__16890\,
            I => \N__16874\
        );

    \I__3888\ : Span4Mux_s3_v
    port map (
            O => \N__16885\,
            I => \N__16871\
        );

    \I__3887\ : InMux
    port map (
            O => \N__16884\,
            I => \N__16864\
        );

    \I__3886\ : InMux
    port map (
            O => \N__16883\,
            I => \N__16864\
        );

    \I__3885\ : InMux
    port map (
            O => \N__16882\,
            I => \N__16864\
        );

    \I__3884\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16857\
        );

    \I__3883\ : InMux
    port map (
            O => \N__16878\,
            I => \N__16857\
        );

    \I__3882\ : InMux
    port map (
            O => \N__16877\,
            I => \N__16857\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__16874\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3880\ : Odrv4
    port map (
            O => \N__16871\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__16864\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3878\ : LocalMux
    port map (
            O => \N__16857\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3877\ : InMux
    port map (
            O => \N__16848\,
            I => \N__16845\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__16845\,
            I => \N__16841\
        );

    \I__3875\ : InMux
    port map (
            O => \N__16844\,
            I => \N__16838\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__16841\,
            I => \Lab_UT.alarmcharZ0Z_1\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__16838\,
            I => \Lab_UT.alarmcharZ0Z_1\
        );

    \I__3872\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16829\
        );

    \I__3871\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16818\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__16829\,
            I => \N__16813\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__16828\,
            I => \N__16807\
        );

    \I__3868\ : InMux
    port map (
            O => \N__16827\,
            I => \N__16800\
        );

    \I__3867\ : InMux
    port map (
            O => \N__16826\,
            I => \N__16800\
        );

    \I__3866\ : InMux
    port map (
            O => \N__16825\,
            I => \N__16800\
        );

    \I__3865\ : InMux
    port map (
            O => \N__16824\,
            I => \N__16795\
        );

    \I__3864\ : InMux
    port map (
            O => \N__16823\,
            I => \N__16795\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \N__16791\
        );

    \I__3862\ : InMux
    port map (
            O => \N__16821\,
            I => \N__16787\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__16818\,
            I => \N__16784\
        );

    \I__3860\ : InMux
    port map (
            O => \N__16817\,
            I => \N__16779\
        );

    \I__3859\ : InMux
    port map (
            O => \N__16816\,
            I => \N__16779\
        );

    \I__3858\ : Span4Mux_v
    port map (
            O => \N__16813\,
            I => \N__16776\
        );

    \I__3857\ : InMux
    port map (
            O => \N__16812\,
            I => \N__16773\
        );

    \I__3856\ : InMux
    port map (
            O => \N__16811\,
            I => \N__16768\
        );

    \I__3855\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16768\
        );

    \I__3854\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16765\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__16800\,
            I => \N__16760\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__16795\,
            I => \N__16760\
        );

    \I__3851\ : InMux
    port map (
            O => \N__16794\,
            I => \N__16753\
        );

    \I__3850\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16753\
        );

    \I__3849\ : InMux
    port map (
            O => \N__16790\,
            I => \N__16753\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__16787\,
            I => \N__16750\
        );

    \I__3847\ : Span4Mux_h
    port map (
            O => \N__16784\,
            I => \N__16747\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__16779\,
            I => \Lab_UT.cnt_3\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__16776\,
            I => \Lab_UT.cnt_3\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__16773\,
            I => \Lab_UT.cnt_3\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__16768\,
            I => \Lab_UT.cnt_3\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__16765\,
            I => \Lab_UT.cnt_3\
        );

    \I__3841\ : Odrv4
    port map (
            O => \N__16760\,
            I => \Lab_UT.cnt_3\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__16753\,
            I => \Lab_UT.cnt_3\
        );

    \I__3839\ : Odrv12
    port map (
            O => \N__16750\,
            I => \Lab_UT.cnt_3\
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__16747\,
            I => \Lab_UT.cnt_3\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__16728\,
            I => \N__16725\
        );

    \I__3836\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16715\
        );

    \I__3835\ : CascadeMux
    port map (
            O => \N__16724\,
            I => \N__16712\
        );

    \I__3834\ : InMux
    port map (
            O => \N__16723\,
            I => \N__16707\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__16722\,
            I => \N__16702\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__16721\,
            I => \N__16699\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__16720\,
            I => \N__16696\
        );

    \I__3830\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16689\
        );

    \I__3829\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16689\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__16715\,
            I => \N__16686\
        );

    \I__3827\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16678\
        );

    \I__3826\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16678\
        );

    \I__3825\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16678\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__16707\,
            I => \N__16675\
        );

    \I__3823\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16668\
        );

    \I__3822\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16668\
        );

    \I__3821\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16668\
        );

    \I__3820\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16661\
        );

    \I__3819\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16661\
        );

    \I__3818\ : InMux
    port map (
            O => \N__16695\,
            I => \N__16661\
        );

    \I__3817\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16658\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__16689\,
            I => \N__16655\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__16686\,
            I => \N__16652\
        );

    \I__3814\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16649\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__16678\,
            I => \N__16640\
        );

    \I__3812\ : Sp12to4
    port map (
            O => \N__16675\,
            I => \N__16640\
        );

    \I__3811\ : LocalMux
    port map (
            O => \N__16668\,
            I => \N__16640\
        );

    \I__3810\ : LocalMux
    port map (
            O => \N__16661\,
            I => \N__16640\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__16658\,
            I => \N__16633\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__16655\,
            I => \N__16633\
        );

    \I__3807\ : Span4Mux_h
    port map (
            O => \N__16652\,
            I => \N__16633\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__16649\,
            I => \Lab_UT.cnt_1\
        );

    \I__3805\ : Odrv12
    port map (
            O => \N__16640\,
            I => \Lab_UT.cnt_1\
        );

    \I__3804\ : Odrv4
    port map (
            O => \N__16633\,
            I => \Lab_UT.cnt_1\
        );

    \I__3803\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16623\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__16623\,
            I => \N__16620\
        );

    \I__3801\ : Span4Mux_h
    port map (
            O => \N__16620\,
            I => \N__16617\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__16617\,
            I => \Lab_UT.bcd2segment1.m42_bmZ0\
        );

    \I__3799\ : IoInMux
    port map (
            O => \N__16614\,
            I => \N__16611\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__16611\,
            I => \N__16608\
        );

    \I__3797\ : IoSpan4Mux
    port map (
            O => \N__16608\,
            I => \N__16603\
        );

    \I__3796\ : SRMux
    port map (
            O => \N__16607\,
            I => \N__16600\
        );

    \I__3795\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16596\
        );

    \I__3794\ : Span4Mux_s1_v
    port map (
            O => \N__16603\,
            I => \N__16593\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__16600\,
            I => \N__16590\
        );

    \I__3792\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16587\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__16596\,
            I => \N__16584\
        );

    \I__3790\ : Span4Mux_v
    port map (
            O => \N__16593\,
            I => \N__16579\
        );

    \I__3789\ : Span4Mux_s3_h
    port map (
            O => \N__16590\,
            I => \N__16579\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__16587\,
            I => \N__16576\
        );

    \I__3787\ : Span12Mux_s6_h
    port map (
            O => \N__16584\,
            I => \N__16573\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__16579\,
            I => \N__16568\
        );

    \I__3785\ : Span4Mux_h
    port map (
            O => \N__16576\,
            I => \N__16568\
        );

    \I__3784\ : Odrv12
    port map (
            O => \N__16573\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__16568\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3782\ : InMux
    port map (
            O => \N__16563\,
            I => \N__16560\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__16560\,
            I => \N__16557\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__16557\,
            I => \buart.Z_rx.bitcount_lm_0\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__16554\,
            I => \buart.Z_rx.un1_sample_0_cascade_\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16551\,
            I => \N__16548\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__16545\,
            I => \Lab_UT.dictrl.next_state_out_3\
        );

    \I__3775\ : SRMux
    port map (
            O => \N__16542\,
            I => \N__16539\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__16539\,
            I => \N__16536\
        );

    \I__3773\ : Span4Mux_h
    port map (
            O => \N__16536\,
            I => \N__16533\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__16533\,
            I => \Lab_UT.m68_0_ns\
        );

    \I__3771\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16527\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__16527\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__3769\ : InMux
    port map (
            O => \N__16524\,
            I => \N__16521\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__16521\,
            I => \N__16518\
        );

    \I__3767\ : Odrv12
    port map (
            O => \N__16518\,
            I => \buart.Z_rx.bitcount_lm_1\
        );

    \I__3766\ : InMux
    port map (
            O => \N__16515\,
            I => \N__16506\
        );

    \I__3765\ : InMux
    port map (
            O => \N__16514\,
            I => \N__16501\
        );

    \I__3764\ : InMux
    port map (
            O => \N__16513\,
            I => \N__16501\
        );

    \I__3763\ : InMux
    port map (
            O => \N__16512\,
            I => \N__16492\
        );

    \I__3762\ : InMux
    port map (
            O => \N__16511\,
            I => \N__16492\
        );

    \I__3761\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16492\
        );

    \I__3760\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16492\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__16506\,
            I => \N__16480\
        );

    \I__3758\ : LocalMux
    port map (
            O => \N__16501\,
            I => \N__16477\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__16492\,
            I => \N__16474\
        );

    \I__3756\ : InMux
    port map (
            O => \N__16491\,
            I => \N__16469\
        );

    \I__3755\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16469\
        );

    \I__3754\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16464\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16488\,
            I => \N__16464\
        );

    \I__3752\ : InMux
    port map (
            O => \N__16487\,
            I => \N__16461\
        );

    \I__3751\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16456\
        );

    \I__3750\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16456\
        );

    \I__3749\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16451\
        );

    \I__3748\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16451\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__16480\,
            I => \N__16448\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__16477\,
            I => \N__16443\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__16474\,
            I => \N__16443\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__16469\,
            I => \N__16438\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__16464\,
            I => \N__16438\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__16461\,
            I => \buart.Z_rx.startbit\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__16456\,
            I => \buart.Z_rx.startbit\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__16451\,
            I => \buart.Z_rx.startbit\
        );

    \I__3739\ : Odrv4
    port map (
            O => \N__16448\,
            I => \buart.Z_rx.startbit\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__16443\,
            I => \buart.Z_rx.startbit\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__16438\,
            I => \buart.Z_rx.startbit\
        );

    \I__3736\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16422\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__16422\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16416\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__16416\,
            I => \N__16413\
        );

    \I__3732\ : Odrv12
    port map (
            O => \N__16413\,
            I => \buart.Z_rx.bitcount_lm_2\
        );

    \I__3731\ : CascadeMux
    port map (
            O => \N__16410\,
            I => \N__16405\
        );

    \I__3730\ : CascadeMux
    port map (
            O => \N__16409\,
            I => \N__16402\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__16408\,
            I => \N__16399\
        );

    \I__3728\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16388\
        );

    \I__3727\ : InMux
    port map (
            O => \N__16402\,
            I => \N__16388\
        );

    \I__3726\ : InMux
    port map (
            O => \N__16399\,
            I => \N__16388\
        );

    \I__3725\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16388\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16384\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16379\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__16387\,
            I => \N__16375\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__16384\,
            I => \N__16370\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__16383\,
            I => \N__16367\
        );

    \I__3719\ : CascadeMux
    port map (
            O => \N__16382\,
            I => \N__16364\
        );

    \I__3718\ : Span4Mux_s2_v
    port map (
            O => \N__16379\,
            I => \N__16357\
        );

    \I__3717\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16354\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16351\
        );

    \I__3715\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16346\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16346\
        );

    \I__3713\ : Span4Mux_h
    port map (
            O => \N__16370\,
            I => \N__16343\
        );

    \I__3712\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16336\
        );

    \I__3711\ : InMux
    port map (
            O => \N__16364\,
            I => \N__16336\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16363\,
            I => \N__16336\
        );

    \I__3709\ : InMux
    port map (
            O => \N__16362\,
            I => \N__16329\
        );

    \I__3708\ : InMux
    port map (
            O => \N__16361\,
            I => \N__16329\
        );

    \I__3707\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16329\
        );

    \I__3706\ : Span4Mux_v
    port map (
            O => \N__16357\,
            I => \N__16326\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__16354\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__16351\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__16346\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3702\ : Odrv4
    port map (
            O => \N__16343\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__16336\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__16329\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__16326\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16308\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__16308\,
            I => \N__16305\
        );

    \I__3696\ : Odrv12
    port map (
            O => \N__16305\,
            I => \Lab_UT.bcd2segment1.N_166\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16302\,
            I => \N__16299\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__16299\,
            I => \N__16296\
        );

    \I__3693\ : Span4Mux_h
    port map (
            O => \N__16296\,
            I => \N__16292\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__16295\,
            I => \N__16289\
        );

    \I__3691\ : Span4Mux_v
    port map (
            O => \N__16292\,
            I => \N__16285\
        );

    \I__3690\ : InMux
    port map (
            O => \N__16289\,
            I => \N__16280\
        );

    \I__3689\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16280\
        );

    \I__3688\ : Span4Mux_s2_h
    port map (
            O => \N__16285\,
            I => \N__16276\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16273\
        );

    \I__3686\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16270\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__16276\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__16273\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__16270\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3682\ : InMux
    port map (
            O => \N__16263\,
            I => \N__16257\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16262\,
            I => \N__16257\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__16257\,
            I => \N__16249\
        );

    \I__3679\ : InMux
    port map (
            O => \N__16256\,
            I => \N__16244\
        );

    \I__3678\ : InMux
    port map (
            O => \N__16255\,
            I => \N__16244\
        );

    \I__3677\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16238\
        );

    \I__3676\ : InMux
    port map (
            O => \N__16253\,
            I => \N__16235\
        );

    \I__3675\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16232\
        );

    \I__3674\ : Span4Mux_h
    port map (
            O => \N__16249\,
            I => \N__16226\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__16244\,
            I => \N__16223\
        );

    \I__3672\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16218\
        );

    \I__3671\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16218\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16215\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__16238\,
            I => \N__16209\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__16235\,
            I => \N__16209\
        );

    \I__3667\ : LocalMux
    port map (
            O => \N__16232\,
            I => \N__16206\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16199\
        );

    \I__3665\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16199\
        );

    \I__3664\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16199\
        );

    \I__3663\ : Span4Mux_v
    port map (
            O => \N__16226\,
            I => \N__16196\
        );

    \I__3662\ : Span4Mux_v
    port map (
            O => \N__16223\,
            I => \N__16193\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__16218\,
            I => \N__16190\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__16215\,
            I => \N__16187\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16214\,
            I => \N__16184\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__16209\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__16206\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__16199\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__16196\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__16193\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__16190\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3652\ : Odrv12
    port map (
            O => \N__16187\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__16184\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16164\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16161\
        );

    \I__3648\ : Span4Mux_h
    port map (
            O => \N__16161\,
            I => \N__16158\
        );

    \I__3647\ : Odrv4
    port map (
            O => \N__16158\,
            I => \Lab_UT.didp.countrce3.q_RNO_0Z0Z_3\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16155\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16152\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__16149\,
            I => \N__16146\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16143\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__16143\,
            I => \N__16140\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__16140\,
            I => \N__16137\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__16137\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__3639\ : InMux
    port map (
            O => \N__16134\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__3638\ : InMux
    port map (
            O => \N__16131\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16125\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__16125\,
            I => \N__16122\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__16122\,
            I => \buart.Z_rx.bitcount_lm_4\
        );

    \I__3634\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16112\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16109\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__16117\,
            I => \N__16105\
        );

    \I__3631\ : CascadeMux
    port map (
            O => \N__16116\,
            I => \N__16099\
        );

    \I__3630\ : InMux
    port map (
            O => \N__16115\,
            I => \N__16096\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__16112\,
            I => \N__16093\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__16109\,
            I => \N__16090\
        );

    \I__3627\ : InMux
    port map (
            O => \N__16108\,
            I => \N__16087\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16105\,
            I => \N__16080\
        );

    \I__3625\ : InMux
    port map (
            O => \N__16104\,
            I => \N__16080\
        );

    \I__3624\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16080\
        );

    \I__3623\ : InMux
    port map (
            O => \N__16102\,
            I => \N__16077\
        );

    \I__3622\ : InMux
    port map (
            O => \N__16099\,
            I => \N__16074\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__16096\,
            I => \N__16069\
        );

    \I__3620\ : Span4Mux_h
    port map (
            O => \N__16093\,
            I => \N__16069\
        );

    \I__3619\ : Span4Mux_h
    port map (
            O => \N__16090\,
            I => \N__16064\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__16087\,
            I => \N__16064\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__16080\,
            I => \N__16059\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__16077\,
            I => \N__16059\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__16074\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__16069\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__16064\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__3612\ : Odrv4
    port map (
            O => \N__16059\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__3611\ : CascadeMux
    port map (
            O => \N__16050\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_\
        );

    \I__3610\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16044\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__16044\,
            I => \uu2.mem0.N_294\
        );

    \I__3608\ : InMux
    port map (
            O => \N__16041\,
            I => \N__16038\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__16038\,
            I => \N__16034\
        );

    \I__3606\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16031\
        );

    \I__3605\ : Odrv4
    port map (
            O => \N__16034\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__16031\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__3603\ : InMux
    port map (
            O => \N__16026\,
            I => \N__16023\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__16023\,
            I => \uu2.mem0.N_271\
        );

    \I__3601\ : InMux
    port map (
            O => \N__16020\,
            I => \N__16017\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__16017\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_80\
        );

    \I__3599\ : InMux
    port map (
            O => \N__16014\,
            I => \N__16011\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__16011\,
            I => \N__16008\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__16008\,
            I => \N__16004\
        );

    \I__3596\ : InMux
    port map (
            O => \N__16007\,
            I => \N__16001\
        );

    \I__3595\ : Odrv4
    port map (
            O => \N__16004\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__16001\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__3593\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15987\
        );

    \I__3592\ : InMux
    port map (
            O => \N__15995\,
            I => \N__15987\
        );

    \I__3591\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15984\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__15993\,
            I => \N__15978\
        );

    \I__3589\ : InMux
    port map (
            O => \N__15992\,
            I => \N__15974\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__15987\,
            I => \N__15970\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__15984\,
            I => \N__15967\
        );

    \I__3586\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15961\
        );

    \I__3585\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15961\
        );

    \I__3584\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15954\
        );

    \I__3583\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15954\
        );

    \I__3582\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15954\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__15974\,
            I => \N__15951\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15973\,
            I => \N__15948\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__15970\,
            I => \N__15943\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__15967\,
            I => \N__15943\
        );

    \I__3577\ : InMux
    port map (
            O => \N__15966\,
            I => \N__15940\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__15961\,
            I => \N__15937\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__15954\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3574\ : Odrv4
    port map (
            O => \N__15951\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__15948\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3572\ : Odrv4
    port map (
            O => \N__15943\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15940\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3570\ : Odrv4
    port map (
            O => \N__15937\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__3569\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15921\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__15921\,
            I => \N__15918\
        );

    \I__3567\ : Span4Mux_v
    port map (
            O => \N__15918\,
            I => \N__15914\
        );

    \I__3566\ : InMux
    port map (
            O => \N__15917\,
            I => \N__15911\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__15914\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__15911\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__3563\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15903\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__15903\,
            I => \N__15900\
        );

    \I__3561\ : Span4Mux_h
    port map (
            O => \N__15900\,
            I => \N__15897\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__15897\,
            I => \uu2.mem0.N_98_0\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__15894\,
            I => \N__15890\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15893\,
            I => \N__15886\
        );

    \I__3557\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15883\
        );

    \I__3556\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15880\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__15886\,
            I => \N__15877\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__15883\,
            I => \N__15872\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__15880\,
            I => \N__15872\
        );

    \I__3552\ : Span4Mux_h
    port map (
            O => \N__15877\,
            I => \N__15869\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__15872\,
            I => \N__15865\
        );

    \I__3550\ : Span4Mux_v
    port map (
            O => \N__15869\,
            I => \N__15862\
        );

    \I__3549\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15859\
        );

    \I__3548\ : Span4Mux_h
    port map (
            O => \N__15865\,
            I => \N__15856\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__15862\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__15859\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__3545\ : Odrv4
    port map (
            O => \N__15856\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \N__15845\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__15848\,
            I => \N__15841\
        );

    \I__3542\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15836\
        );

    \I__3541\ : InMux
    port map (
            O => \N__15844\,
            I => \N__15836\
        );

    \I__3540\ : InMux
    port map (
            O => \N__15841\,
            I => \N__15831\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__15836\,
            I => \N__15828\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15825\
        );

    \I__3537\ : InMux
    port map (
            O => \N__15834\,
            I => \N__15821\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__15831\,
            I => \N__15818\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__15828\,
            I => \N__15815\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__15825\,
            I => \N__15812\
        );

    \I__3533\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15809\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__15821\,
            I => \N__15806\
        );

    \I__3531\ : Odrv4
    port map (
            O => \N__15818\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__3530\ : Odrv4
    port map (
            O => \N__15815\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__3529\ : Odrv12
    port map (
            O => \N__15812\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__15809\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__3527\ : Odrv4
    port map (
            O => \N__15806\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__3526\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15789\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15789\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__15789\,
            I => \N__15782\
        );

    \I__3523\ : InMux
    port map (
            O => \N__15788\,
            I => \N__15773\
        );

    \I__3522\ : InMux
    port map (
            O => \N__15787\,
            I => \N__15773\
        );

    \I__3521\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15773\
        );

    \I__3520\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15773\
        );

    \I__3519\ : Odrv12
    port map (
            O => \N__15782\,
            I => \uu2.trig_rd_is_det\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__15773\,
            I => \uu2.trig_rd_is_det\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15765\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15761\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__15764\,
            I => \N__15758\
        );

    \I__3514\ : Span4Mux_v
    port map (
            O => \N__15761\,
            I => \N__15755\
        );

    \I__3513\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15751\
        );

    \I__3512\ : IoSpan4Mux
    port map (
            O => \N__15755\,
            I => \N__15748\
        );

    \I__3511\ : InMux
    port map (
            O => \N__15754\,
            I => \N__15745\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__15751\,
            I => \N__15738\
        );

    \I__3509\ : Span4Mux_s0_h
    port map (
            O => \N__15748\,
            I => \N__15738\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15738\
        );

    \I__3507\ : Span4Mux_h
    port map (
            O => \N__15738\,
            I => \N__15733\
        );

    \I__3506\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15728\
        );

    \I__3505\ : InMux
    port map (
            O => \N__15736\,
            I => \N__15728\
        );

    \I__3504\ : Span4Mux_h
    port map (
            O => \N__15733\,
            I => \N__15725\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__15728\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__15725\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__15720\,
            I => \uu2.N_12_i_cascade_\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15717\,
            I => \N__15708\
        );

    \I__3499\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15701\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15701\
        );

    \I__3497\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15701\
        );

    \I__3496\ : InMux
    port map (
            O => \N__15713\,
            I => \N__15698\
        );

    \I__3495\ : InMux
    port map (
            O => \N__15712\,
            I => \N__15693\
        );

    \I__3494\ : InMux
    port map (
            O => \N__15711\,
            I => \N__15693\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__15708\,
            I => \N__15688\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__15701\,
            I => \N__15688\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__15698\,
            I => \uu2.N_67\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15693\,
            I => \uu2.N_67\
        );

    \I__3489\ : Odrv12
    port map (
            O => \N__15688\,
            I => \uu2.N_67\
        );

    \I__3488\ : InMux
    port map (
            O => \N__15681\,
            I => \N__15665\
        );

    \I__3487\ : InMux
    port map (
            O => \N__15680\,
            I => \N__15665\
        );

    \I__3486\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15665\
        );

    \I__3485\ : InMux
    port map (
            O => \N__15678\,
            I => \N__15662\
        );

    \I__3484\ : InMux
    port map (
            O => \N__15677\,
            I => \N__15659\
        );

    \I__3483\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15654\
        );

    \I__3482\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15654\
        );

    \I__3481\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15644\
        );

    \I__3480\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15644\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15672\,
            I => \N__15644\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15636\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15633\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__15659\,
            I => \N__15630\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__15654\,
            I => \N__15627\
        );

    \I__3474\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15620\
        );

    \I__3473\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15620\
        );

    \I__3472\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15620\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__15644\,
            I => \N__15617\
        );

    \I__3470\ : InMux
    port map (
            O => \N__15643\,
            I => \N__15612\
        );

    \I__3469\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15612\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15605\
        );

    \I__3467\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15605\
        );

    \I__3466\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15605\
        );

    \I__3465\ : Span4Mux_h
    port map (
            O => \N__15636\,
            I => \N__15598\
        );

    \I__3464\ : Span4Mux_h
    port map (
            O => \N__15633\,
            I => \N__15598\
        );

    \I__3463\ : Span4Mux_h
    port map (
            O => \N__15630\,
            I => \N__15598\
        );

    \I__3462\ : Span4Mux_v
    port map (
            O => \N__15627\,
            I => \N__15591\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__15620\,
            I => \N__15591\
        );

    \I__3460\ : Span4Mux_s3_h
    port map (
            O => \N__15617\,
            I => \N__15591\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__15612\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__15605\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3457\ : Odrv4
    port map (
            O => \N__15598\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__15591\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15574\
        );

    \I__3454\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15570\
        );

    \I__3453\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15567\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__15579\,
            I => \N__15564\
        );

    \I__3451\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15561\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15577\,
            I => \N__15557\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__15574\,
            I => \N__15554\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15573\,
            I => \N__15551\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__15570\,
            I => \N__15547\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__15567\,
            I => \N__15544\
        );

    \I__3445\ : InMux
    port map (
            O => \N__15564\,
            I => \N__15534\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__15561\,
            I => \N__15531\
        );

    \I__3443\ : InMux
    port map (
            O => \N__15560\,
            I => \N__15528\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__15557\,
            I => \N__15521\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__15554\,
            I => \N__15521\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__15551\,
            I => \N__15521\
        );

    \I__3439\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15518\
        );

    \I__3438\ : Span4Mux_h
    port map (
            O => \N__15547\,
            I => \N__15515\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__15544\,
            I => \N__15512\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15503\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15503\
        );

    \I__3434\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15503\
        );

    \I__3433\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15503\
        );

    \I__3432\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15496\
        );

    \I__3431\ : InMux
    port map (
            O => \N__15538\,
            I => \N__15496\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15537\,
            I => \N__15496\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__15534\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3428\ : Odrv12
    port map (
            O => \N__15531\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__15528\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3426\ : Odrv4
    port map (
            O => \N__15521\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__15518\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3424\ : Odrv4
    port map (
            O => \N__15515\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3423\ : Odrv4
    port map (
            O => \N__15512\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__15503\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__15496\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__3420\ : InMux
    port map (
            O => \N__15477\,
            I => \N__15467\
        );

    \I__3419\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15460\
        );

    \I__3418\ : InMux
    port map (
            O => \N__15475\,
            I => \N__15460\
        );

    \I__3417\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15460\
        );

    \I__3416\ : InMux
    port map (
            O => \N__15473\,
            I => \N__15453\
        );

    \I__3415\ : InMux
    port map (
            O => \N__15472\,
            I => \N__15453\
        );

    \I__3414\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15453\
        );

    \I__3413\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15448\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15445\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__15460\,
            I => \N__15442\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15439\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15434\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15451\,
            I => \N__15434\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__15448\,
            I => \N__15431\
        );

    \I__3406\ : Span4Mux_v
    port map (
            O => \N__15445\,
            I => \N__15419\
        );

    \I__3405\ : Span4Mux_s3_h
    port map (
            O => \N__15442\,
            I => \N__15419\
        );

    \I__3404\ : Span4Mux_v
    port map (
            O => \N__15439\,
            I => \N__15419\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__15434\,
            I => \N__15419\
        );

    \I__3402\ : Span4Mux_h
    port map (
            O => \N__15431\,
            I => \N__15416\
        );

    \I__3401\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15411\
        );

    \I__3400\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15411\
        );

    \I__3399\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15408\
        );

    \I__3398\ : Odrv4
    port map (
            O => \N__15419\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3397\ : Odrv4
    port map (
            O => \N__15416\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__15411\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__15408\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15393\
        );

    \I__3393\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15390\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__15397\,
            I => \N__15387\
        );

    \I__3391\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15381\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15381\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15378\
        );

    \I__3388\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15375\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__15386\,
            I => \N__15370\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__15381\,
            I => \N__15367\
        );

    \I__3385\ : Span4Mux_v
    port map (
            O => \N__15378\,
            I => \N__15364\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__15375\,
            I => \N__15361\
        );

    \I__3383\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15356\
        );

    \I__3382\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15356\
        );

    \I__3381\ : InMux
    port map (
            O => \N__15370\,
            I => \N__15353\
        );

    \I__3380\ : Span4Mux_v
    port map (
            O => \N__15367\,
            I => \N__15348\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__15364\,
            I => \N__15348\
        );

    \I__3378\ : Odrv12
    port map (
            O => \N__15361\,
            I => \uu2.N_12_i\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__15356\,
            I => \uu2.N_12_i\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__15353\,
            I => \uu2.N_12_i\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__15348\,
            I => \uu2.N_12_i\
        );

    \I__3374\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15336\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__15336\,
            I => \N__15325\
        );

    \I__3372\ : InMux
    port map (
            O => \N__15335\,
            I => \N__15322\
        );

    \I__3371\ : InMux
    port map (
            O => \N__15334\,
            I => \N__15317\
        );

    \I__3370\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15317\
        );

    \I__3369\ : InMux
    port map (
            O => \N__15332\,
            I => \N__15314\
        );

    \I__3368\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15306\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15303\
        );

    \I__3366\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15300\
        );

    \I__3365\ : InMux
    port map (
            O => \N__15328\,
            I => \N__15297\
        );

    \I__3364\ : Span4Mux_h
    port map (
            O => \N__15325\,
            I => \N__15292\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__15322\,
            I => \N__15292\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__15317\,
            I => \N__15287\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__15314\,
            I => \N__15287\
        );

    \I__3360\ : InMux
    port map (
            O => \N__15313\,
            I => \N__15284\
        );

    \I__3359\ : CascadeMux
    port map (
            O => \N__15312\,
            I => \N__15278\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__15311\,
            I => \N__15275\
        );

    \I__3357\ : InMux
    port map (
            O => \N__15310\,
            I => \N__15270\
        );

    \I__3356\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15267\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__15306\,
            I => \N__15262\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15262\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__15300\,
            I => \N__15256\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__15297\,
            I => \N__15253\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__15292\,
            I => \N__15250\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__15287\,
            I => \N__15245\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__15284\,
            I => \N__15245\
        );

    \I__3348\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15232\
        );

    \I__3347\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15232\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15232\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15278\,
            I => \N__15232\
        );

    \I__3344\ : InMux
    port map (
            O => \N__15275\,
            I => \N__15232\
        );

    \I__3343\ : InMux
    port map (
            O => \N__15274\,
            I => \N__15232\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15229\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__15270\,
            I => \N__15222\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__15267\,
            I => \N__15222\
        );

    \I__3339\ : Span4Mux_h
    port map (
            O => \N__15262\,
            I => \N__15222\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15215\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15215\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15259\,
            I => \N__15215\
        );

    \I__3335\ : Odrv4
    port map (
            O => \N__15256\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3334\ : Odrv4
    port map (
            O => \N__15253\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3333\ : Odrv4
    port map (
            O => \N__15250\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3332\ : Odrv4
    port map (
            O => \N__15245\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__15232\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__15229\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3329\ : Odrv4
    port map (
            O => \N__15222\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__15215\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__3327\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15193\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15197\,
            I => \N__15184\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__15196\,
            I => \N__15180\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__15193\,
            I => \N__15176\
        );

    \I__3323\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15173\
        );

    \I__3322\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15170\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__15190\,
            I => \N__15167\
        );

    \I__3320\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15162\
        );

    \I__3319\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15162\
        );

    \I__3318\ : InMux
    port map (
            O => \N__15187\,
            I => \N__15159\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__15184\,
            I => \N__15153\
        );

    \I__3316\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15150\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15180\,
            I => \N__15144\
        );

    \I__3314\ : InMux
    port map (
            O => \N__15179\,
            I => \N__15144\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__15176\,
            I => \N__15139\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15139\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15170\,
            I => \N__15136\
        );

    \I__3310\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15133\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__15162\,
            I => \N__15128\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__15159\,
            I => \N__15128\
        );

    \I__3307\ : CascadeMux
    port map (
            O => \N__15158\,
            I => \N__15125\
        );

    \I__3306\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15119\
        );

    \I__3305\ : InMux
    port map (
            O => \N__15156\,
            I => \N__15119\
        );

    \I__3304\ : Span4Mux_h
    port map (
            O => \N__15153\,
            I => \N__15114\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__15150\,
            I => \N__15114\
        );

    \I__3302\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15107\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__15144\,
            I => \N__15104\
        );

    \I__3300\ : Span4Mux_h
    port map (
            O => \N__15139\,
            I => \N__15101\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__15136\,
            I => \N__15098\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__15133\,
            I => \N__15093\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__15128\,
            I => \N__15093\
        );

    \I__3296\ : InMux
    port map (
            O => \N__15125\,
            I => \N__15090\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15124\,
            I => \N__15087\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__15119\,
            I => \N__15082\
        );

    \I__3293\ : Span4Mux_h
    port map (
            O => \N__15114\,
            I => \N__15082\
        );

    \I__3292\ : InMux
    port map (
            O => \N__15113\,
            I => \N__15073\
        );

    \I__3291\ : InMux
    port map (
            O => \N__15112\,
            I => \N__15073\
        );

    \I__3290\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15073\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15073\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15107\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3287\ : Odrv4
    port map (
            O => \N__15104\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3286\ : Odrv4
    port map (
            O => \N__15101\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__15098\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__15093\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__15090\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__15087\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3281\ : Odrv4
    port map (
            O => \N__15082\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__15073\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__3279\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15045\
        );

    \I__3278\ : InMux
    port map (
            O => \N__15053\,
            I => \N__15045\
        );

    \I__3277\ : InMux
    port map (
            O => \N__15052\,
            I => \N__15040\
        );

    \I__3276\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15035\
        );

    \I__3275\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15035\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__15045\,
            I => \N__15032\
        );

    \I__3273\ : InMux
    port map (
            O => \N__15044\,
            I => \N__15029\
        );

    \I__3272\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15026\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__15040\,
            I => \N__15023\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__15035\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__15032\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__15029\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15026\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3266\ : Odrv12
    port map (
            O => \N__15023\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__3265\ : CascadeMux
    port map (
            O => \N__15012\,
            I => \uu2.N_272_cascade_\
        );

    \I__3264\ : InMux
    port map (
            O => \N__15009\,
            I => \N__15006\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15006\,
            I => \uu2.mem0.m317_0_a6_1_0\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15003\,
            I => \N__15000\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__15000\,
            I => \uu2.mem0.N_13\
        );

    \I__3260\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14994\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__14994\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__3258\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14967\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14967\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14989\,
            I => \N__14967\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14988\,
            I => \N__14960\
        );

    \I__3254\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14960\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14960\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14953\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14953\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14953\
        );

    \I__3249\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14942\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14942\
        );

    \I__3247\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14937\
        );

    \I__3246\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14937\
        );

    \I__3245\ : InMux
    port map (
            O => \N__14978\,
            I => \N__14927\
        );

    \I__3244\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14927\
        );

    \I__3243\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14927\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14922\
        );

    \I__3241\ : InMux
    port map (
            O => \N__14974\,
            I => \N__14922\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14967\,
            I => \N__14919\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__14960\,
            I => \N__14914\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__14953\,
            I => \N__14914\
        );

    \I__3237\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14903\
        );

    \I__3236\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14903\
        );

    \I__3235\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14903\
        );

    \I__3234\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14903\
        );

    \I__3233\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14903\
        );

    \I__3232\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14897\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__14942\,
            I => \N__14892\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__14937\,
            I => \N__14892\
        );

    \I__3229\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14887\
        );

    \I__3228\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14887\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__14934\,
            I => \N__14883\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__14927\,
            I => \N__14878\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__14922\,
            I => \N__14878\
        );

    \I__3224\ : Span4Mux_s3_v
    port map (
            O => \N__14919\,
            I => \N__14873\
        );

    \I__3223\ : Span4Mux_h
    port map (
            O => \N__14914\,
            I => \N__14873\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__14903\,
            I => \N__14870\
        );

    \I__3221\ : InMux
    port map (
            O => \N__14902\,
            I => \N__14863\
        );

    \I__3220\ : InMux
    port map (
            O => \N__14901\,
            I => \N__14863\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14900\,
            I => \N__14863\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__14897\,
            I => \N__14860\
        );

    \I__3217\ : Span4Mux_v
    port map (
            O => \N__14892\,
            I => \N__14855\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__14887\,
            I => \N__14855\
        );

    \I__3215\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14850\
        );

    \I__3214\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14850\
        );

    \I__3213\ : Span12Mux_s10_v
    port map (
            O => \N__14878\,
            I => \N__14847\
        );

    \I__3212\ : Span4Mux_v
    port map (
            O => \N__14873\,
            I => \N__14840\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__14870\,
            I => \N__14840\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__14863\,
            I => \N__14840\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__14860\,
            I => \N__14837\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__14855\,
            I => \N__14832\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__14850\,
            I => \N__14832\
        );

    \I__3206\ : Odrv12
    port map (
            O => \N__14847\,
            I => \Lab_UT.Run\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__14840\,
            I => \Lab_UT.Run\
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__14837\,
            I => \Lab_UT.Run\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__14832\,
            I => \Lab_UT.Run\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14820\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__14820\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__3200\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14811\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14811\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__3197\ : Odrv12
    port map (
            O => \N__14808\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__14805\,
            I => \N__14799\
        );

    \I__3195\ : InMux
    port map (
            O => \N__14804\,
            I => \N__14794\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14794\
        );

    \I__3193\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14790\
        );

    \I__3192\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14787\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__14794\,
            I => \N__14781\
        );

    \I__3190\ : InMux
    port map (
            O => \N__14793\,
            I => \N__14778\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__14790\,
            I => \N__14775\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__14787\,
            I => \N__14772\
        );

    \I__3187\ : InMux
    port map (
            O => \N__14786\,
            I => \N__14769\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14785\,
            I => \N__14766\
        );

    \I__3185\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14763\
        );

    \I__3184\ : Span4Mux_h
    port map (
            O => \N__14781\,
            I => \N__14758\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__14778\,
            I => \N__14758\
        );

    \I__3182\ : Span4Mux_v
    port map (
            O => \N__14775\,
            I => \N__14753\
        );

    \I__3181\ : Span4Mux_v
    port map (
            O => \N__14772\,
            I => \N__14753\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__14769\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__14766\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__14763\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__14758\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__14753\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__3175\ : InMux
    port map (
            O => \N__14742\,
            I => \N__14739\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__14739\,
            I => \uu2.N_272\
        );

    \I__3173\ : InMux
    port map (
            O => \N__14736\,
            I => \N__14733\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__14733\,
            I => \N__14728\
        );

    \I__3171\ : InMux
    port map (
            O => \N__14732\,
            I => \N__14725\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14731\,
            I => \N__14722\
        );

    \I__3169\ : Span4Mux_v
    port map (
            O => \N__14728\,
            I => \N__14717\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__14725\,
            I => \N__14717\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14722\,
            I => \N__14714\
        );

    \I__3166\ : Span4Mux_h
    port map (
            O => \N__14717\,
            I => \N__14711\
        );

    \I__3165\ : Span12Mux_s10_h
    port map (
            O => \N__14714\,
            I => \N__14708\
        );

    \I__3164\ : Span4Mux_s2_h
    port map (
            O => \N__14711\,
            I => \N__14705\
        );

    \I__3163\ : Odrv12
    port map (
            O => \N__14708\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__3162\ : Odrv4
    port map (
            O => \N__14705\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__14700\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_\
        );

    \I__3160\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14694\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__14694\,
            I => \uu2.mem0.bitmap_pmux_u_i_4_0\
        );

    \I__3158\ : InMux
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__14688\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_69\
        );

    \I__3156\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14677\
        );

    \I__3155\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14677\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__14683\,
            I => \N__14674\
        );

    \I__3153\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14671\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14665\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14662\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__14671\,
            I => \N__14659\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__14670\,
            I => \N__14656\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__14669\,
            I => \N__14653\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14646\
        );

    \I__3146\ : Span4Mux_v
    port map (
            O => \N__14665\,
            I => \N__14641\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__14662\,
            I => \N__14641\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__14659\,
            I => \N__14638\
        );

    \I__3143\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14635\
        );

    \I__3142\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14632\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14629\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__14651\,
            I => \N__14626\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__14650\,
            I => \N__14622\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__14649\,
            I => \N__14617\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__14646\,
            I => \N__14614\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__14641\,
            I => \N__14611\
        );

    \I__3135\ : Span4Mux_h
    port map (
            O => \N__14638\,
            I => \N__14602\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__14635\,
            I => \N__14602\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__14632\,
            I => \N__14602\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__14629\,
            I => \N__14602\
        );

    \I__3131\ : InMux
    port map (
            O => \N__14626\,
            I => \N__14589\
        );

    \I__3130\ : InMux
    port map (
            O => \N__14625\,
            I => \N__14589\
        );

    \I__3129\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14589\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14589\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14589\
        );

    \I__3126\ : InMux
    port map (
            O => \N__14617\,
            I => \N__14589\
        );

    \I__3125\ : Odrv12
    port map (
            O => \N__14614\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__14611\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__14602\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__14589\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__3121\ : CEMux
    port map (
            O => \N__14580\,
            I => \N__14575\
        );

    \I__3120\ : CEMux
    port map (
            O => \N__14579\,
            I => \N__14572\
        );

    \I__3119\ : CEMux
    port map (
            O => \N__14578\,
            I => \N__14569\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14566\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__14572\,
            I => \N__14563\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14569\,
            I => \N__14560\
        );

    \I__3115\ : Span4Mux_h
    port map (
            O => \N__14566\,
            I => \N__14557\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__14563\,
            I => \N__14554\
        );

    \I__3113\ : Span4Mux_v
    port map (
            O => \N__14560\,
            I => \N__14551\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__14557\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__14554\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__3110\ : Odrv4
    port map (
            O => \N__14551\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__14544\,
            I => \uu2.mem0.G_13_0_a2_1_cascade_\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14541\,
            I => \N__14538\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__14538\,
            I => \N__14535\
        );

    \I__3106\ : Odrv12
    port map (
            O => \N__14535\,
            I => \uu2.mem0.G_13_0_a3_1_2\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__14532\,
            I => \N__14522\
        );

    \I__3104\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14516\
        );

    \I__3103\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14513\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14510\
        );

    \I__3101\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14505\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14527\,
            I => \N__14505\
        );

    \I__3099\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14498\
        );

    \I__3098\ : InMux
    port map (
            O => \N__14525\,
            I => \N__14498\
        );

    \I__3097\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14493\
        );

    \I__3096\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14493\
        );

    \I__3095\ : InMux
    port map (
            O => \N__14520\,
            I => \N__14488\
        );

    \I__3094\ : InMux
    port map (
            O => \N__14519\,
            I => \N__14488\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__14516\,
            I => \N__14481\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__14513\,
            I => \N__14481\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__14510\,
            I => \N__14478\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14475\
        );

    \I__3089\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14470\
        );

    \I__3088\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14470\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__14498\,
            I => \N__14463\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__14493\,
            I => \N__14463\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__14488\,
            I => \N__14463\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14457\
        );

    \I__3083\ : InMux
    port map (
            O => \N__14486\,
            I => \N__14454\
        );

    \I__3082\ : Span4Mux_v
    port map (
            O => \N__14481\,
            I => \N__14451\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__14478\,
            I => \N__14442\
        );

    \I__3080\ : Span4Mux_v
    port map (
            O => \N__14475\,
            I => \N__14442\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14470\,
            I => \N__14442\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__14463\,
            I => \N__14442\
        );

    \I__3077\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14437\
        );

    \I__3076\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14437\
        );

    \I__3075\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14434\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__14457\,
            I => \L3_tx_data_rdy\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__14454\,
            I => \L3_tx_data_rdy\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__14451\,
            I => \L3_tx_data_rdy\
        );

    \I__3071\ : Odrv4
    port map (
            O => \N__14442\,
            I => \L3_tx_data_rdy\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__14437\,
            I => \L3_tx_data_rdy\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__14434\,
            I => \L3_tx_data_rdy\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14421\,
            I => \N__14418\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__14418\,
            I => \N__14415\
        );

    \I__3066\ : Span4Mux_h
    port map (
            O => \N__14415\,
            I => \N__14410\
        );

    \I__3065\ : InMux
    port map (
            O => \N__14414\,
            I => \N__14405\
        );

    \I__3064\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14405\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__14410\,
            I => \L3_tx_data_1\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__14405\,
            I => \L3_tx_data_1\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__14400\,
            I => \uu2.mem0.G_13_0_a2_2_cascade_\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14391\
        );

    \I__3059\ : InMux
    port map (
            O => \N__14396\,
            I => \N__14381\
        );

    \I__3058\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14376\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14376\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14391\,
            I => \N__14371\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14390\,
            I => \N__14362\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14362\
        );

    \I__3053\ : InMux
    port map (
            O => \N__14388\,
            I => \N__14362\
        );

    \I__3052\ : InMux
    port map (
            O => \N__14387\,
            I => \N__14362\
        );

    \I__3051\ : InMux
    port map (
            O => \N__14386\,
            I => \N__14357\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14385\,
            I => \N__14357\
        );

    \I__3049\ : InMux
    port map (
            O => \N__14384\,
            I => \N__14354\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__14381\,
            I => \N__14348\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14345\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14375\,
            I => \N__14340\
        );

    \I__3045\ : InMux
    port map (
            O => \N__14374\,
            I => \N__14340\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14337\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14362\,
            I => \N__14332\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14332\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__14354\,
            I => \N__14329\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14353\,
            I => \N__14325\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14352\,
            I => \N__14320\
        );

    \I__3038\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14320\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__14348\,
            I => \N__14313\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__14345\,
            I => \N__14313\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14313\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__14337\,
            I => \N__14308\
        );

    \I__3033\ : Span4Mux_h
    port map (
            O => \N__14332\,
            I => \N__14308\
        );

    \I__3032\ : Span4Mux_h
    port map (
            O => \N__14329\,
            I => \N__14305\
        );

    \I__3031\ : InMux
    port map (
            O => \N__14328\,
            I => \N__14302\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__14325\,
            I => \N_96\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__14320\,
            I => \N_96\
        );

    \I__3028\ : Odrv4
    port map (
            O => \N__14313\,
            I => \N_96\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__14308\,
            I => \N_96\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__14305\,
            I => \N_96\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__14302\,
            I => \N_96\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14289\,
            I => \N__14286\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__14286\,
            I => \N__14283\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__14283\,
            I => \N__14280\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__14280\,
            I => \uu2.mem0.G_13_0_0\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14274\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__14274\,
            I => \N__14271\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__14271\,
            I => \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0\
        );

    \I__3017\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14261\
        );

    \I__3016\ : InMux
    port map (
            O => \N__14267\,
            I => \N__14261\
        );

    \I__3015\ : InMux
    port map (
            O => \N__14266\,
            I => \N__14256\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__14261\,
            I => \N__14252\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14247\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14259\,
            I => \N__14247\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14256\,
            I => \N__14238\
        );

    \I__3010\ : InMux
    port map (
            O => \N__14255\,
            I => \N__14235\
        );

    \I__3009\ : Span4Mux_h
    port map (
            O => \N__14252\,
            I => \N__14232\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__14247\,
            I => \N__14229\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14246\,
            I => \N__14224\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14245\,
            I => \N__14224\
        );

    \I__3005\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14217\
        );

    \I__3004\ : InMux
    port map (
            O => \N__14243\,
            I => \N__14217\
        );

    \I__3003\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14217\
        );

    \I__3002\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14213\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__14238\,
            I => \N__14208\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__14235\,
            I => \N__14208\
        );

    \I__2999\ : Span4Mux_v
    port map (
            O => \N__14232\,
            I => \N__14205\
        );

    \I__2998\ : Span4Mux_v
    port map (
            O => \N__14229\,
            I => \N__14202\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14224\,
            I => \N__14197\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__14217\,
            I => \N__14197\
        );

    \I__2995\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14194\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14213\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__14208\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2992\ : Odrv4
    port map (
            O => \N__14205\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__14202\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2990\ : Odrv12
    port map (
            O => \N__14197\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__14194\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__2988\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14172\
        );

    \I__2987\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14172\
        );

    \I__2986\ : InMux
    port map (
            O => \N__14179\,
            I => \N__14167\
        );

    \I__2985\ : InMux
    port map (
            O => \N__14178\,
            I => \N__14167\
        );

    \I__2984\ : InMux
    port map (
            O => \N__14177\,
            I => \N__14163\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__14172\,
            I => \N__14155\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__14167\,
            I => \N__14155\
        );

    \I__2981\ : InMux
    port map (
            O => \N__14166\,
            I => \N__14151\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__14163\,
            I => \N__14148\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14162\,
            I => \N__14143\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14161\,
            I => \N__14143\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14160\,
            I => \N__14140\
        );

    \I__2976\ : Span4Mux_h
    port map (
            O => \N__14155\,
            I => \N__14137\
        );

    \I__2975\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14133\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__14151\,
            I => \N__14130\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__14148\,
            I => \N__14125\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14143\,
            I => \N__14125\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14120\
        );

    \I__2970\ : Span4Mux_v
    port map (
            O => \N__14137\,
            I => \N__14120\
        );

    \I__2969\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14117\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__14133\,
            I => \N__14114\
        );

    \I__2967\ : Odrv4
    port map (
            O => \N__14130\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__14125\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2965\ : Odrv4
    port map (
            O => \N__14120\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__14117\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2963\ : Odrv12
    port map (
            O => \N__14114\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__2962\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14095\
        );

    \I__2961\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14092\
        );

    \I__2960\ : CascadeMux
    port map (
            O => \N__14101\,
            I => \N__14089\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__14100\,
            I => \N__14086\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__14099\,
            I => \N__14080\
        );

    \I__2957\ : CascadeMux
    port map (
            O => \N__14098\,
            I => \N__14077\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__14095\,
            I => \N__14073\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__14092\,
            I => \N__14070\
        );

    \I__2954\ : InMux
    port map (
            O => \N__14089\,
            I => \N__14065\
        );

    \I__2953\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14065\
        );

    \I__2952\ : CascadeMux
    port map (
            O => \N__14085\,
            I => \N__14062\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__14084\,
            I => \N__14059\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__14083\,
            I => \N__14054\
        );

    \I__2949\ : InMux
    port map (
            O => \N__14080\,
            I => \N__14049\
        );

    \I__2948\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14049\
        );

    \I__2947\ : InMux
    port map (
            O => \N__14076\,
            I => \N__14046\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__14073\,
            I => \N__14043\
        );

    \I__2945\ : Span12Mux_v
    port map (
            O => \N__14070\,
            I => \N__14038\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__14065\,
            I => \N__14038\
        );

    \I__2943\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14033\
        );

    \I__2942\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14033\
        );

    \I__2941\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14026\
        );

    \I__2940\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14026\
        );

    \I__2939\ : InMux
    port map (
            O => \N__14054\,
            I => \N__14026\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__14049\,
            I => \N__14021\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__14046\,
            I => \N__14021\
        );

    \I__2936\ : Odrv4
    port map (
            O => \N__14043\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2935\ : Odrv12
    port map (
            O => \N__14038\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__14033\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__14026\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2932\ : Odrv12
    port map (
            O => \N__14021\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__14010\,
            I => \Lab_UT.bcd2segment1.N_248_cascade_\
        );

    \I__2930\ : InMux
    port map (
            O => \N__14007\,
            I => \N__14004\
        );

    \I__2929\ : LocalMux
    port map (
            O => \N__14004\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14001\,
            I => \N__13998\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__13998\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13992\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__13992\,
            I => \uu2.m76_bm_1_0\
        );

    \I__2924\ : InMux
    port map (
            O => \N__13989\,
            I => \N__13986\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__13986\,
            I => \N__13982\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__13985\,
            I => \N__13977\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__13982\,
            I => \N__13974\
        );

    \I__2920\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13971\
        );

    \I__2919\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13966\
        );

    \I__2918\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13966\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__13974\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__13971\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__13966\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__2914\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13956\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13953\
        );

    \I__2912\ : Span4Mux_h
    port map (
            O => \N__13953\,
            I => \N__13950\
        );

    \I__2911\ : Span4Mux_h
    port map (
            O => \N__13950\,
            I => \N__13947\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__13947\,
            I => \uu2.mem0.g1_2_2\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13944\,
            I => \N__13941\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__13941\,
            I => \N__13938\
        );

    \I__2907\ : Span12Mux_s8_h
    port map (
            O => \N__13938\,
            I => \N__13935\
        );

    \I__2906\ : Odrv12
    port map (
            O => \N__13935\,
            I => \uu2.mem0.g2_0_0_0_0\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13932\,
            I => \N__13929\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13929\,
            I => \N__13926\
        );

    \I__2903\ : Span4Mux_h
    port map (
            O => \N__13926\,
            I => \N__13923\
        );

    \I__2902\ : Odrv4
    port map (
            O => \N__13923\,
            I => \uu2.mem0.g2_2\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__13920\,
            I => \N__13914\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__13919\,
            I => \N__13909\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__13918\,
            I => \N__13905\
        );

    \I__2898\ : CascadeMux
    port map (
            O => \N__13917\,
            I => \N__13901\
        );

    \I__2897\ : InMux
    port map (
            O => \N__13914\,
            I => \N__13897\
        );

    \I__2896\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13894\
        );

    \I__2895\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13891\
        );

    \I__2894\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13888\
        );

    \I__2893\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13884\
        );

    \I__2892\ : InMux
    port map (
            O => \N__13905\,
            I => \N__13881\
        );

    \I__2891\ : InMux
    port map (
            O => \N__13904\,
            I => \N__13874\
        );

    \I__2890\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13874\
        );

    \I__2889\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13874\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__13897\,
            I => \N__13871\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__13894\,
            I => \N__13868\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13865\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__13888\,
            I => \N__13862\
        );

    \I__2884\ : InMux
    port map (
            O => \N__13887\,
            I => \N__13859\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__13884\,
            I => \N__13856\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__13881\,
            I => \N__13851\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__13874\,
            I => \N__13851\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__13871\,
            I => \N__13842\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__13868\,
            I => \N__13842\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__13865\,
            I => \N__13842\
        );

    \I__2877\ : Span4Mux_h
    port map (
            O => \N__13862\,
            I => \N__13842\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__13859\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__13856\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__2874\ : Odrv4
    port map (
            O => \N__13851\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__13842\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__2872\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__13830\,
            I => \N__13823\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13820\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__13828\,
            I => \N__13817\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__13827\,
            I => \N__13812\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13807\
        );

    \I__2866\ : Span4Mux_h
    port map (
            O => \N__13823\,
            I => \N__13804\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__13820\,
            I => \N__13801\
        );

    \I__2864\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13794\
        );

    \I__2863\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13794\
        );

    \I__2862\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13794\
        );

    \I__2861\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13787\
        );

    \I__2860\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13787\
        );

    \I__2859\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13787\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__13807\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2857\ : Odrv4
    port map (
            O => \N__13804\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__13801\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__13794\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__13787\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2853\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13773\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__13773\,
            I => \N__13767\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__13772\,
            I => \N__13763\
        );

    \I__2850\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13758\
        );

    \I__2849\ : InMux
    port map (
            O => \N__13770\,
            I => \N__13755\
        );

    \I__2848\ : Span4Mux_h
    port map (
            O => \N__13767\,
            I => \N__13752\
        );

    \I__2847\ : InMux
    port map (
            O => \N__13766\,
            I => \N__13749\
        );

    \I__2846\ : InMux
    port map (
            O => \N__13763\,
            I => \N__13742\
        );

    \I__2845\ : InMux
    port map (
            O => \N__13762\,
            I => \N__13742\
        );

    \I__2844\ : InMux
    port map (
            O => \N__13761\,
            I => \N__13742\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__13758\,
            I => \Lab_UT.state_2\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__13755\,
            I => \Lab_UT.state_2\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__13752\,
            I => \Lab_UT.state_2\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__13749\,
            I => \Lab_UT.state_2\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__13742\,
            I => \Lab_UT.state_2\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13731\,
            I => \N__13728\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__13728\,
            I => \Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\
        );

    \I__2835\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13719\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__13719\,
            I => \N__13716\
        );

    \I__2833\ : Span4Mux_s3_v
    port map (
            O => \N__13716\,
            I => \N__13713\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__13713\,
            I => \N__13710\
        );

    \I__2831\ : Odrv4
    port map (
            O => \N__13710\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_1\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13707\,
            I => \N__13704\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__13704\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2828\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13698\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__13698\,
            I => \uu2.m76_am_1\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__13695\,
            I => \N__13692\
        );

    \I__2825\ : InMux
    port map (
            O => \N__13692\,
            I => \N__13689\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__13689\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2823\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13683\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__13683\,
            I => \N__13680\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__13680\,
            I => \Lab_UT.bcd2segment1.N_244\
        );

    \I__2820\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13673\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13670\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__13673\,
            I => \N__13667\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__13670\,
            I => \N__13664\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__13667\,
            I => \N__13661\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__13664\,
            I => \N__13658\
        );

    \I__2814\ : Odrv4
    port map (
            O => \N__13661\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2813\ : Odrv4
    port map (
            O => \N__13658\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__13653\,
            I => \Lab_UT.bcd2segment1.N_246_cascade_\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__13650\,
            I => \Lab_UT.dictrl.un1_state_11_cascade_\
        );

    \I__2810\ : SRMux
    port map (
            O => \N__13647\,
            I => \N__13644\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__13644\,
            I => \N__13641\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__13641\,
            I => \N__13637\
        );

    \I__2807\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13634\
        );

    \I__2806\ : Odrv4
    port map (
            O => \N__13637\,
            I => \Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__13634\,
            I => \Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1\
        );

    \I__2804\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13623\
        );

    \I__2803\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13618\
        );

    \I__2802\ : InMux
    port map (
            O => \N__13627\,
            I => \N__13618\
        );

    \I__2801\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13615\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__13623\,
            I => \N__13612\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__13618\,
            I => \N__13609\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__13615\,
            I => \N__13602\
        );

    \I__2797\ : Span4Mux_h
    port map (
            O => \N__13612\,
            I => \N__13602\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__13609\,
            I => \N__13602\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__13602\,
            I => \N__13599\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__13599\,
            I => \Lab_UT.bcd2segment1.N_264\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__13596\,
            I => \Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_\
        );

    \I__2792\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13590\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13587\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__13587\,
            I => \N__13582\
        );

    \I__2789\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13579\
        );

    \I__2788\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13576\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__13582\,
            I => \Lab_UT.dictrl.next_state16Z0Z_5\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__13579\,
            I => \Lab_UT.dictrl.next_state16Z0Z_5\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__13576\,
            I => \Lab_UT.dictrl.next_state16Z0Z_5\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__13569\,
            I => \Lab_UT.m68_0_ns_cascade_\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13566\,
            I => \N__13561\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13565\,
            I => \N__13558\
        );

    \I__2781\ : InMux
    port map (
            O => \N__13564\,
            I => \N__13555\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__13561\,
            I => \Lab_UT.dictrl.next_state16Z0Z_4\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__13558\,
            I => \Lab_UT.dictrl.next_state16Z0Z_4\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__13555\,
            I => \Lab_UT.dictrl.next_state16Z0Z_4\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13545\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__13545\,
            I => \N__13539\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13532\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13532\
        );

    \I__2773\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13532\
        );

    \I__2772\ : Sp12to4
    port map (
            O => \N__13539\,
            I => \N__13526\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13526\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13531\,
            I => \N__13523\
        );

    \I__2769\ : Odrv12
    port map (
            O => \N__13526\,
            I => \Lab_UT.state_3\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__13523\,
            I => \Lab_UT.state_3\
        );

    \I__2767\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13511\
        );

    \I__2766\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13511\
        );

    \I__2765\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13508\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__13511\,
            I => \N__13499\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__13508\,
            I => \N__13499\
        );

    \I__2762\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13496\
        );

    \I__2761\ : InMux
    port map (
            O => \N__13506\,
            I => \N__13489\
        );

    \I__2760\ : InMux
    port map (
            O => \N__13505\,
            I => \N__13489\
        );

    \I__2759\ : InMux
    port map (
            O => \N__13504\,
            I => \N__13489\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__13499\,
            I => \Lab_UT.state_1\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__13496\,
            I => \Lab_UT.state_1\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__13489\,
            I => \Lab_UT.state_1\
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__13482\,
            I => \Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__13479\,
            I => \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__13476\,
            I => \N__13472\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__13475\,
            I => \N__13469\
        );

    \I__2751\ : InMux
    port map (
            O => \N__13472\,
            I => \N__13466\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13469\,
            I => \N__13463\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__13466\,
            I => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__13463\,
            I => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\
        );

    \I__2747\ : InMux
    port map (
            O => \N__13458\,
            I => \N__13453\
        );

    \I__2746\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13448\
        );

    \I__2745\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13448\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__13453\,
            I => \N__13445\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13442\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__13445\,
            I => \N__13439\
        );

    \I__2741\ : Span4Mux_h
    port map (
            O => \N__13442\,
            I => \N__13436\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__13439\,
            I => \Lab_UT.dictrl.next_state_set\
        );

    \I__2739\ : Odrv4
    port map (
            O => \N__13436\,
            I => \Lab_UT.dictrl.next_state_set\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__13431\,
            I => \buart.Z_rx.bitcount_lm_3_cascade_\
        );

    \I__2737\ : SRMux
    port map (
            O => \N__13428\,
            I => \N__13424\
        );

    \I__2736\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13421\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__13424\,
            I => \N__13418\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__13421\,
            I => \N__13415\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__13418\,
            I => \Lab_UT.m72_0\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__13415\,
            I => \Lab_UT.m72_0\
        );

    \I__2731\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13400\
        );

    \I__2730\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13400\
        );

    \I__2729\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13400\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13397\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__13400\,
            I => \N__13394\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__13397\,
            I => \Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__13394\,
            I => \Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__13389\,
            I => \N__13386\
        );

    \I__2723\ : InMux
    port map (
            O => \N__13386\,
            I => \N__13383\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__13383\,
            I => \Lab_UT.un1_state_13\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__13380\,
            I => \Lab_UT.un1_state_13_cascade_\
        );

    \I__2720\ : InMux
    port map (
            O => \N__13377\,
            I => \N__13373\
        );

    \I__2719\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13370\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__13373\,
            I => \N__13365\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13370\,
            I => \N__13365\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__13365\,
            I => \N__13362\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__13362\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13359\,
            I => \N__13355\
        );

    \I__2713\ : InMux
    port map (
            O => \N__13358\,
            I => \N__13352\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__13355\,
            I => \N__13349\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__13352\,
            I => \N__13346\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__13349\,
            I => \N__13343\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__13346\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__13343\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__2707\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13335\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13335\,
            I => \Lab_UT.dictrl.un1_state_11\
        );

    \I__2705\ : CascadeMux
    port map (
            O => \N__13332\,
            I => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_\
        );

    \I__2704\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13326\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13323\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__13323\,
            I => \N__13320\
        );

    \I__2701\ : Odrv4
    port map (
            O => \N__13320\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__13317\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__2698\ : InMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__13305\,
            I => \N__13301\
        );

    \I__2695\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13298\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__13301\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__13298\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__2692\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13289\
        );

    \I__2691\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13286\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13283\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__13286\,
            I => \N__13280\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__13283\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__2687\ : Odrv4
    port map (
            O => \N__13280\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__13275\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3_cascade_\
        );

    \I__2685\ : InMux
    port map (
            O => \N__13272\,
            I => \N__13269\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__13269\,
            I => \N__13266\
        );

    \I__2683\ : Span4Mux_h
    port map (
            O => \N__13266\,
            I => \N__13261\
        );

    \I__2682\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13256\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13256\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__13261\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__13256\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__2678\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13248\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13248\,
            I => \N__13245\
        );

    \I__2676\ : Span4Mux_h
    port map (
            O => \N__13245\,
            I => \N__13242\
        );

    \I__2675\ : Odrv4
    port map (
            O => \N__13242\,
            I => \Lab_UT.dictrl.dicRun_2_reti\
        );

    \I__2674\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13236\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__13236\,
            I => \Lab_UT.dictrl.next_state_out_0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__13233\,
            I => \N__13229\
        );

    \I__2671\ : InMux
    port map (
            O => \N__13232\,
            I => \N__13226\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__13229\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__13226\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__13221\,
            I => \N__13218\
        );

    \I__2667\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13213\
        );

    \I__2666\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13210\
        );

    \I__2665\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13207\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__13213\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__13210\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13207\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__13200\,
            I => \Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_\
        );

    \I__2659\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13187\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__13190\,
            I => \N__13184\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__13187\,
            I => \N__13179\
        );

    \I__2655\ : InMux
    port map (
            O => \N__13184\,
            I => \N__13174\
        );

    \I__2654\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13174\
        );

    \I__2653\ : InMux
    port map (
            O => \N__13182\,
            I => \N__13171\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__13179\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__13174\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__13171\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__13164\,
            I => \N__13159\
        );

    \I__2648\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13155\
        );

    \I__2647\ : InMux
    port map (
            O => \N__13162\,
            I => \N__13148\
        );

    \I__2646\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13148\
        );

    \I__2645\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13148\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__13155\,
            I => \N__13145\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__13148\,
            I => \N__13142\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__13145\,
            I => \N__13139\
        );

    \I__2641\ : Span4Mux_h
    port map (
            O => \N__13142\,
            I => \N__13136\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__13139\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2639\ : Odrv4
    port map (
            O => \N__13136\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__2638\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13127\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13119\
        );

    \I__2636\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13119\
        );

    \I__2635\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13119\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__2633\ : Odrv12
    port map (
            O => \N__13116\,
            I => \Lab_UT.N_9_0\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__13113\,
            I => \N__13110\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13107\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13107\,
            I => \N__13103\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__13106\,
            I => \N__13099\
        );

    \I__2628\ : Sp12to4
    port map (
            O => \N__13103\,
            I => \N__13095\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13088\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13099\,
            I => \N__13088\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13098\,
            I => \N__13088\
        );

    \I__2624\ : Odrv12
    port map (
            O => \N__13095\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__13088\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13080\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__13080\,
            I => \N__13077\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__13077\,
            I => \Lab_UT.bcd2segment1.N_181\
        );

    \I__2619\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13071\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13068\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__13068\,
            I => \Lab_UT.bcd2segment1.N_229\
        );

    \I__2616\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13053\
        );

    \I__2615\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13053\
        );

    \I__2614\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13053\
        );

    \I__2613\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13053\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__13053\,
            I => \N__13045\
        );

    \I__2611\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13037\
        );

    \I__2610\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13037\
        );

    \I__2609\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13034\
        );

    \I__2608\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13031\
        );

    \I__2607\ : InMux
    port map (
            O => \N__13048\,
            I => \N__13028\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__13045\,
            I => \N__13025\
        );

    \I__2605\ : InMux
    port map (
            O => \N__13044\,
            I => \N__13018\
        );

    \I__2604\ : InMux
    port map (
            O => \N__13043\,
            I => \N__13018\
        );

    \I__2603\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13018\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__13037\,
            I => \N__13015\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__13034\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__13031\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__13028\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2598\ : Odrv4
    port map (
            O => \N__13025\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__13018\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__13015\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__2595\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12990\
        );

    \I__2594\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12990\
        );

    \I__2593\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12990\
        );

    \I__2592\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12990\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__12990\,
            I => \N__12982\
        );

    \I__2590\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12973\
        );

    \I__2589\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12973\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12973\
        );

    \I__2587\ : InMux
    port map (
            O => \N__12986\,
            I => \N__12973\
        );

    \I__2586\ : InMux
    port map (
            O => \N__12985\,
            I => \N__12968\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__12982\,
            I => \N__12963\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__12973\,
            I => \N__12960\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12954\
        );

    \I__2582\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12954\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__12968\,
            I => \N__12951\
        );

    \I__2580\ : InMux
    port map (
            O => \N__12967\,
            I => \N__12946\
        );

    \I__2579\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12946\
        );

    \I__2578\ : Sp12to4
    port map (
            O => \N__12963\,
            I => \N__12943\
        );

    \I__2577\ : Span4Mux_h
    port map (
            O => \N__12960\,
            I => \N__12940\
        );

    \I__2576\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12937\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__12954\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2574\ : Odrv4
    port map (
            O => \N__12951\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__12946\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__12943\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__12940\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__12937\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__12924\,
            I => \N__12917\
        );

    \I__2568\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12914\
        );

    \I__2567\ : InMux
    port map (
            O => \N__12922\,
            I => \N__12903\
        );

    \I__2566\ : InMux
    port map (
            O => \N__12921\,
            I => \N__12903\
        );

    \I__2565\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12903\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12903\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__12914\,
            I => \N__12898\
        );

    \I__2562\ : InMux
    port map (
            O => \N__12913\,
            I => \N__12893\
        );

    \I__2561\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12893\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__12903\,
            I => \N__12890\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__12902\,
            I => \N__12884\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__12901\,
            I => \N__12880\
        );

    \I__2557\ : Span4Mux_h
    port map (
            O => \N__12898\,
            I => \N__12877\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__12893\,
            I => \N__12872\
        );

    \I__2555\ : Span12Mux_s9_v
    port map (
            O => \N__12890\,
            I => \N__12872\
        );

    \I__2554\ : InMux
    port map (
            O => \N__12889\,
            I => \N__12863\
        );

    \I__2553\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12863\
        );

    \I__2552\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12863\
        );

    \I__2551\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12863\
        );

    \I__2550\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12858\
        );

    \I__2549\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12858\
        );

    \I__2548\ : Odrv4
    port map (
            O => \N__12877\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__12872\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__12863\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__12858\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__2544\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12846\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12846\,
            I => \N__12843\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__12843\,
            I => \Lab_UT.bcd2segment1.N_233\
        );

    \I__2541\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12836\
        );

    \I__2540\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12833\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__12836\,
            I => \N__12829\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__12833\,
            I => \N__12826\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12823\
        );

    \I__2536\ : Span4Mux_h
    port map (
            O => \N__12829\,
            I => \N__12820\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__12826\,
            I => \N__12817\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__12823\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__12820\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2532\ : Odrv4
    port map (
            O => \N__12817\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__2530\ : InMux
    port map (
            O => \N__12809\,
            I => \N__12797\
        );

    \I__2529\ : InMux
    port map (
            O => \N__12808\,
            I => \N__12797\
        );

    \I__2528\ : InMux
    port map (
            O => \N__12807\,
            I => \N__12797\
        );

    \I__2527\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12794\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12791\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__12794\,
            I => \N__12788\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__12791\,
            I => \N__12785\
        );

    \I__2523\ : Span4Mux_h
    port map (
            O => \N__12788\,
            I => \N__12782\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__12785\,
            I => \uu2.N_115\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__12782\,
            I => \uu2.N_115\
        );

    \I__2520\ : CascadeMux
    port map (
            O => \N__12777\,
            I => \N__12773\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12763\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12763\
        );

    \I__2517\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12763\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__12771\,
            I => \N__12760\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__12770\,
            I => \N__12756\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__12763\,
            I => \N__12750\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12760\,
            I => \N__12747\
        );

    \I__2512\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12744\
        );

    \I__2511\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12741\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__12755\,
            I => \N__12738\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__12754\,
            I => \N__12733\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__12753\,
            I => \N__12728\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__12750\,
            I => \N__12722\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__12747\,
            I => \N__12722\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__12744\,
            I => \N__12717\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__12741\,
            I => \N__12717\
        );

    \I__2503\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12710\
        );

    \I__2502\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12710\
        );

    \I__2501\ : InMux
    port map (
            O => \N__12736\,
            I => \N__12710\
        );

    \I__2500\ : InMux
    port map (
            O => \N__12733\,
            I => \N__12707\
        );

    \I__2499\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12700\
        );

    \I__2498\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12700\
        );

    \I__2497\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12700\
        );

    \I__2496\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12697\
        );

    \I__2495\ : Span4Mux_h
    port map (
            O => \N__12722\,
            I => \N__12694\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__12717\,
            I => \N__12691\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__12710\,
            I => \N__12686\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__12707\,
            I => \N__12686\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__12700\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__12697\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__12694\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__12691\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__12686\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__12675\,
            I => \Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_\
        );

    \I__2485\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12669\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__12669\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_0\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__12666\,
            I => \Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__12663\,
            I => \N__12660\
        );

    \I__2481\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12657\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__12657\,
            I => \N__12654\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__12654\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2478\ : InMux
    port map (
            O => \N__12651\,
            I => \N__12647\
        );

    \I__2477\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12644\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__12647\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__12644\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__12639\,
            I => \uu2.mem0.m317_0_a6_0_cascade_\
        );

    \I__2473\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12633\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__12630\,
            I => \uu2.mem0.N_6_0\
        );

    \I__2470\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__12624\,
            I => \uu2.mem0.m317_0_0\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__12621\,
            I => \uu2.mem0.N_11_0_0_cascade_\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12615\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__12615\,
            I => \N__12612\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__12612\,
            I => \uu2.mem0.N_6_0_0_0\
        );

    \I__2464\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12602\
        );

    \I__2463\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12602\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__12607\,
            I => \N__12596\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__12602\,
            I => \N__12591\
        );

    \I__2460\ : InMux
    port map (
            O => \N__12601\,
            I => \N__12582\
        );

    \I__2459\ : InMux
    port map (
            O => \N__12600\,
            I => \N__12582\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12582\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12582\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12577\
        );

    \I__2455\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12577\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__12591\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__12582\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__12577\,
            I => \uu2.w_addr_displaying_4_repZ0Z1\
        );

    \I__2451\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12567\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__12567\,
            I => \uu2.mem0.N_5_0\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12561\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__12561\,
            I => \uu2.mem0.N_14\
        );

    \I__2447\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12555\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N__12552\
        );

    \I__2445\ : Odrv12
    port map (
            O => \N__12552\,
            I => \uu2.mem0.g1_2_2_2_1\
        );

    \I__2444\ : InMux
    port map (
            O => \N__12549\,
            I => \N__12545\
        );

    \I__2443\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12542\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__12545\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__12542\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__12531\,
            I => \N__12528\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__12528\,
            I => \Lab_UT.bcd2segment1.N_239\
        );

    \I__2436\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12521\
        );

    \I__2435\ : InMux
    port map (
            O => \N__12524\,
            I => \N__12518\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__12521\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__12518\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__12513\,
            I => \N__12508\
        );

    \I__2431\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12505\
        );

    \I__2430\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12500\
        );

    \I__2429\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12500\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__12505\,
            I => \N__12495\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__12500\,
            I => \N__12495\
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__12495\,
            I => \uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8\
        );

    \I__2425\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12488\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12485\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__12488\,
            I => \N__12482\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__12485\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2421\ : Odrv4
    port map (
            O => \N__12482\,
            I => \uu2.w_addr_displaying_fastZ0Z_4\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__12477\,
            I => \N__12468\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12476\,
            I => \N__12465\
        );

    \I__2418\ : InMux
    port map (
            O => \N__12475\,
            I => \N__12462\
        );

    \I__2417\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12459\
        );

    \I__2416\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12456\
        );

    \I__2415\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12453\
        );

    \I__2414\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12448\
        );

    \I__2413\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12448\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__12465\,
            I => \N__12444\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__12462\,
            I => \N__12441\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__12459\,
            I => \N__12434\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__12456\,
            I => \N__12434\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__12453\,
            I => \N__12434\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__12448\,
            I => \N__12429\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12447\,
            I => \N__12421\
        );

    \I__2405\ : Span4Mux_h
    port map (
            O => \N__12444\,
            I => \N__12418\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__12441\,
            I => \N__12415\
        );

    \I__2403\ : Span4Mux_v
    port map (
            O => \N__12434\,
            I => \N__12412\
        );

    \I__2402\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12409\
        );

    \I__2401\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12406\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__12429\,
            I => \N__12403\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12398\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12398\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12426\,
            I => \N__12391\
        );

    \I__2396\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12391\
        );

    \I__2395\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12391\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12421\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__12418\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2392\ : Odrv4
    port map (
            O => \N__12415\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__12412\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__12409\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__12406\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2388\ : Odrv4
    port map (
            O => \N__12403\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__12398\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12391\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2385\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12369\,
            I => \N__12364\
        );

    \I__2383\ : InMux
    port map (
            O => \N__12368\,
            I => \N__12361\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__12367\,
            I => \N__12355\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__12364\,
            I => \N__12348\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__12361\,
            I => \N__12348\
        );

    \I__2379\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12345\
        );

    \I__2378\ : InMux
    port map (
            O => \N__12359\,
            I => \N__12342\
        );

    \I__2377\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12332\
        );

    \I__2376\ : InMux
    port map (
            O => \N__12355\,
            I => \N__12332\
        );

    \I__2375\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12332\
        );

    \I__2374\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12332\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__12348\,
            I => \N__12321\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__12345\,
            I => \N__12316\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12316\
        );

    \I__2370\ : InMux
    port map (
            O => \N__12341\,
            I => \N__12313\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__12332\,
            I => \N__12310\
        );

    \I__2368\ : InMux
    port map (
            O => \N__12331\,
            I => \N__12303\
        );

    \I__2367\ : InMux
    port map (
            O => \N__12330\,
            I => \N__12303\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12303\
        );

    \I__2365\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12300\
        );

    \I__2364\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12293\
        );

    \I__2363\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12293\
        );

    \I__2362\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12293\
        );

    \I__2361\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12290\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__12321\,
            I => \N__12287\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__12316\,
            I => \N__12282\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12282\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__12310\,
            I => \N__12279\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12276\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__12300\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__12293\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__12290\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__12287\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__12282\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__12279\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__12276\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12261\,
            I => \N__12258\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__12258\,
            I => \N__12254\
        );

    \I__2346\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12251\
        );

    \I__2345\ : Odrv12
    port map (
            O => \N__12254\,
            I => \uu2.N_9_i\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__12251\,
            I => \uu2.N_9_i\
        );

    \I__2343\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12242\
        );

    \I__2342\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12239\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__12242\,
            I => \N__12234\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__12239\,
            I => \N__12234\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__12234\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__12231\,
            I => \uu2.mem0.N_9_cascade_\
        );

    \I__2337\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12225\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__12225\,
            I => \uu2.mem0.N_15\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12217\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12210\
        );

    \I__2333\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12204\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__12217\,
            I => \N__12201\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12196\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12196\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12214\,
            I => \N__12193\
        );

    \I__2328\ : InMux
    port map (
            O => \N__12213\,
            I => \N__12188\
        );

    \I__2327\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12188\
        );

    \I__2326\ : InMux
    port map (
            O => \N__12209\,
            I => \N__12181\
        );

    \I__2325\ : InMux
    port map (
            O => \N__12208\,
            I => \N__12181\
        );

    \I__2324\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12181\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__12204\,
            I => \N__12178\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__12201\,
            I => \N__12173\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__12196\,
            I => \N__12173\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12193\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__12188\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__12181\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2317\ : Odrv12
    port map (
            O => \N__12178\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__12173\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__2315\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12159\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__12159\,
            I => \N__12156\
        );

    \I__2313\ : Odrv4
    port map (
            O => \N__12156\,
            I => \uu2.mem0.N_7\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \uu2.N_126_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12150\,
            I => \N__12143\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12139\
        );

    \I__2309\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12136\
        );

    \I__2308\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12131\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12146\,
            I => \N__12131\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12143\,
            I => \N__12128\
        );

    \I__2305\ : InMux
    port map (
            O => \N__12142\,
            I => \N__12125\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__12139\,
            I => \N__12120\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__12136\,
            I => \N__12120\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__12131\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2301\ : Odrv12
    port map (
            O => \N__12128\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__12125\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2299\ : Odrv4
    port map (
            O => \N__12120\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__2298\ : CascadeMux
    port map (
            O => \N__12111\,
            I => \N__12108\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12108\,
            I => \N__12105\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__12105\,
            I => \N__12102\
        );

    \I__2295\ : Odrv12
    port map (
            O => \N__12102\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0\
        );

    \I__2294\ : InMux
    port map (
            O => \N__12099\,
            I => \N__12096\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__12096\,
            I => \N__12093\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__12090\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_67\
        );

    \I__2290\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12084\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__12084\,
            I => \N__12081\
        );

    \I__2288\ : Span4Mux_h
    port map (
            O => \N__12081\,
            I => \N__12078\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__12078\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_66\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12071\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12068\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__12071\,
            I => \N__12065\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__12068\,
            I => \N__12060\
        );

    \I__2282\ : Span4Mux_h
    port map (
            O => \N__12065\,
            I => \N__12057\
        );

    \I__2281\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12052\
        );

    \I__2280\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12052\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__12060\,
            I => \uu2.N_126\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__12057\,
            I => \uu2.N_126\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__12052\,
            I => \uu2.N_126\
        );

    \I__2276\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12042\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__12042\,
            I => \N__12039\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__12039\,
            I => \N__12036\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__12036\,
            I => \N__12033\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__12033\,
            I => \uu2.mem0.g0_7_0_0\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__12030\,
            I => \uu2.mem0.N_57_cascade_\
        );

    \I__2270\ : InMux
    port map (
            O => \N__12027\,
            I => \N__12024\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__12024\,
            I => \uu2.mem0.bitmap_pmux_u_i_5_1\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12021\,
            I => \N__12018\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__12018\,
            I => \uu2.mem0.g0_7_0_3\
        );

    \I__2266\ : InMux
    port map (
            O => \N__12015\,
            I => \N__12012\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__12012\,
            I => \uu2.N_16\
        );

    \I__2264\ : CascadeMux
    port map (
            O => \N__12009\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_\
        );

    \I__2263\ : InMux
    port map (
            O => \N__12006\,
            I => \N__12003\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__12003\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_57\
        );

    \I__2261\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11997\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__11997\,
            I => \uu2.mem0.N_13_0\
        );

    \I__2259\ : InMux
    port map (
            O => \N__11994\,
            I => \N__11990\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11987\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__11990\,
            I => \uu2.N_8\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__11987\,
            I => \uu2.N_8\
        );

    \I__2255\ : CascadeMux
    port map (
            O => \N__11982\,
            I => \Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__11979\,
            I => \uu2.N_1580_0_cascade_\
        );

    \I__2253\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11973\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11969\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__11972\,
            I => \N__11966\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__11969\,
            I => \N__11963\
        );

    \I__2249\ : InMux
    port map (
            O => \N__11966\,
            I => \N__11960\
        );

    \I__2248\ : Odrv4
    port map (
            O => \N__11963\,
            I => \uu2.N_77_0\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__11960\,
            I => \uu2.N_77_0\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11947\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11947\
        );

    \I__2244\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11944\
        );

    \I__2243\ : InMux
    port map (
            O => \N__11952\,
            I => \N__11940\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__11947\,
            I => \N__11933\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__11944\,
            I => \N__11930\
        );

    \I__2240\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11927\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__11940\,
            I => \N__11924\
        );

    \I__2238\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11919\
        );

    \I__2237\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11919\
        );

    \I__2236\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11914\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11914\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__11933\,
            I => \N__11911\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__11930\,
            I => \N__11908\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__11927\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__11924\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11919\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__11914\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__11911\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__11908\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__2226\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__11892\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__11889\,
            I => \N__11886\
        );

    \I__2223\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__11883\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11877\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11877\,
            I => \uu2.N_1581_0\
        );

    \I__2219\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11871\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__11871\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2217\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11865\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__2215\ : Span4Mux_h
    port map (
            O => \N__11862\,
            I => \N__11857\
        );

    \I__2214\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11852\
        );

    \I__2213\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11852\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__11857\,
            I => \L3_tx_data_5\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__11852\,
            I => \L3_tx_data_5\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__11847\,
            I => \uu2.mem0.N_134_mux_cascade_\
        );

    \I__2209\ : InMux
    port map (
            O => \N__11844\,
            I => \N__11840\
        );

    \I__2208\ : InMux
    port map (
            O => \N__11843\,
            I => \N__11837\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11840\,
            I => \N__11831\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__11837\,
            I => \N__11828\
        );

    \I__2205\ : InMux
    port map (
            O => \N__11836\,
            I => \N__11821\
        );

    \I__2204\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11821\
        );

    \I__2203\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11821\
        );

    \I__2202\ : Span4Mux_h
    port map (
            O => \N__11831\,
            I => \N__11818\
        );

    \I__2201\ : Span4Mux_h
    port map (
            O => \N__11828\,
            I => \N__11813\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11813\
        );

    \I__2199\ : Odrv4
    port map (
            O => \N__11818\,
            I => \uu2.w_data_i_0_tzZ0Z_0\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__11813\,
            I => \uu2.w_data_i_0_tzZ0Z_0\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__2195\ : Span12Mux_s7_h
    port map (
            O => \N__11802\,
            I => \N__11799\
        );

    \I__2194\ : Odrv12
    port map (
            O => \N__11799\,
            I => \uu2.mem0.N_60_0_i\
        );

    \I__2193\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11793\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__11793\,
            I => \uu2.mem0.N_55_0\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__11790\,
            I => \Lab_UT.bcd2segment1.N_127_mux_cascade_\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__11787\,
            I => \Lab_UT.bcd2segment1.N_235_cascade_\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \Lab_UT.bcd2segment1.N_237_cascade_\
        );

    \I__2188\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__11778\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__2186\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__11772\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__2184\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__2183\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11763\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__11763\,
            I => \uu2.N_101_0\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \Lab_UT.bcd2segment1.N_242_cascade_\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__2178\ : Odrv12
    port map (
            O => \N__11751\,
            I => \resetGen.escKeyZ0Z_5\
        );

    \I__2177\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__11745\,
            I => \Lab_UT.dictrl.next_state_set_0_1\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__11742\,
            I => \N__11737\
        );

    \I__2174\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11734\
        );

    \I__2173\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11728\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11725\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__11734\,
            I => \N__11722\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11733\,
            I => \N__11715\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11732\,
            I => \N__11715\
        );

    \I__2168\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11715\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__11728\,
            I => bu_rx_data_6
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__11725\,
            I => bu_rx_data_6
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__11722\,
            I => bu_rx_data_6
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__11715\,
            I => bu_rx_data_6
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__11706\,
            I => \N__11699\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__11705\,
            I => \N__11696\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__11704\,
            I => \N__11693\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__11703\,
            I => \N__11689\
        );

    \I__2159\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11684\
        );

    \I__2158\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11684\
        );

    \I__2157\ : InMux
    port map (
            O => \N__11696\,
            I => \N__11681\
        );

    \I__2156\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11674\
        );

    \I__2155\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11674\
        );

    \I__2154\ : InMux
    port map (
            O => \N__11689\,
            I => \N__11674\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__11684\,
            I => bu_rx_data_7
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__11681\,
            I => bu_rx_data_7
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__11674\,
            I => bu_rx_data_7
        );

    \I__2150\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11662\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__11666\,
            I => \N__11657\
        );

    \I__2148\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11653\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__11662\,
            I => \N__11650\
        );

    \I__2146\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11647\
        );

    \I__2145\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11640\
        );

    \I__2144\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11640\
        );

    \I__2143\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11640\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__11653\,
            I => bu_rx_data_4
        );

    \I__2141\ : Odrv4
    port map (
            O => \N__11650\,
            I => bu_rx_data_4
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__11647\,
            I => bu_rx_data_4
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__11640\,
            I => bu_rx_data_4
        );

    \I__2138\ : InMux
    port map (
            O => \N__11631\,
            I => \N__11628\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__11628\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__11625\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_\
        );

    \I__2135\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11616\
        );

    \I__2134\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11616\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__11616\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__11613\,
            I => \Lab_UT.dictrl.un1_state_16_cascade_\
        );

    \I__2131\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11607\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11604\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__11604\,
            I => \N__11596\
        );

    \I__2128\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11591\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11591\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11588\
        );

    \I__2125\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11583\
        );

    \I__2124\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11583\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__11596\,
            I => bu_rx_data_5
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__11591\,
            I => bu_rx_data_5
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__11588\,
            I => bu_rx_data_5
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__11583\,
            I => bu_rx_data_5
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11571\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11571\,
            I => \N__11566\
        );

    \I__2117\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11563\
        );

    \I__2116\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11556\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__11566\,
            I => \N__11551\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__11563\,
            I => \N__11551\
        );

    \I__2113\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11546\
        );

    \I__2112\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11546\
        );

    \I__2111\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11541\
        );

    \I__2110\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11541\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__11556\,
            I => bu_rx_data_1
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__11551\,
            I => bu_rx_data_1
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__11546\,
            I => bu_rx_data_1
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__11541\,
            I => bu_rx_data_1
        );

    \I__2105\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11525\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11521\
        );

    \I__2103\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11514\
        );

    \I__2102\ : InMux
    port map (
            O => \N__11529\,
            I => \N__11514\
        );

    \I__2101\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11514\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__11525\,
            I => \N__11511\
        );

    \I__2099\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11508\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11503\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__11514\,
            I => \N__11503\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__11511\,
            I => bu_rx_data_0
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__11508\,
            I => bu_rx_data_0
        );

    \I__2094\ : Odrv4
    port map (
            O => \N__11503\,
            I => bu_rx_data_0
        );

    \I__2093\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11492\
        );

    \I__2092\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11489\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__11492\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__11489\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2089\ : InMux
    port map (
            O => \N__11484\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__2088\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11478\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__11478\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__11475\,
            I => \N__11472\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11469\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__11469\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\
        );

    \I__2083\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11462\
        );

    \I__2082\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11459\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__11462\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11459\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2079\ : InMux
    port map (
            O => \N__11454\,
            I => \N__11451\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__11451\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__11448\,
            I => \N__11444\
        );

    \I__2076\ : InMux
    port map (
            O => \N__11447\,
            I => \N__11441\
        );

    \I__2075\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11438\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__11441\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__11438\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2072\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11430\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__11430\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_1\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__11424\,
            I => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_\
        );

    \I__2068\ : InMux
    port map (
            O => \N__11421\,
            I => \N__11418\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__11418\,
            I => \Lab_UT.dictrl.next_state_out_1\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \Lab_UT.dictrl.N_97_cascade_\
        );

    \I__2065\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_\
        );

    \I__2064\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11404\
        );

    \I__2063\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11401\
        );

    \I__2062\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11398\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__11404\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__11401\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__11398\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__11391\,
            I => \N__11385\
        );

    \I__2057\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11382\
        );

    \I__2056\ : InMux
    port map (
            O => \N__11389\,
            I => \N__11379\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11376\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11385\,
            I => \N__11373\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__11382\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__11379\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__11376\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__11373\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2049\ : InMux
    port map (
            O => \N__11364\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11358\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__11358\,
            I => \N__11354\
        );

    \I__2046\ : InMux
    port map (
            O => \N__11357\,
            I => \N__11351\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__11354\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11351\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2043\ : InMux
    port map (
            O => \N__11346\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__2042\ : InMux
    port map (
            O => \N__11343\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \Lab_UT.didp.did_alarmMatch_1_cascade_\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11334\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__11334\,
            I => \Lab_UT.zero\
        );

    \I__2038\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11325\
        );

    \I__2037\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11325\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__11325\,
            I => \Lab_UT.alarmMatch\
        );

    \I__2035\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11319\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11319\,
            I => \Lab_UT.didp.countrce3.did_alarmMatch_0\
        );

    \I__2033\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11313\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__11313\,
            I => \Lab_UT.q_5_3\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__11310\,
            I => \Lab_UT.q_5_0_cascade_\
        );

    \I__2030\ : InMux
    port map (
            O => \N__11307\,
            I => \N__11304\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11304\,
            I => \Lab_UT.q_5_2\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__11301\,
            I => \N__11298\
        );

    \I__2027\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11292\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11292\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__11292\,
            I => \N__11289\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__11289\,
            I => \N__11286\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__11286\,
            I => \Lab_UT.N_27_i\
        );

    \I__2022\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11280\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11280\,
            I => \N__11277\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__11277\,
            I => \N__11274\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__11274\,
            I => \resetGen.escKeyZ0Z_4\
        );

    \I__2018\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__11268\,
            I => \N__11261\
        );

    \I__2016\ : InMux
    port map (
            O => \N__11267\,
            I => \N__11252\
        );

    \I__2015\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11252\
        );

    \I__2014\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11252\
        );

    \I__2013\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11252\
        );

    \I__2012\ : Span4Mux_v
    port map (
            O => \N__11261\,
            I => \N__11247\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__11252\,
            I => \N__11247\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__11247\,
            I => \resetGen.escKeyZ0\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__11244\,
            I => \Lab_UT.bcd2segment1.i2_mux_cascade_\
        );

    \I__2008\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11238\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11234\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11231\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__11234\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__11231\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__11226\,
            I => \N__11223\
        );

    \I__2002\ : InMux
    port map (
            O => \N__11223\,
            I => \N__11217\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11217\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__11217\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__11214\,
            I => \uu2.m95_i_m2_i_m2_1_cascade_\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \uu2.N_16_cascade_\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__11208\,
            I => \N__11205\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11200\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__11204\,
            I => \N__11197\
        );

    \I__1994\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11194\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__11200\,
            I => \N__11191\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11188\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__11194\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__11191\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__11188\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__11181\,
            I => \N__11173\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__11180\,
            I => \N__11169\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \N__11165\
        );

    \I__1985\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11156\
        );

    \I__1984\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11156\
        );

    \I__1983\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11156\
        );

    \I__1982\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11153\
        );

    \I__1981\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11142\
        );

    \I__1980\ : InMux
    port map (
            O => \N__11169\,
            I => \N__11142\
        );

    \I__1979\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11142\
        );

    \I__1978\ : InMux
    port map (
            O => \N__11165\,
            I => \N__11142\
        );

    \I__1977\ : InMux
    port map (
            O => \N__11164\,
            I => \N__11139\
        );

    \I__1976\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11135\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__11156\,
            I => \N__11132\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11127\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11122\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11122\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11117\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__11139\,
            I => \N__11117\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11114\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__11135\,
            I => \N__11111\
        );

    \I__1967\ : Span4Mux_v
    port map (
            O => \N__11132\,
            I => \N__11108\
        );

    \I__1966\ : InMux
    port map (
            O => \N__11131\,
            I => \N__11103\
        );

    \I__1965\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11103\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__11127\,
            I => \N__11096\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__11122\,
            I => \N__11096\
        );

    \I__1962\ : Span4Mux_h
    port map (
            O => \N__11117\,
            I => \N__11096\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11114\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__11111\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__11108\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__11103\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__11096\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__1956\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__11082\,
            I => \N__11079\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__11079\,
            I => \uu2.N_67_1_0\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__11076\,
            I => \uu2.N_67_1_0_cascade_\
        );

    \I__1952\ : InMux
    port map (
            O => \N__11073\,
            I => \N__11070\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11067\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__11067\,
            I => \uu2.mem0.N_55_0_0_0\
        );

    \I__1949\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__11061\,
            I => \uu2.mem0.g2_1\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \Lab_UT.bcd2segment1.N_250_cascade_\
        );

    \I__1946\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__11052\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_34\
        );

    \I__1944\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__11046\,
            I => \N__11043\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__11043\,
            I => \N__11038\
        );

    \I__1941\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11033\
        );

    \I__1940\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11033\
        );

    \I__1939\ : Odrv4
    port map (
            O => \N__11038\,
            I => \L3_tx_data_2\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__11033\,
            I => \L3_tx_data_2\
        );

    \I__1937\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11025\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__11025\,
            I => \N__11022\
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__11022\,
            I => \uu2.mem0.N_93_i\
        );

    \I__1934\ : InMux
    port map (
            O => \N__11019\,
            I => \N__11016\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11016\,
            I => \uu2.mem0.N_57_0_0\
        );

    \I__1932\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11010\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__11010\,
            I => \uu2.mem0.N_67_0\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__11007\,
            I => \uu2.mem0.g0_1_cascade_\
        );

    \I__1929\ : InMux
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__11001\,
            I => \uu2.mem0.g0_2\
        );

    \I__1927\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10995\,
            I => \uu2.mem0.i14_mux\
        );

    \I__1925\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10989\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10986\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__10983\,
            I => \uu2.mem0.N_126_0\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__10980\,
            I => \uu2.mem0.g0_1_3_cascade_\
        );

    \I__1920\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__10974\,
            I => \uu2.mem0.G_13_0_a2_0_1\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__10971\,
            I => \uu2.mem0.N_22_cascade_\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__10965\,
            I => \N__10962\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__10962\,
            I => \N__10959\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__10959\,
            I => \uu2.mem0.N_66_0_i\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__10953\,
            I => \uu2.mem0.g0_i_m2_1\
        );

    \I__1911\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10944\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__10944\,
            I => \N__10941\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__10941\,
            I => \uu2.mem0.g2_0_0_0\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__1906\ : InMux
    port map (
            O => \N__10935\,
            I => \N__10932\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__10932\,
            I => \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__10929\,
            I => \uu2.mem0.N_92_0_cascade_\
        );

    \I__1903\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__10923\,
            I => \uu2.mem0.m73_ns_1_0\
        );

    \I__1901\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10917\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__10917\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_1_4\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__10914\,
            I => \N__10911\
        );

    \I__1898\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10905\
        );

    \I__1897\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10905\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__10905\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__1895\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10896\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10896\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__10896\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__10893\,
            I => \uu2.mem0.N_92_0_0_cascade_\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__10890\,
            I => \N__10887\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10884\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10881\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__10881\,
            I => \uu2.mem0.m73_ns_1_0_0_1\
        );

    \I__1887\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10875\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__10875\,
            I => \uu2.mem0.N_74_0\
        );

    \I__1885\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10869\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__10869\,
            I => \N__10866\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__10866\,
            I => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__10863\,
            I => \Lab_UT.bcd2segment1.N_194_cascade_\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__10860\,
            I => \buart.Z_rx.ser_clk_2_cascade_\
        );

    \I__1880\ : CascadeMux
    port map (
            O => \N__10857\,
            I => \Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__10854\,
            I => \N__10851\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10848\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__10848\,
            I => \N__10843\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10840\
        );

    \I__1875\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10837\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__10843\,
            I => \N__10834\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10840\,
            I => \N__10829\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__10837\,
            I => \N__10829\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__10834\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z4\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__10829\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z4\
        );

    \I__1869\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10821\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__10821\,
            I => \Lab_UT.dictrl.next_alarmstate4Z0Z_0\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__10818\,
            I => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__10815\,
            I => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__10812\,
            I => \Lab_UT.bcd2segment1.N_222_cascade_\
        );

    \I__1864\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10804\
        );

    \I__1863\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10798\
        );

    \I__1862\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10795\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__10804\,
            I => \N__10792\
        );

    \I__1860\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10785\
        );

    \I__1859\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10785\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10801\,
            I => \N__10785\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__10798\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__10795\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__10792\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__10785\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_1\
        );

    \I__1853\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10773\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__1851\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10764\
        );

    \I__1850\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10759\
        );

    \I__1849\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10759\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__10767\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__10764\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__10759\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__1845\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10748\
        );

    \I__1844\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10745\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__10748\,
            I => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__10745\,
            I => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\
        );

    \I__1841\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10735\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10732\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10738\,
            I => \N__10729\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__10735\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__10732\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__10729\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1835\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10718\
        );

    \I__1834\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10712\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__10718\,
            I => \N__10709\
        );

    \I__1832\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10702\
        );

    \I__1831\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10702\
        );

    \I__1830\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10702\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__10712\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__10709\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__10702\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__10695\,
            I => \N__10691\
        );

    \I__1825\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10686\
        );

    \I__1824\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10686\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10682\
        );

    \I__1822\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10679\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__10682\,
            I => \N__10676\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__10679\,
            I => \N__10671\
        );

    \I__1819\ : Sp12to4
    port map (
            O => \N__10676\,
            I => \N__10671\
        );

    \I__1818\ : Odrv12
    port map (
            O => \N__10671\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__10668\,
            I => \Lab_UT.q_5_1_cascade_\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__10665\,
            I => \Lab_UT.bcd2segment1.i5_mux_cascade_\
        );

    \I__1815\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10653\
        );

    \I__1814\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10648\
        );

    \I__1813\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10648\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10645\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10640\
        );

    \I__1810\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10640\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__10656\,
            I => \N__10636\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10631\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__10648\,
            I => \N__10624\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10645\,
            I => \N__10624\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__10640\,
            I => \N__10624\
        );

    \I__1804\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10617\
        );

    \I__1803\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10617\
        );

    \I__1802\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10617\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10614\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__10631\,
            I => \N__10611\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__10624\,
            I => \N__10608\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10617\,
            I => \Lab_UT.cnt_2\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10614\,
            I => \Lab_UT.cnt_2\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__10611\,
            I => \Lab_UT.cnt_2\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__10608\,
            I => \Lab_UT.cnt_2\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__10599\,
            I => \Lab_UT.bcd2segment1.m42_amZ0_cascade_\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__10593\,
            I => \Lab_UT.bcd2segment1.m52_bmZ0\
        );

    \I__1791\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10587\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__10587\,
            I => \Lab_UT.bcd2segment1.N_42_i\
        );

    \I__1789\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10579\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10576\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10573\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__10579\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_0\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10576\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_0\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__10573\,
            I => \Lab_UT.dictrl.alarmstateZ0Z_0\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__10566\,
            I => \Lab_UT.dictrl.idle_cascade_\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10556\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10556\
        );

    \I__1780\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10553\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__10556\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__10553\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10545\
        );

    \I__1776\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10542\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__10542\,
            I => \N__10539\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__10539\,
            I => \N__10536\
        );

    \I__1773\ : Odrv4
    port map (
            O => \N__10536\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_0\
        );

    \I__1772\ : IoInMux
    port map (
            O => \N__10533\,
            I => \N__10529\
        );

    \I__1771\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10526\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10529\,
            I => \N__10523\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__10526\,
            I => \N__10520\
        );

    \I__1768\ : Span12Mux_s9_v
    port map (
            O => \N__10523\,
            I => \N__10517\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__10520\,
            I => \N__10514\
        );

    \I__1766\ : Odrv12
    port map (
            O => \N__10517\,
            I => clk
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__10514\,
            I => clk
        );

    \I__1764\ : SRMux
    port map (
            O => \N__10509\,
            I => \N__10505\
        );

    \I__1763\ : CEMux
    port map (
            O => \N__10508\,
            I => \N__10502\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10505\,
            I => \N__10499\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__10502\,
            I => \N__10496\
        );

    \I__1760\ : Span4Mux_h
    port map (
            O => \N__10499\,
            I => \N__10491\
        );

    \I__1759\ : Span4Mux_h
    port map (
            O => \N__10496\,
            I => \N__10491\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__10491\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__10488\,
            I => \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_\
        );

    \I__1756\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10482\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__10482\,
            I => \N__10479\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__10479\,
            I => \N__10476\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__10476\,
            I => \uu2.mem0.g1_2_0\
        );

    \I__1752\ : InMux
    port map (
            O => \N__10473\,
            I => \N__10470\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__10470\,
            I => \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10464\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__10464\,
            I => \uu2.mem0.g0_7_0_0_1\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__10461\,
            I => \Lab_UT.alarmchar9_cascade_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__10458\,
            I => \N__10455\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10452\
        );

    \I__1745\ : Span4Mux_h
    port map (
            O => \N__10452\,
            I => \N__10449\
        );

    \I__1744\ : Odrv4
    port map (
            O => \N__10449\,
            I => \Lab_UT.alarmcharZ0Z_2\
        );

    \I__1743\ : InMux
    port map (
            O => \N__10446\,
            I => \N__10443\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10443\,
            I => \Lab_UT.bcd2segment1.N_160\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__10440\,
            I => \uu2.mem0.N_3_0_cascade_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10437\,
            I => \N__10434\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__10434\,
            I => \uu2.mem0.N_98_0_0_0\
        );

    \I__1738\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10426\
        );

    \I__1737\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10423\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10429\,
            I => \N__10420\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__10426\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__10423\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__10420\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1732\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10407\
        );

    \I__1731\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10407\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__10407\,
            I => \uu2.N_1585_0_0\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__10404\,
            I => \Lab_UT.bcd2segment1.i6_mux_cascade_\
        );

    \I__1728\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10398\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__10398\,
            I => \Lab_UT.bcd2segment1.m68_amZ0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10392\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10392\,
            I => \N__10384\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10375\
        );

    \I__1723\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10375\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10375\
        );

    \I__1721\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10375\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10372\
        );

    \I__1719\ : Span4Mux_h
    port map (
            O => \N__10384\,
            I => \N__10369\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__10375\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__10372\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__10369\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__1715\ : IoInMux
    port map (
            O => \N__10362\,
            I => \N__10359\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__10359\,
            I => \N__10354\
        );

    \I__1713\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10351\
        );

    \I__1712\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10346\
        );

    \I__1711\ : IoSpan4Mux
    port map (
            O => \N__10354\,
            I => \N__10343\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10351\,
            I => \N__10340\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10334\
        );

    \I__1708\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10334\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10329\
        );

    \I__1706\ : Span4Mux_s1_h
    port map (
            O => \N__10343\,
            I => \N__10329\
        );

    \I__1705\ : Span4Mux_v
    port map (
            O => \N__10340\,
            I => \N__10326\
        );

    \I__1704\ : InMux
    port map (
            O => \N__10339\,
            I => \N__10323\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10318\
        );

    \I__1702\ : Span4Mux_h
    port map (
            O => \N__10329\,
            I => \N__10318\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__10326\,
            I => rst
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__10323\,
            I => rst
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__10318\,
            I => rst
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__10311\,
            I => \N__10307\
        );

    \I__1697\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10302\
        );

    \I__1696\ : InMux
    port map (
            O => \N__10307\,
            I => \N__10298\
        );

    \I__1695\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10295\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__10305\,
            I => \N__10292\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__10302\,
            I => \N__10289\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10286\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__10298\,
            I => \N__10283\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__10295\,
            I => \N__10280\
        );

    \I__1689\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10277\
        );

    \I__1688\ : Span4Mux_v
    port map (
            O => \N__10289\,
            I => \N__10274\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__10286\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__10283\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__10280\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__10277\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1683\ : Odrv4
    port map (
            O => \N__10274\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__10263\,
            I => \uu2.mem0.N_17_0_cascade_\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__10260\,
            I => \N__10257\
        );

    \I__1680\ : InMux
    port map (
            O => \N__10257\,
            I => \N__10252\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__10256\,
            I => \N__10246\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__10255\,
            I => \N__10243\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__10252\,
            I => \N__10240\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__10251\,
            I => \N__10237\
        );

    \I__1675\ : InMux
    port map (
            O => \N__10250\,
            I => \N__10230\
        );

    \I__1674\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10230\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10230\
        );

    \I__1672\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10227\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__10240\,
            I => \N__10224\
        );

    \I__1670\ : InMux
    port map (
            O => \N__10237\,
            I => \N__10221\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__10230\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__10227\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__10224\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__10221\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__1664\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__10203\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_5\
        );

    \I__1661\ : InMux
    port map (
            O => \N__10200\,
            I => \N__10197\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10194\,
            I => \uu2.mem0.N_107_0_0\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__1657\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10185\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__10185\,
            I => \uu2.mem0.N_74_0_0_1\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__10182\,
            I => \uu2.mem0.g0_7_0_0_2_cascade_\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__10179\,
            I => \Lab_UT.bcd2segment1.N_187_cascade_\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__10176\,
            I => \Lab_UT.bcd2segment1.N_189_cascade_\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10167\
        );

    \I__1651\ : InMux
    port map (
            O => \N__10172\,
            I => \N__10167\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__10167\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__1648\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10155\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10155\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__10155\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__10152\,
            I => \uu2.mem0.N_107_0_cascade_\
        );

    \I__1644\ : InMux
    port map (
            O => \N__10149\,
            I => \N__10143\
        );

    \I__1643\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10140\
        );

    \I__1642\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10135\
        );

    \I__1641\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10135\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__10143\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__10140\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__10135\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__10128\,
            I => \N__10125\
        );

    \I__1636\ : InMux
    port map (
            O => \N__10125\,
            I => \N__10122\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__10122\,
            I => \N__10119\
        );

    \I__1634\ : Span4Mux_s3_h
    port map (
            O => \N__10119\,
            I => \N__10116\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__10116\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_1\
        );

    \I__1632\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10110\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10106\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__10109\,
            I => \N__10102\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__10106\,
            I => \N__10099\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10094\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10094\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__10099\,
            I => \L3_tx_data_6\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10094\,
            I => \L3_tx_data_6\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__10089\,
            I => \uu2.mem0.N_130_mux_cascade_\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10080\
        );

    \I__1621\ : Span4Mux_h
    port map (
            O => \N__10080\,
            I => \N__10077\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__10077\,
            I => \uu2.mem0.N_54_0_i\
        );

    \I__1619\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10070\
        );

    \I__1618\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10066\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__10070\,
            I => \N__10063\
        );

    \I__1616\ : InMux
    port map (
            O => \N__10069\,
            I => \N__10060\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__10066\,
            I => \N__10052\
        );

    \I__1614\ : Span4Mux_v
    port map (
            O => \N__10063\,
            I => \N__10052\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__10060\,
            I => \N__10052\
        );

    \I__1612\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10049\
        );

    \I__1611\ : Span4Mux_h
    port map (
            O => \N__10052\,
            I => \N__10046\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__10049\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__10046\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1608\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10036\
        );

    \I__1607\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10031\
        );

    \I__1606\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10031\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__10036\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__10031\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10021\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10016\
        );

    \I__1601\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10016\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10021\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__10016\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10011\,
            I => \N__10008\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__10008\,
            I => \N__10004\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10007\,
            I => \N__10001\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__10004\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10001\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1593\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9993\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9990\
        );

    \I__1591\ : Span4Mux_h
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__9987\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__9984\,
            I => \N__9981\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9977\
        );

    \I__1587\ : InMux
    port map (
            O => \N__9980\,
            I => \N__9974\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9977\,
            I => \uu2.un284_ci\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__9974\,
            I => \uu2.un284_ci\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__9969\,
            I => \N__9962\
        );

    \I__1583\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9959\
        );

    \I__1582\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9956\
        );

    \I__1581\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9951\
        );

    \I__1580\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9951\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9948\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__9959\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__9956\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__9951\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__9948\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9936\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__9936\,
            I => \N__9933\
        );

    \I__1572\ : Span4Mux_h
    port map (
            O => \N__9933\,
            I => \N__9930\
        );

    \I__1571\ : IoSpan4Mux
    port map (
            O => \N__9930\,
            I => \N__9927\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__9927\,
            I => \uart_RXD\
        );

    \I__1569\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9920\
        );

    \I__1568\ : InMux
    port map (
            O => \N__9923\,
            I => \N__9917\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9914\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9917\,
            I => \uu2.un350_ci\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__9914\,
            I => \uu2.un350_ci\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__9909\,
            I => \N__9904\
        );

    \I__1563\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9901\
        );

    \I__1562\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9898\
        );

    \I__1561\ : InMux
    port map (
            O => \N__9904\,
            I => \N__9895\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__9901\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__9898\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9895\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__9888\,
            I => \N__9885\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9880\
        );

    \I__1555\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9875\
        );

    \I__1554\ : InMux
    port map (
            O => \N__9883\,
            I => \N__9875\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__9880\,
            I => \N__9868\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9868\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9863\
        );

    \I__1550\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9863\
        );

    \I__1549\ : Span4Mux_h
    port map (
            O => \N__9868\,
            I => \N__9860\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9857\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__9860\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__9857\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__1545\ : CEMux
    port map (
            O => \N__9852\,
            I => \N__9849\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9846\
        );

    \I__1543\ : Sp12to4
    port map (
            O => \N__9846\,
            I => \N__9843\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__9843\,
            I => \Lab_UT.dictrl.G_74\
        );

    \I__1541\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9833\
        );

    \I__1540\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9833\
        );

    \I__1539\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9830\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__9833\,
            I => \N__9822\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9822\
        );

    \I__1536\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9815\
        );

    \I__1535\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9815\
        );

    \I__1534\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9815\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__9822\,
            I => \Lab_UT.dictrl.un1_next_alarmstate21_0\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__9815\,
            I => \Lab_UT.dictrl.un1_next_alarmstate21_0\
        );

    \I__1531\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9806\
        );

    \I__1530\ : InMux
    port map (
            O => \N__9809\,
            I => \N__9803\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9798\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__9803\,
            I => \N__9798\
        );

    \I__1527\ : Span12Mux_s9_v
    port map (
            O => \N__9798\,
            I => \N__9792\
        );

    \I__1526\ : InMux
    port map (
            O => \N__9797\,
            I => \N__9785\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9785\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9795\,
            I => \N__9785\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__9792\,
            I => \Lab_UT.cnt_0\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__9785\,
            I => \Lab_UT.cnt_0\
        );

    \I__1521\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9771\
        );

    \I__1520\ : InMux
    port map (
            O => \N__9779\,
            I => \N__9771\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9778\,
            I => \N__9768\
        );

    \I__1518\ : InMux
    port map (
            O => \N__9777\,
            I => \N__9763\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9776\,
            I => \N__9763\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__9771\,
            I => \N__9760\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__9768\,
            I => \uu2.un306_ci\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9763\,
            I => \uu2.un306_ci\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__9760\,
            I => \uu2.un306_ci\
        );

    \I__1512\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9750\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__9750\,
            I => \N__9743\
        );

    \I__1510\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9738\
        );

    \I__1509\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9738\
        );

    \I__1508\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9733\
        );

    \I__1507\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9733\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__9743\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__9738\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__9733\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1503\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9723\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__9723\,
            I => \N__9716\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9722\,
            I => \N__9709\
        );

    \I__1500\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9709\
        );

    \I__1499\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9709\
        );

    \I__1498\ : InMux
    port map (
            O => \N__9719\,
            I => \N__9706\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__9716\,
            I => \N__9696\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9691\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__9706\,
            I => \N__9691\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9686\
        );

    \I__1493\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9686\
        );

    \I__1492\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9679\
        );

    \I__1491\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9679\
        );

    \I__1490\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9679\
        );

    \I__1489\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9674\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9699\,
            I => \N__9674\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__9696\,
            I => \uu0.un4_l_count_0\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__9691\,
            I => \uu0.un4_l_count_0\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__9686\,
            I => \uu0.un4_l_count_0\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__9679\,
            I => \uu0.un4_l_count_0\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__9674\,
            I => \uu0.un4_l_count_0\
        );

    \I__1482\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9660\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__9660\,
            I => \N__9656\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9653\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__9656\,
            I => \N__9647\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9647\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9644\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__9647\,
            I => \N__9638\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9638\
        );

    \I__1474\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9635\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__9638\,
            I => \N__9632\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__9635\,
            I => \o_One_Sec_Pulse\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__9632\,
            I => \o_One_Sec_Pulse\
        );

    \I__1470\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__1468\ : Odrv4
    port map (
            O => \N__9621\,
            I => \Lab_UT.bcd2segment1.m59_bmZ0\
        );

    \I__1467\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__9615\,
            I => \Lab_UT.bcd2segment1.m52_amZ0\
        );

    \I__1465\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9609\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__9606\,
            I => \Lab_UT.alarmcharZ0Z_0\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__9603\,
            I => \N__9600\
        );

    \I__1461\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9594\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9591\
        );

    \I__1458\ : Span4Mux_h
    port map (
            O => \N__9591\,
            I => \N__9587\
        );

    \I__1457\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9584\
        );

    \I__1456\ : Odrv4
    port map (
            O => \N__9587\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9584\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0\
        );

    \I__1454\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9573\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9573\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__9573\,
            I => \N__9570\
        );

    \I__1451\ : Span4Mux_h
    port map (
            O => \N__9570\,
            I => \N__9565\
        );

    \I__1450\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9562\
        );

    \I__1449\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9559\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__9565\,
            I => \Lab_UT.dictrl.next_alarmstate_1\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__9562\,
            I => \Lab_UT.dictrl.next_alarmstate_1\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__9559\,
            I => \Lab_UT.dictrl.next_alarmstate_1\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__9552\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9546\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__9546\,
            I => \N__9543\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__9543\,
            I => \Lab_UT.bcd2segment1.m59_amZ0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9537\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__9537\,
            I => \Lab_UT.bcd2segment1.m68_bmZ0\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9531\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__9531\,
            I => \uu2.un28_w_addr_user_i_0_a2Z0Z_4\
        );

    \I__1437\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9525\,
            I => \N__9520\
        );

    \I__1435\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9517\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9514\
        );

    \I__1433\ : Odrv4
    port map (
            O => \N__9520\,
            I => \L3_tx_data_3\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__9517\,
            I => \L3_tx_data_3\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__9514\,
            I => \L3_tx_data_3\
        );

    \I__1430\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9503\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__9506\,
            I => \N__9499\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9496\
        );

    \I__1427\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9493\
        );

    \I__1426\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9490\
        );

    \I__1425\ : Odrv4
    port map (
            O => \N__9496\,
            I => \L3_tx_data_4\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__9493\,
            I => \L3_tx_data_4\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9490\,
            I => \L3_tx_data_4\
        );

    \I__1422\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9478\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9475\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9472\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__9478\,
            I => \L3_tx_data_0\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__9475\,
            I => \L3_tx_data_0\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__9472\,
            I => \L3_tx_data_0\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__9465\,
            I => \uu2.w_data_i_o2_4Z0Z_0_cascade_\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__9462\,
            I => \N_96_cascade_\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__9459\,
            I => \uu2.un21_w_addr_displaying_i_cascade_\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__9456\,
            I => \N__9453\
        );

    \I__1412\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9450\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9450\,
            I => \N__9447\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__9447\,
            I => \N__9444\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__9444\,
            I => \Lab_UT.alarmcharZ0Z_5\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__9438\,
            I => \uu2.mem0.N_13_1_0_0\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__9435\,
            I => \uu2.mem0.i14_mux_0_0_0_cascade_\
        );

    \I__1405\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9429\,
            I => \uu2.mem0.N_8_0_0_1\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__1402\ : InMux
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__9420\,
            I => \Lab_UT.alarmcharZ0Z_6\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__9417\,
            I => \N__9413\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__9416\,
            I => \N__9410\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9405\
        );

    \I__1397\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9405\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__9405\,
            I => \N__9401\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9398\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__9401\,
            I => \uu2.N_155\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9398\,
            I => \uu2.N_155\
        );

    \I__1392\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9386\
        );

    \I__1391\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9386\
        );

    \I__1390\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9383\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9386\,
            I => \uu2.N_106\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__9383\,
            I => \uu2.N_106\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__9378\,
            I => \N__9373\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9369\
        );

    \I__1385\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9366\
        );

    \I__1384\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9361\
        );

    \I__1383\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9361\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__9369\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__9366\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__9361\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__9354\,
            I => \N__9351\
        );

    \I__1378\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9348\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__9348\,
            I => \N__9343\
        );

    \I__1376\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9340\
        );

    \I__1375\ : InMux
    port map (
            O => \N__9346\,
            I => \N__9337\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__9343\,
            I => \uu2.N_102\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__9340\,
            I => \uu2.N_102\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__9337\,
            I => \uu2.N_102\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__9330\,
            I => \N__9326\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__9329\,
            I => \N__9321\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9317\
        );

    \I__1368\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9312\
        );

    \I__1367\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9312\
        );

    \I__1366\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9309\
        );

    \I__1365\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9305\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__9317\,
            I => \N__9302\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9297\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__9309\,
            I => \N__9297\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9294\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__9305\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__9302\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1358\ : Odrv12
    port map (
            O => \N__9297\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__9294\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1356\ : InMux
    port map (
            O => \N__9285\,
            I => \N__9276\
        );

    \I__1355\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9265\
        );

    \I__1354\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9265\
        );

    \I__1353\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9265\
        );

    \I__1352\ : InMux
    port map (
            O => \N__9281\,
            I => \N__9265\
        );

    \I__1351\ : InMux
    port map (
            O => \N__9280\,
            I => \N__9265\
        );

    \I__1350\ : CascadeMux
    port map (
            O => \N__9279\,
            I => \N__9262\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__9276\,
            I => \N__9254\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9265\,
            I => \N__9254\
        );

    \I__1347\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9245\
        );

    \I__1346\ : InMux
    port map (
            O => \N__9261\,
            I => \N__9245\
        );

    \I__1345\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9245\
        );

    \I__1344\ : InMux
    port map (
            O => \N__9259\,
            I => \N__9245\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__9254\,
            I => \uu2.N_97\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__9245\,
            I => \uu2.N_97\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__1340\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9228\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9228\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9225\
        );

    \I__1337\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9222\
        );

    \I__1336\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9219\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__9228\,
            I => \N__9216\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__9225\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__9222\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__9219\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__9216\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__1330\ : CEMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1328\ : Span4Mux_v
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__1327\ : Span4Mux_s2_v
    port map (
            O => \N__9198\,
            I => \N__9195\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__9195\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__1325\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9189\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9186\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__9186\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_12\
        );

    \I__1322\ : CascadeMux
    port map (
            O => \N__9183\,
            I => \uu2.N_41_0_cascade_\
        );

    \I__1321\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9177\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__9177\,
            I => \uu2.N_132_mux\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__9174\,
            I => \uu2.N_132_mux_cascade_\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9168\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__1316\ : Span4Mux_h
    port map (
            O => \N__9165\,
            I => \N__9162\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__9162\,
            I => \uu2.mem0.N_94_i\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__1313\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9153\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__9153\,
            I => \N__9149\
        );

    \I__1311\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9146\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__9149\,
            I => \N__9143\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__9146\,
            I => \uu2.N_15_i\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__9143\,
            I => \uu2.N_15_i\
        );

    \I__1307\ : InMux
    port map (
            O => \N__9138\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9135\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__9132\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__1304\ : InMux
    port map (
            O => \N__9129\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__1302\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9117\
        );

    \I__1301\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9117\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__9117\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__1298\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9105\
        );

    \I__1297\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9105\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__9105\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__9102\,
            I => \N__9098\
        );

    \I__1294\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9095\
        );

    \I__1293\ : InMux
    port map (
            O => \N__9098\,
            I => \N__9092\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__9095\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9092\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__9087\,
            I => \N__9084\
        );

    \I__1289\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9078\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9083\,
            I => \N__9078\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__9078\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__1286\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9069\
        );

    \I__1285\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9069\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__9069\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__1283\ : InMux
    port map (
            O => \N__9066\,
            I => \N__9058\
        );

    \I__1282\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9058\
        );

    \I__1281\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9055\
        );

    \I__1280\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9052\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__9058\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__9055\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__9052\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__9045\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__9042\,
            I => \N__9038\
        );

    \I__1274\ : InMux
    port map (
            O => \N__9041\,
            I => \N__9034\
        );

    \I__1273\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9029\
        );

    \I__1272\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9029\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__9034\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9029\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__1269\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9018\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9011\
        );

    \I__1267\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9011\
        );

    \I__1266\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9011\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__9008\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__9011\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__9008\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__9000\,
            I => \N__8995\
        );

    \I__1260\ : CascadeMux
    port map (
            O => \N__8999\,
            I => \N__8992\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__8998\,
            I => \N__8989\
        );

    \I__1258\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8982\
        );

    \I__1257\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8982\
        );

    \I__1256\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8982\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__8982\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__8979\,
            I => \N__8975\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8971\
        );

    \I__1252\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8966\
        );

    \I__1251\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8966\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__8971\,
            I => \N__8963\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8966\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__8963\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8958\,
            I => \N__8952\
        );

    \I__1246\ : InMux
    port map (
            O => \N__8957\,
            I => \N__8952\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__8952\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__1244\ : InMux
    port map (
            O => \N__8949\,
            I => \N__8940\
        );

    \I__1243\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8940\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8937\
        );

    \I__1241\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8932\
        );

    \I__1240\ : InMux
    port map (
            O => \N__8945\,
            I => \N__8932\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__8940\,
            I => \N__8929\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__8937\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__8932\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__8929\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8914\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8914\
        );

    \I__1233\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8907\
        );

    \I__1232\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8907\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__8914\,
            I => \N__8904\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8899\
        );

    \I__1229\ : InMux
    port map (
            O => \N__8912\,
            I => \N__8899\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__8907\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__8904\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__8899\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1225\ : InMux
    port map (
            O => \N__8892\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8889\,
            I => \N__8878\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__8888\,
            I => \N__8875\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8853\
        );

    \I__1221\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8853\
        );

    \I__1220\ : InMux
    port map (
            O => \N__8885\,
            I => \N__8853\
        );

    \I__1219\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8853\
        );

    \I__1218\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8853\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8882\,
            I => \N__8853\
        );

    \I__1216\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8853\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__8878\,
            I => \N__8850\
        );

    \I__1214\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8845\
        );

    \I__1213\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8845\
        );

    \I__1212\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8838\
        );

    \I__1211\ : InMux
    port map (
            O => \N__8872\,
            I => \N__8838\
        );

    \I__1210\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8838\
        );

    \I__1209\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8835\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8832\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__8868\,
            I => \N__8829\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__8853\,
            I => \N__8826\
        );

    \I__1205\ : Span4Mux_s2_h
    port map (
            O => \N__8850\,
            I => \N__8821\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__8845\,
            I => \N__8821\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__8838\,
            I => \N__8818\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8813\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__8832\,
            I => \N__8813\
        );

    \I__1200\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8810\
        );

    \I__1199\ : Span4Mux_s3_h
    port map (
            O => \N__8826\,
            I => \N__8807\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__8821\,
            I => \N__8804\
        );

    \I__1197\ : Span4Mux_s3_h
    port map (
            O => \N__8818\,
            I => \N__8801\
        );

    \I__1196\ : Span4Mux_h
    port map (
            O => \N__8813\,
            I => \N__8798\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__8810\,
            I => vbuf_tx_data_rdy
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__8807\,
            I => vbuf_tx_data_rdy
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__8804\,
            I => vbuf_tx_data_rdy
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__8801\,
            I => vbuf_tx_data_rdy
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__8798\,
            I => vbuf_tx_data_rdy
        );

    \I__1190\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8783\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__8786\,
            I => \N__8780\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8775\
        );

    \I__1187\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8770\
        );

    \I__1186\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8770\
        );

    \I__1185\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8767\
        );

    \I__1184\ : Odrv4
    port map (
            O => \N__8775\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8770\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__8767\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1181\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8757\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__8757\,
            I => \N__8751\
        );

    \I__1179\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8746\
        );

    \I__1178\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8743\
        );

    \I__1177\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8740\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__8751\,
            I => \N__8737\
        );

    \I__1175\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8732\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8732\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__8746\,
            I => \N__8727\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__8743\,
            I => \N__8727\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__8740\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__8737\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__8732\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1168\ : Odrv4
    port map (
            O => \N__8727\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1167\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8715\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__8715\,
            I => \N__8711\
        );

    \I__1165\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8705\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__8711\,
            I => \N__8702\
        );

    \I__1163\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8697\
        );

    \I__1162\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8697\
        );

    \I__1161\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8694\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__8705\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__8702\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__8697\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8694\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1156\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8682\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__1154\ : Span4Mux_s3_h
    port map (
            O => \N__8679\,
            I => \N__8676\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__8676\,
            I => \uu0.un143_ci_0\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__8673\,
            I => \uu2.un1_l_count_1_2_0_cascade_\
        );

    \I__1151\ : InMux
    port map (
            O => \N__8670\,
            I => \N__8666\
        );

    \I__1150\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8663\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8660\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8655\
        );

    \I__1147\ : Span4Mux_s3_h
    port map (
            O => \N__8660\,
            I => \N__8655\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__8655\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__8652\,
            I => \uu2.un1_l_count_2_2_cascade_\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__8649\,
            I => \resetGen.reset_count_2_0_4_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8646\,
            I => \N__8643\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__8643\,
            I => \N__8640\
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__8640\,
            I => \Lab_UT.alarmchar10\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1139\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8631\,
            I => \Lab_UT.alarmcharZ0Z_4\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__8628\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__1136\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8621\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8618\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__8621\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__8618\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8606\
        );

    \I__1131\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8606\
        );

    \I__1130\ : InMux
    port map (
            O => \N__8611\,
            I => \N__8603\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__8606\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__8603\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1127\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__8595\,
            I => \resetGen.un241_ci\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__8592\,
            I => \resetGen.un241_ci_cascade_\
        );

    \I__1124\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8584\
        );

    \I__1123\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8581\
        );

    \I__1122\ : InMux
    port map (
            O => \N__8587\,
            I => \N__8578\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__8584\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__8581\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8578\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__1117\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8556\
        );

    \I__1116\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8556\
        );

    \I__1115\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8556\
        );

    \I__1114\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8556\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__8556\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__8553\,
            I => \uu2.un28_w_addr_user_i_0_cascade_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8547\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8547\,
            I => \N__8541\
        );

    \I__1109\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8536\
        );

    \I__1108\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8536\
        );

    \I__1107\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8533\
        );

    \I__1106\ : Odrv4
    port map (
            O => \N__8541\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__8536\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8533\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__1103\ : InMux
    port map (
            O => \N__8526\,
            I => \N__8523\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8523\,
            I => \N__8520\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__8520\,
            I => \uu2.N_105\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__1099\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8508\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8503\
        );

    \I__1097\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8503\
        );

    \I__1096\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8500\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8495\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8503\,
            I => \N__8495\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__8500\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__8495\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__8490\,
            I => \uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_\
        );

    \I__1090\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8484\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8481\
        );

    \I__1088\ : Odrv4
    port map (
            O => \N__8481\,
            I => \Lab_UT.alarmchar_2_1_1\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__8478\,
            I => \N__8475\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__8472\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_4\
        );

    \I__1084\ : InMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__8466\,
            I => \uu2.w_addr_user_3_i_a2_3_6\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \uu2.mem0.g1_3_0_cascade_\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8457\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__8457\,
            I => \uu2.mem0.N_63_0_i\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8451\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__8451\,
            I => \uu2.mem0.G_17_0_0_0\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__8448\,
            I => \N__8444\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__8447\,
            I => \N__8441\
        );

    \I__1075\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8436\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8436\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__8436\,
            I => \N_72_mux\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8430\
        );

    \I__1071\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__1069\ : Span4Mux_s3_h
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__1068\ : Odrv4
    port map (
            O => \N__8421\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_3\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8415\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__8415\,
            I => \uu2.w_addr_user_3_i_a2_2_6\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1064\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__8406\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_2\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1061\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__8397\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_6\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__8394\,
            I => \N__8391\
        );

    \I__1058\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8388\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8388\,
            I => \N__8385\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__8385\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_7\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__8382\,
            I => \uu2.N_102_cascade_\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__8379\,
            I => \N__8376\
        );

    \I__1053\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__8373\,
            I => \uu2.N_61_i\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__8370\,
            I => \N__8364\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8361\
        );

    \I__1049\ : InMux
    port map (
            O => \N__8368\,
            I => \N__8358\
        );

    \I__1048\ : InMux
    port map (
            O => \N__8367\,
            I => \N__8351\
        );

    \I__1047\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8351\
        );

    \I__1046\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8351\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__8358\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8351\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__8346\,
            I => \buart.Z_tx.un1_bitcount_c3_cascade_\
        );

    \I__1042\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8339\
        );

    \I__1041\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8336\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__8339\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__8336\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__8331\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8321\
        );

    \I__1036\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8318\
        );

    \I__1035\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8311\
        );

    \I__1034\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8311\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8311\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__8321\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__8318\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8311\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1029\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8292\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8292\
        );

    \I__1027\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8292\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8292\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__8292\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__8289\,
            I => \N__8284\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8279\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8274\
        );

    \I__1021\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8274\
        );

    \I__1020\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8269\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8269\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8279\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__8274\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__8269\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__8262\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__8259\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\
        );

    \I__1013\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8247\
        );

    \I__1012\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8247\
        );

    \I__1011\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8247\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__8247\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8241\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__8241\,
            I => \N__8238\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__8238\,
            I => \N__8235\
        );

    \I__1006\ : Span4Mux_v
    port map (
            O => \N__8235\,
            I => \N__8232\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__8232\,
            I => \Lab_UT.alarmchar10_i_2\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__8229\,
            I => \N__8224\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8219\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8219\
        );

    \I__1001\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8216\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8219\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__8216\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__8211\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__997\ : InMux
    port map (
            O => \N__8208\,
            I => \N__8204\
        );

    \I__996\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8201\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__8204\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__8201\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__993\ : CEMux
    port map (
            O => \N__8196\,
            I => \N__8181\
        );

    \I__992\ : CEMux
    port map (
            O => \N__8195\,
            I => \N__8181\
        );

    \I__991\ : CEMux
    port map (
            O => \N__8194\,
            I => \N__8181\
        );

    \I__990\ : CEMux
    port map (
            O => \N__8193\,
            I => \N__8181\
        );

    \I__989\ : CEMux
    port map (
            O => \N__8192\,
            I => \N__8181\
        );

    \I__988\ : GlobalMux
    port map (
            O => \N__8181\,
            I => \N__8178\
        );

    \I__987\ : gio2CtrlBuf
    port map (
            O => \N__8178\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__8175\,
            I => \N__8170\
        );

    \I__985\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8165\
        );

    \I__984\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8165\
        );

    \I__983\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8162\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8165\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__8162\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__979\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8141\
        );

    \I__978\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8141\
        );

    \I__977\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8141\
        );

    \I__976\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8141\
        );

    \I__975\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8138\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__8141\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__8138\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__972\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8123\
        );

    \I__971\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8123\
        );

    \I__970\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8123\
        );

    \I__969\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8120\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__8123\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__8120\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__966\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8109\
        );

    \I__965\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8100\
        );

    \I__964\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8100\
        );

    \I__963\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8100\
        );

    \I__962\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8100\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__8100\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__960\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8081\
        );

    \I__959\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8081\
        );

    \I__958\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8081\
        );

    \I__957\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8081\
        );

    \I__956\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8081\
        );

    \I__955\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8078\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__8081\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__8078\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__8073\,
            I => \N__8070\
        );

    \I__951\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8062\
        );

    \I__950\ : InMux
    port map (
            O => \N__8069\,
            I => \N__8062\
        );

    \I__949\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8059\
        );

    \I__948\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8056\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8051\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__8059\,
            I => \N__8051\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__8056\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__8051\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__8046\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__942\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8033\
        );

    \I__941\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8033\
        );

    \I__940\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8033\
        );

    \I__939\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8030\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__8033\,
            I => \N__8027\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__8030\,
            I => \N__8024\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__8027\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__8024\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__934\ : InMux
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__8016\,
            I => \uu0.un4_l_count_18\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__8013\,
            I => \N__8006\
        );

    \I__931\ : InMux
    port map (
            O => \N__8012\,
            I => \N__7992\
        );

    \I__930\ : InMux
    port map (
            O => \N__8011\,
            I => \N__7992\
        );

    \I__929\ : InMux
    port map (
            O => \N__8010\,
            I => \N__7992\
        );

    \I__928\ : InMux
    port map (
            O => \N__8009\,
            I => \N__7992\
        );

    \I__927\ : InMux
    port map (
            O => \N__8006\,
            I => \N__7992\
        );

    \I__926\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7992\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__7992\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__924\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7985\
        );

    \I__923\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7982\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__7985\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__7982\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__920\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__7974\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__918\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7967\
        );

    \I__917\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__7967\,
            I => \N__7961\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7964\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__7961\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__913\ : InMux
    port map (
            O => \N__7956\,
            I => \N__7953\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7950\
        );

    \I__911\ : Odrv4
    port map (
            O => \N__7950\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__910\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__7944\,
            I => \uu0.un55_ci\
        );

    \I__908\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7936\
        );

    \I__907\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7933\
        );

    \I__906\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7930\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__7936\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__7933\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__7930\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7919\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7916\
        );

    \I__900\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7912\
        );

    \I__899\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7909\
        );

    \I__898\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7906\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__7912\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__7909\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7906\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__7899\,
            I => \N__7891\
        );

    \I__893\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7881\
        );

    \I__892\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7881\
        );

    \I__891\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7876\
        );

    \I__890\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7876\
        );

    \I__889\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7871\
        );

    \I__888\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7871\
        );

    \I__887\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7868\
        );

    \I__886\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7859\
        );

    \I__885\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7859\
        );

    \I__884\ : InMux
    port map (
            O => \N__7887\,
            I => \N__7859\
        );

    \I__883\ : InMux
    port map (
            O => \N__7886\,
            I => \N__7859\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7854\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7876\,
            I => \N__7854\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__7871\,
            I => \uu0.un110_ci\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7868\,
            I => \uu0.un110_ci\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__7859\,
            I => \uu0.un110_ci\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__7854\,
            I => \uu0.un110_ci\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__7845\,
            I => \N__7841\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__7844\,
            I => \N__7837\
        );

    \I__874\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7834\
        );

    \I__873\ : InMux
    port map (
            O => \N__7840\,
            I => \N__7829\
        );

    \I__872\ : InMux
    port map (
            O => \N__7837\,
            I => \N__7829\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__7834\,
            I => \uu0.un198_ci_2\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7829\,
            I => \uu0.un198_ci_2\
        );

    \I__869\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7820\
        );

    \I__868\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7817\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__7820\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__7817\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__865\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7807\
        );

    \I__864\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7802\
        );

    \I__863\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7802\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__7807\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__7802\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__859\ : InMux
    port map (
            O => \N__7794\,
            I => \N__7790\
        );

    \I__858\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7785\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__7790\,
            I => \N__7782\
        );

    \I__856\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7777\
        );

    \I__855\ : InMux
    port map (
            O => \N__7788\,
            I => \N__7777\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__7785\,
            I => \N__7774\
        );

    \I__853\ : Odrv12
    port map (
            O => \N__7782\,
            I => \uu0.un154_ci_9\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7777\,
            I => \uu0.un154_ci_9\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__7774\,
            I => \uu0.un154_ci_9\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__7767\,
            I => \N__7764\
        );

    \I__849\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7761\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__7761\,
            I => \uu0.un165_ci_0\
        );

    \I__847\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7755\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__7755\,
            I => \N__7752\
        );

    \I__845\ : Span4Mux_h
    port map (
            O => \N__7752\,
            I => \N__7749\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__7749\,
            I => \uu0.sec_clkDZ0\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__7746\,
            I => \N__7743\
        );

    \I__842\ : InMux
    port map (
            O => \N__7743\,
            I => \N__7738\
        );

    \I__841\ : InMux
    port map (
            O => \N__7742\,
            I => \N__7732\
        );

    \I__840\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7732\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__7738\,
            I => \N__7729\
        );

    \I__838\ : InMux
    port map (
            O => \N__7737\,
            I => \N__7726\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__7732\,
            I => \N__7723\
        );

    \I__836\ : Odrv4
    port map (
            O => \N__7729\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__7726\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__7723\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__7716\,
            I => \N__7711\
        );

    \I__832\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7705\
        );

    \I__831\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7705\
        );

    \I__830\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7700\
        );

    \I__829\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7700\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__7705\,
            I => \N__7697\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7694\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__7697\,
            I => \uu2.un404_ci\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__7694\,
            I => \uu2.un404_ci\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__823\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7679\
        );

    \I__822\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7674\
        );

    \I__821\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7674\
        );

    \I__820\ : InMux
    port map (
            O => \N__7683\,
            I => \N__7669\
        );

    \I__819\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7669\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__7679\,
            I => \N__7664\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__7674\,
            I => \N__7664\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__7669\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__7664\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__814\ : CEMux
    port map (
            O => \N__7659\,
            I => \N__7656\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7656\,
            I => \N__7652\
        );

    \I__812\ : CEMux
    port map (
            O => \N__7655\,
            I => \N__7649\
        );

    \I__811\ : Span4Mux_h
    port map (
            O => \N__7652\,
            I => \N__7644\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7644\
        );

    \I__809\ : Sp12to4
    port map (
            O => \N__7644\,
            I => \N__7641\
        );

    \I__808\ : Odrv12
    port map (
            O => \N__7641\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__7638\,
            I => \N__7635\
        );

    \I__806\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7631\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__7634\,
            I => \N__7627\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7624\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__7630\,
            I => \N__7621\
        );

    \I__802\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7618\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__7624\,
            I => \N__7615\
        );

    \I__800\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7612\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__7618\,
            I => \N__7609\
        );

    \I__798\ : Odrv4
    port map (
            O => \N__7615\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__7612\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__796\ : Odrv4
    port map (
            O => \N__7609\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__7602\,
            I => \uu2.un404_ci_cascade_\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__793\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7592\
        );

    \I__792\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7588\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7592\,
            I => \N__7585\
        );

    \I__790\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7582\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__7588\,
            I => \N__7579\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__7585\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__7582\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__786\ : Odrv4
    port map (
            O => \N__7579\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__7572\,
            I => \N__7568\
        );

    \I__784\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__783\ : InMux
    port map (
            O => \N__7568\,
            I => \N__7560\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__7565\,
            I => \N__7557\
        );

    \I__781\ : InMux
    port map (
            O => \N__7564\,
            I => \N__7552\
        );

    \I__780\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7552\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__7560\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__778\ : Odrv4
    port map (
            O => \N__7557\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__7552\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__776\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__7542\,
            I => \N__7539\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__7539\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__773\ : InMux
    port map (
            O => \N__7536\,
            I => \N__7533\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__7533\,
            I => \N__7530\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__7530\,
            I => vbuf_tx_data_5
        );

    \I__770\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7524\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__7524\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__768\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__766\ : Odrv4
    port map (
            O => \N__7515\,
            I => vbuf_tx_data_6
        );

    \I__765\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__7509\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__763\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__7503\,
            I => \N__7500\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__7500\,
            I => vbuf_tx_data_7
        );

    \I__760\ : InMux
    port map (
            O => \N__7497\,
            I => \N__7494\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__7491\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__757\ : CEMux
    port map (
            O => \N__7488\,
            I => \N__7485\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7485\,
            I => \N__7481\
        );

    \I__755\ : CEMux
    port map (
            O => \N__7484\,
            I => \N__7478\
        );

    \I__754\ : Span4Mux_v
    port map (
            O => \N__7481\,
            I => \N__7475\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7472\
        );

    \I__752\ : Span4Mux_s1_h
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__750\ : Odrv4
    port map (
            O => \N__7469\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__749\ : Odrv4
    port map (
            O => \N__7466\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__748\ : CEMux
    port map (
            O => \N__7461\,
            I => \N__7458\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__7458\,
            I => \N__7454\
        );

    \I__746\ : CEMux
    port map (
            O => \N__7457\,
            I => \N__7451\
        );

    \I__745\ : Span4Mux_v
    port map (
            O => \N__7454\,
            I => \N__7448\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7445\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__7448\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__742\ : Odrv12
    port map (
            O => \N__7445\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__741\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7437\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__7437\,
            I => \uu2.r_data_wire_0\
        );

    \I__739\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__7431\,
            I => vbuf_tx_data_0
        );

    \I__737\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7425\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__7425\,
            I => \N__7422\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__7422\,
            I => \uu2.r_data_wire_1\
        );

    \I__734\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7416\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__7416\,
            I => vbuf_tx_data_1
        );

    \I__732\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7410\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__7410\,
            I => \uu2.r_data_wire_2\
        );

    \I__730\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__7404\,
            I => vbuf_tx_data_2
        );

    \I__728\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7398\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__7398\,
            I => \uu2.r_data_wire_3\
        );

    \I__726\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7392\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__7392\,
            I => vbuf_tx_data_3
        );

    \I__724\ : InMux
    port map (
            O => \N__7389\,
            I => \N__7386\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7386\,
            I => \uu2.r_data_wire_5\
        );

    \I__722\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__7380\,
            I => \uu2.r_data_wire_6\
        );

    \I__720\ : InMux
    port map (
            O => \N__7377\,
            I => \N__7374\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__7374\,
            I => \uu2.r_data_wire_7\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__7371\,
            I => \N__7368\
        );

    \I__717\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7362\
        );

    \I__716\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7362\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__7362\,
            I => \N__7359\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__7359\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__713\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7351\
        );

    \I__712\ : InMux
    port map (
            O => \N__7355\,
            I => \N__7348\
        );

    \I__711\ : InMux
    port map (
            O => \N__7354\,
            I => \N__7345\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__7351\,
            I => \N__7339\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7339\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__7345\,
            I => \N__7336\
        );

    \I__707\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7333\
        );

    \I__706\ : Odrv12
    port map (
            O => \N__7339\,
            I => \uu0.un66_ci\
        );

    \I__705\ : Odrv4
    port map (
            O => \N__7336\,
            I => \uu0.un66_ci\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__7333\,
            I => \uu0.un66_ci\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__7326\,
            I => \N__7322\
        );

    \I__702\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7319\
        );

    \I__701\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7316\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7311\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__7316\,
            I => \N__7311\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__7311\,
            I => \uu0.un88_ci_3\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__7308\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__696\ : InMux
    port map (
            O => \N__7305\,
            I => \N__7301\
        );

    \I__695\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7296\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__7301\,
            I => \N__7293\
        );

    \I__693\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7288\
        );

    \I__692\ : InMux
    port map (
            O => \N__7299\,
            I => \N__7288\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__7296\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__690\ : Odrv12
    port map (
            O => \N__7293\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7288\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__688\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7276\
        );

    \I__687\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7271\
        );

    \I__686\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7271\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__7276\,
            I => \N__7268\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__7271\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__683\ : Odrv12
    port map (
            O => \N__7268\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__7263\,
            I => \N__7257\
        );

    \I__681\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7247\
        );

    \I__680\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7247\
        );

    \I__679\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7247\
        );

    \I__678\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7247\
        );

    \I__677\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7244\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__7247\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__7244\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__674\ : InMux
    port map (
            O => \N__7239\,
            I => \N__7236\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__672\ : Odrv4
    port map (
            O => \N__7233\,
            I => \uu0.un4_l_count_12\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__7230\,
            I => \N__7227\
        );

    \I__670\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7223\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__7226\,
            I => \N__7220\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__7223\,
            I => \N__7217\
        );

    \I__667\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7214\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__7217\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__7214\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__7209\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__663\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7196\
        );

    \I__662\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7196\
        );

    \I__661\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7196\
        );

    \I__660\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7193\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__7196\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__7193\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__7188\,
            I => \N__7183\
        );

    \I__656\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7178\
        );

    \I__655\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7178\
        );

    \I__654\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7175\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__7178\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__7175\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__651\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7164\
        );

    \I__650\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7161\
        );

    \I__649\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7158\
        );

    \I__648\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7155\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__7164\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__7161\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__7158\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__7155\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__7146\,
            I => \uu0.un4_l_count_13_cascade_\
        );

    \I__642\ : CascadeMux
    port map (
            O => \N__7143\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__641\ : IoInMux
    port map (
            O => \N__7140\,
            I => \N__7137\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__7137\,
            I => \uu0.un11_l_count_i\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__7134\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__638\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7128\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__7128\,
            I => \uu0.un4_l_count_16\
        );

    \I__636\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7118\
        );

    \I__635\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7118\
        );

    \I__634\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7115\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__7118\,
            I => \N__7112\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__7115\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__7112\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__7107\,
            I => \uu0.un88_ci_3_cascade_\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__7104\,
            I => \N__7101\
        );

    \I__628\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7098\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__7098\,
            I => \uu0.un99_ci_0\
        );

    \I__626\ : CascadeMux
    port map (
            O => \N__7095\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__625\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7089\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__7089\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__623\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7083\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__7083\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__621\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7077\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__7077\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__619\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7071\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__7071\,
            I => vbuf_tx_data_4
        );

    \I__617\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7065\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__7065\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__615\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7059\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__7059\,
            I => \N__7056\
        );

    \I__613\ : Span4Mux_v
    port map (
            O => \N__7056\,
            I => \N__7053\
        );

    \I__612\ : Odrv4
    port map (
            O => \N__7053\,
            I => \uu2.r_data_wire_4\
        );

    \I__611\ : InMux
    port map (
            O => \N__7050\,
            I => \N__7047\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__7047\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7041\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__7041\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__607\ : IoInMux
    port map (
            O => \N__7038\,
            I => \N__7035\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__7035\,
            I => \N__7032\
        );

    \I__605\ : IoSpan4Mux
    port map (
            O => \N__7032\,
            I => \N__7029\
        );

    \I__604\ : Span4Mux_s0_h
    port map (
            O => \N__7029\,
            I => \N__7026\
        );

    \I__603\ : Odrv4
    port map (
            O => \N__7026\,
            I => o_serial_data_c
        );

    \I__602\ : IoInMux
    port map (
            O => \N__7023\,
            I => \N__7020\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__7020\,
            I => \N__7017\
        );

    \I__600\ : IoSpan4Mux
    port map (
            O => \N__7017\,
            I => \N__7014\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__7014\,
            I => clk_in_c
        );

    \INVuu2.bitmap_58C\ : INV
    port map (
            O => \INVuu2.bitmap_58C_net\,
            I => \N__18484\
        );

    \INVuu2.w_addr_displaying_7_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_7_rep1C_net\,
            I => \N__18492\
        );

    \INVuu2.w_addr_displaying_ness_6C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_ness_6C_net\,
            I => \N__18499\
        );

    \INVuu2.bitmap_168C\ : INV
    port map (
            O => \INVuu2.bitmap_168C_net\,
            I => \N__18504\
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__18507\
        );

    \INVuu2.bitmap_180C\ : INV
    port map (
            O => \INVuu2.bitmap_180C_net\,
            I => \N__18460\
        );

    \INVuu2.bitmap_34C\ : INV
    port map (
            O => \INVuu2.bitmap_34C_net\,
            I => \N__18467\
        );

    \INVuu2.w_addr_displaying_4_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4_rep1C_net\,
            I => \N__18483\
        );

    \INVuu2.bitmap_75C\ : INV
    port map (
            O => \INVuu2.bitmap_75C_net\,
            I => \N__18498\
        );

    \INVuu2.bitmap_162C\ : INV
    port map (
            O => \INVuu2.bitmap_162C_net\,
            I => \N__18503\
        );

    \INVuu2.w_addr_displaying_3_rep1_nesrC\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            I => \N__18459\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__18466\
        );

    \INVuu2.w_addr_displaying_1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_1C_net\,
            I => \N__18475\
        );

    \INVuu2.bitmap_90C\ : INV
    port map (
            O => \INVuu2.bitmap_90C_net\,
            I => \N__18497\
        );

    \INVuu2.w_addr_displaying_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_3C_net\,
            I => \N__18448\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__18477\
        );

    \INVuu2.w_addr_displaying_0C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_0C_net\,
            I => \N__18474\
        );

    \INVuu2.w_addr_user_nesr_0C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_0C_net\,
            I => \N__18482\
        );

    \INVuu2.w_addr_user_1C\ : INV
    port map (
            O => \INVuu2.w_addr_user_1C_net\,
            I => \N__18473\
        );

    \INVuu2.w_addr_user_8C\ : INV
    port map (
            O => \INVuu2.w_addr_user_8C_net\,
            I => \N__18489\
        );

    \INVuu2.bitmap_111C\ : INV
    port map (
            O => \INVuu2.bitmap_111C_net\,
            I => \N__18472\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__18501\
        );

    \INVuu2.r_data_reg_4C\ : INV
    port map (
            O => \INVuu2.r_data_reg_4C_net\,
            I => \N__18505\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_9_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_10_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_12_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10533\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7140\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10362\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7062\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_4C_net\,
            ce => \N__7461\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8883\,
            in1 => \N__7092\,
            in2 => \_gnd_net_\,
            in3 => \N__7434\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.shifter_0_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7050\,
            in2 => \_gnd_net_\,
            in3 => \N__8881\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.uart_tx_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7044\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.shifter_2_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7086\,
            in1 => \N__8884\,
            in2 => \_gnd_net_\,
            in3 => \N__7419\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.shifter_3_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8885\,
            in1 => \N__7080\,
            in2 => \_gnd_net_\,
            in3 => \N__7407\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.shifter_4_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7068\,
            in1 => \N__8886\,
            in2 => \_gnd_net_\,
            in3 => \N__7395\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \buart.Z_tx.shifter_5_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8887\,
            in1 => \N__7527\,
            in2 => \_gnd_net_\,
            in3 => \N__7074\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18500\,
            ce => \N__7484\,
            sr => \N__18700\
        );

    \uu0.l_count_13_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7895\,
            in1 => \N__9721\,
            in2 => \N__7767\,
            in3 => \N__7824\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18493\,
            ce => \N__8195\,
            sr => \N__18698\
        );

    \uu0.l_count_7_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9722\,
            in1 => \N__7356\,
            in2 => \N__7104\,
            in3 => \N__7123\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18493\,
            ce => \N__8195\,
            sr => \N__18698\
        );

    \uu0.l_count_12_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9720\,
            in1 => \N__7896\,
            in2 => \N__7797\,
            in3 => \N__7812\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18493\,
            ce => \N__8195\,
            sr => \N__18698\
        );

    \uu0.l_count_16_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7897\,
            in1 => \N__9719\,
            in2 => \N__7845\,
            in3 => \N__8067\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18487\,
            ce => \N__8193\,
            sr => \N__18697\
        );

    \uu0.l_count_8_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7898\,
            in2 => \_gnd_net_\,
            in3 => \N__8754\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18487\,
            ce => \N__8193\,
            sr => \N__18697\
        );

    \uu0.l_count_5_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__7280\,
            in1 => \N__7355\,
            in2 => \_gnd_net_\,
            in3 => \N__7170\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18487\,
            ce => \N__8193\,
            sr => \N__18697\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7168\,
            in2 => \_gnd_net_\,
            in3 => \N__7279\,
            lcout => \uu0.un88_ci_3\,
            ltout => \uu0.un88_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7107\,
            in3 => \N__7305\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7988\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7977\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_10_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__8750\,
            in1 => \N__7894\,
            in2 => \N__8786\,
            in3 => \N__8710\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18479\,
            ce => \N__8192\,
            sr => \N__18699\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__7788\,
            in2 => \_gnd_net_\,
            in3 => \N__8042\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7890\,
            in1 => \N__9704\,
            in2 => \N__7095\,
            in3 => \N__7187\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18479\,
            ce => \N__8192\,
            sr => \N__18699\
        );

    \uu0.l_count_14_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__7206\,
            in1 => \N__8043\,
            in2 => \N__7899\,
            in3 => \N__7789\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18479\,
            ce => \N__8192\,
            sr => \N__18699\
        );

    \uu0.l_count_4_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__7354\,
            in1 => \N__9705\,
            in2 => \_gnd_net_\,
            in3 => \N__7169\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18479\,
            ce => \N__8192\,
            sr => \N__18699\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8709\,
            in1 => \N__8779\,
            in2 => \N__7922\,
            in3 => \N__8749\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8041\,
            in1 => \N__7186\,
            in2 => \N__7209\,
            in3 => \N__7204\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIGTCU_15_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8778\,
            in1 => \N__7203\,
            in2 => \N__7188\,
            in3 => \N__7167\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_15_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7239\,
            in1 => \N__7131\,
            in2 => \N__7146\,
            in3 => \N__8019\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_RNILLLG7_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9996\,
            in2 => \N__7143\,
            in3 => \N__10007\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9663\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.sec_clkDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18471\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8708\,
            in1 => \N__7124\,
            in2 => \N__8229\,
            in3 => \N__7939\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIOIDD2_18_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7915\,
            in1 => \N__8207\,
            in2 => \N__7134\,
            in3 => \N__7299\,
            lcout => \uu0.un4_l_count_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7125\,
            in1 => \N__7344\,
            in2 => \N__7326\,
            in3 => \N__7300\,
            lcout => \uu0.un110_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8097\,
            in1 => \N__7262\,
            in2 => \_gnd_net_\,
            in3 => \N__8133\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18462\,
            ce => \N__8194\,
            sr => \N__18701\
        );

    \uu0.l_count_1_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7261\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8096\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18462\,
            ce => \N__8194\,
            sr => \N__18701\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__7260\,
            in2 => \_gnd_net_\,
            in3 => \N__8132\,
            lcout => \uu0.un55_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__9699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8095\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18462\,
            ce => \N__8194\,
            sr => \N__18701\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8131\,
            in1 => \N__7940\,
            in2 => \N__7263\,
            in3 => \N__8093\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_6_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7325\,
            in1 => \N__9700\,
            in2 => \N__7308\,
            in3 => \N__7304\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18462\,
            ce => \N__8194\,
            sr => \N__18701\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8869\,
            in2 => \_gnd_net_\,
            in3 => \N__8327\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8150\,
            in1 => \N__7281\,
            in2 => \N__8175\,
            in3 => \N__7256\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__7545\,
            in1 => \N__7367\,
            in2 => \N__7226\,
            in3 => \N__7714\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18506\,
            ce => \N__7659\,
            sr => \N__18689\
        );

    \uu2.r_addr_esr_3_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15893\,
            in1 => \N__15768\,
            in2 => \N__7630\,
            in3 => \N__15835\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18506\,
            ce => \N__7659\,
            sr => \N__18689\
        );

    \uu2.r_addr_esr_7_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7715\,
            in1 => \N__7591\,
            in2 => \N__7371\,
            in3 => \N__7571\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18506\,
            ce => \N__7659\,
            sr => \N__18689\
        );

    \uu2.r_data_reg_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7440\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7428\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7401\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7383\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7377\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7457\,
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7741\,
            in2 => \_gnd_net_\,
            in3 => \N__7684\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15889\,
            in1 => \N__15754\,
            in2 => \N__7634\,
            in3 => \N__15834\,
            lcout => \uu2.un404_ci\,
            ltout => \uu2.un404_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__7564\,
            in1 => \N__7742\,
            in2 => \N__7602\,
            in3 => \N__7685\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18494\,
            ce => \N__7655\,
            sr => \N__18688\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7595\,
            in2 => \_gnd_net_\,
            in3 => \N__7563\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI83ID7_8_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__9152\,
            in1 => \N__14682\,
            in2 => \N__12810\,
            in3 => \N__11844\,
            lcout => \uu2.w_addr_displaying_nesr_RNI83ID7Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_6_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7512\,
            in1 => \N__8872\,
            in2 => \_gnd_net_\,
            in3 => \N__7536\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18488\,
            ce => \N__7488\,
            sr => \N__18742\
        );

    \buart.Z_tx.shifter_7_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8873\,
            in1 => \N__7497\,
            in2 => \_gnd_net_\,
            in3 => \N__7521\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18488\,
            ce => \N__7488\,
            sr => \N__18742\
        );

    \buart.Z_tx.shifter_8_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8871\,
            in2 => \_gnd_net_\,
            in3 => \N__7506\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18488\,
            ce => \N__7488\,
            sr => \N__18742\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7956\,
            in1 => \N__7971\,
            in2 => \_gnd_net_\,
            in3 => \N__18741\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIMBBL2_7_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15398\,
            in1 => \N__15197\,
            in2 => \_gnd_net_\,
            in3 => \N__15339\,
            lcout => \uu2.N_15_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIFAQ9_13_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7823\,
            in2 => \_gnd_net_\,
            in3 => \N__7810\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7811\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7793\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7758\,
            in2 => \_gnd_net_\,
            in3 => \N__9659\,
            lcout => \oneSecStrb_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_5_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15788\,
            in1 => \N__7683\,
            in2 => \N__7716\,
            in3 => \N__7737\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \uu2.r_addr_4_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__7682\,
            in1 => \N__7710\,
            in2 => \_gnd_net_\,
            in3 => \N__15787\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__15785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18747\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_0_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15824\,
            in2 => \_gnd_net_\,
            in3 => \N__15786\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \Lab_UT.dictrl.alarmstate_ret_1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9599\,
            in2 => \_gnd_net_\,
            in3 => \N__9578\,
            lcout => \Lab_UT.alarmchar10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \Lab_UT.dictrl.alarmstate_ret_2_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__9579\,
            in1 => \_gnd_net_\,
            in2 => \N__9603\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmchar10_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \uu2.trig_rd_det_0_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10074\,
            in2 => \_gnd_net_\,
            in3 => \N__8670\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \uu2.trig_rd_det_1_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7989\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18480\,
            ce => 'H',
            sr => \N__18687\
        );

    \uu2.bitmap_111_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9652\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__18648\
        );

    \uu2.vram_rd_clk_det_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10069\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__18648\
        );

    \uu2.vram_rd_clk_det_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7970\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__18648\
        );

    \uu0.l_count_3_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__7947\,
            in1 => \N__9703\,
            in2 => \_gnd_net_\,
            in3 => \N__7941\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18463\,
            ce => \N__8196\,
            sr => \N__18702\
        );

    \uu0.l_count_9_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7887\,
            in1 => \N__8756\,
            in2 => \_gnd_net_\,
            in3 => \N__8714\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18463\,
            ce => \N__8196\,
            sr => \N__18702\
        );

    \uu0.l_count_17_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__8228\,
            in1 => \N__7840\,
            in2 => \N__8073\,
            in3 => \N__7889\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18463\,
            ce => \N__8196\,
            sr => \N__18702\
        );

    \uu0.l_count_11_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__8685\,
            in1 => \N__9701\,
            in2 => \N__7923\,
            in3 => \N__7888\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18463\,
            ce => \N__8196\,
            sr => \N__18702\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7886\,
            in1 => \N__8069\,
            in2 => \N__7844\,
            in3 => \N__8227\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000010010"
        )
    port map (
            in0 => \N__8208\,
            in1 => \N__9702\,
            in2 => \N__8211\,
            in3 => \_gnd_net_\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18463\,
            ce => \N__8196\,
            sr => \N__18702\
        );

    \uu0.delay_line_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8173\,
            in1 => \N__8151\,
            in2 => \N__8013\,
            in3 => \N__8112\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18456\,
            ce => 'H',
            sr => \N__18703\
        );

    \uu0.l_precount_3_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8114\,
            in1 => \N__8012\,
            in2 => \N__8157\,
            in3 => \N__8174\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18456\,
            ce => 'H',
            sr => \N__18703\
        );

    \uu0.l_precount_1_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8152\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8010\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18456\,
            ce => 'H',
            sr => \N__18703\
        );

    \uu0.l_precount_2_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8011\,
            in1 => \N__8153\,
            in2 => \_gnd_net_\,
            in3 => \N__8113\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18456\,
            ce => 'H',
            sr => \N__18703\
        );

    \uu0.l_precount_RNI3Q7K1_2_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8755\,
            in1 => \N__8130\,
            in2 => \N__8115\,
            in3 => \N__8092\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIO2782_16_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8005\,
            in1 => \N__8068\,
            in2 => \N__8046\,
            in3 => \N__8040\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_0_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8009\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18456\,
            ce => 'H',
            sr => \N__18703\
        );

    \buart.Z_tx.bitcount_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__8870\,
            in1 => \N__8288\,
            in2 => \_gnd_net_\,
            in3 => \N__8328\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18449\,
            ce => 'H',
            sr => \N__18704\
        );

    \buart.Z_tx.bitcount_1_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110110"
        )
    port map (
            in0 => \N__8325\,
            in1 => \N__8304\,
            in2 => \N__8888\,
            in3 => \N__8287\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18442\,
            ce => 'H',
            sr => \N__18706\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__8303\,
            in1 => \N__8256\,
            in2 => \N__8289\,
            in3 => \N__8324\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110111011110"
        )
    port map (
            in0 => \N__8326\,
            in1 => \N__8889\,
            in2 => \N__8346\,
            in3 => \N__8343\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18442\,
            ce => 'H',
            sr => \N__18706\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8282\,
            in2 => \_gnd_net_\,
            in3 => \N__8342\,
            lcout => OPEN,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__8254\,
            in1 => \N__8301\,
            in2 => \N__8331\,
            in3 => \N__9024\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100010000"
        )
    port map (
            in0 => \N__8302\,
            in1 => \N__8283\,
            in2 => \N__8262\,
            in3 => \N__8255\,
            lcout => OPEN,
            ltout => \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__8874\,
            in1 => \_gnd_net_\,
            in2 => \N__8259\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18442\,
            ce => 'H',
            sr => \N__18706\
        );

    \Lab_UT.alarmchar_5_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8244\,
            lcout => \Lab_UT.alarmcharZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18502\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNO_0_8_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001100110011"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__8368\,
            in2 => \N__10255\,
            in3 => \N__9376\,
            lcout => \uu2.N_61_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14529\,
            in1 => \N__12372\,
            in2 => \N__9329\,
            in3 => \N__14396\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14527\,
            in1 => \N__15198\,
            in2 => \N__9378\,
            in3 => \N__14395\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__14394\,
            in1 => \N__14528\,
            in2 => \N__8370\,
            in3 => \N__14668\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIK9E4_2_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__12148\,
            in1 => \N__10306\,
            in2 => \_gnd_net_\,
            in3 => \N__10147\,
            lcout => \uu2.N_102\,
            ltout => \uu2.N_102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIQ6EA_5_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__9233\,
            in1 => \N__8513\,
            in2 => \N__8382\,
            in3 => \N__9324\,
            lcout => \uu2.N_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_8_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__8367\,
            in1 => \N__9285\,
            in2 => \N__8379\,
            in3 => \N__8550\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_8C_net\,
            ce => 'H',
            sr => \N__18652\
        );

    \uu2.w_addr_user_RNO_0_5_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__9346\,
            in1 => \N__9234\,
            in2 => \_gnd_net_\,
            in3 => \N__9325\,
            lcout => \uu2.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI86V6_2_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8512\,
            in1 => \N__9372\,
            in2 => \N__8369\,
            in3 => \N__10146\,
            lcout => \uu2.w_addr_user_3_i_a2_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIR7FF7_6_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10357\,
            in2 => \_gnd_net_\,
            in3 => \N__8544\,
            lcout => \uu2.un28_w_addr_user_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_6_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8487\,
            lcout => \Lab_UT.alarmcharZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18481\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__14375\,
            in1 => \N__14504\,
            in2 => \N__8517\,
            in3 => \N__15578\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI2UTD_1_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8469\,
            in1 => \N__12142\,
            in2 => \N__10305\,
            in3 => \N__8418\,
            lcout => \uu2.N_155\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__13944\,
            in1 => \N__11085\,
            in2 => \N__8448\,
            in3 => \N__10950\,
            lcout => OPEN,
            ltout => \uu2.mem0.g1_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__10485\,
            in1 => \N__8454\,
            in2 => \N__8463\,
            in3 => \N__9432\,
            lcout => \uu2.mem0.N_63_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__11073\,
            in1 => \N__13959\,
            in2 => \N__8447\,
            in3 => \N__9528\,
            lcout => \uu2.mem0.G_17_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_RNIGIDK3_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14374\,
            lcout => \N_72_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14462\,
            in1 => \N__12474\,
            in2 => \N__9240\,
            in3 => \N__14353\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI0FF3_4_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9236\,
            in2 => \_gnd_net_\,
            in3 => \N__9308\,
            lcout => \uu2.w_addr_user_3_i_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNINEKD7_6_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__9404\,
            in1 => \N__9259\,
            in2 => \N__10260\,
            in3 => \N__14461\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => \uu2.un28_w_addr_user_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_1_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001110001001100"
        )
    port map (
            in0 => \N__9260\,
            in1 => \N__10301\,
            in2 => \N__8553\,
            in3 => \N__12149\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__18649\
        );

    \uu2.w_addr_user_3_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000110101010"
        )
    port map (
            in0 => \N__9320\,
            in1 => \N__9261\,
            in2 => \N__9354\,
            in3 => \N__8545\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__18649\
        );

    \uu2.w_addr_user_5_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100000010"
        )
    port map (
            in0 => \N__8546\,
            in1 => \N__8526\,
            in2 => \N__9279\,
            in3 => \N__8511\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__18649\
        );

    \uu2.un28_w_addr_user_i_0_a2_0_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9524\,
            in2 => \_gnd_net_\,
            in3 => \N__9482\,
            lcout => OPEN,
            ltout => \uu2.un28_w_addr_user_i_0_a2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_o4_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__9534\,
            in1 => \N__9502\,
            in2 => \N__8490\,
            in3 => \N__14328\,
            lcout => \uu2.N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000100010"
        )
    port map (
            in0 => \N__10659\,
            in1 => \N__16723\,
            in2 => \N__8637\,
            in3 => \N__16833\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10809\,
            in2 => \_gnd_net_\,
            in3 => \N__10776\,
            lcout => \Lab_UT.alarmchar_2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_RNO_0_4_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8624\,
            in2 => \_gnd_net_\,
            in3 => \N__8587\,
            lcout => OPEN,
            ltout => \resetGen.reset_count_2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101010"
        )
    port map (
            in0 => \N__10387\,
            in1 => \N__8598\,
            in2 => \N__8649\,
            in3 => \N__11271\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_4_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8646\,
            lcout => \Lab_UT.alarmcharZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_3_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__9569\,
            in2 => \_gnd_net_\,
            in3 => \N__10358\,
            lcout => \Lab_UT.dictrl.un1_next_alarmstate21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18464\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__11265\,
            in1 => \N__10391\,
            in2 => \N__8571\,
            in3 => \N__8613\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8612\,
            in1 => \N__8566\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__11267\,
            in1 => \N__10390\,
            in2 => \N__8628\,
            in3 => \N__8625\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8611\,
            in2 => \_gnd_net_\,
            in3 => \N__8565\,
            lcout => \resetGen.un241_ci\,
            ltout => \resetGen.un241_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010100"
        )
    port map (
            in0 => \N__11266\,
            in1 => \N__8589\,
            in2 => \N__8592\,
            in3 => \N__10389\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__10388\,
            in1 => \N__8567\,
            in2 => \_gnd_net_\,
            in3 => \N__11264\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__10073\,
            in1 => \N__8669\,
            in2 => \N__8868\,
            in3 => \N__18748\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8787\,
            in1 => \N__8760\,
            in2 => \_gnd_net_\,
            in3 => \N__8718\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_1_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8920\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8947\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18450\,
            ce => 'H',
            sr => \N__18705\
        );

    \uu2.l_count_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8919\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18450\,
            ce => 'H',
            sr => \N__18705\
        );

    \uu2.l_count_7_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9780\,
            in1 => \N__10694\,
            in2 => \N__8979\,
            in3 => \N__9749\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18450\,
            ce => 'H',
            sr => \N__18705\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9748\,
            in1 => \N__8974\,
            in2 => \N__10695\,
            in3 => \N__9779\,
            lcout => \uu2.un350_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9746\,
            in1 => \N__10715\,
            in2 => \N__8998\,
            in3 => \N__8912\,
            lcout => OPEN,
            ltout => \uu2.un1_l_count_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9965\,
            in1 => \N__8945\,
            in2 => \N__8673\,
            in3 => \N__8958\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_9_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9747\,
            in1 => \N__10716\,
            in2 => \N__8999\,
            in3 => \N__8913\,
            lcout => OPEN,
            ltout => \uu2.un1_l_count_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9966\,
            in1 => \N__8946\,
            in2 => \N__8652\,
            in3 => \N__8957\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10717\,
            in2 => \N__9003\,
            in3 => \N__9778\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18443\,
            ce => 'H',
            sr => \N__18707\
        );

    \uu2.l_count_9_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__9908\,
            in1 => \N__9923\,
            in2 => \N__9000\,
            in3 => \N__10041\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18443\,
            ce => 'H',
            sr => \N__18707\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9065\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8949\,
            in2 => \_gnd_net_\,
            in3 => \N__8922\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIFGGK1_3_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10738\,
            in1 => \N__8978\,
            in2 => \N__9909\,
            in3 => \N__10024\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9066\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9041\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18436\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10025\,
            in1 => \N__8948\,
            in2 => \N__9969\,
            in3 => \N__8921\,
            lcout => \uu2.un306_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9064\,
            in2 => \N__9042\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_13_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9087\,
            in3 => \N__8892\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__18431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9022\,
            in1 => \N__9075\,
            in2 => \_gnd_net_\,
            in3 => \N__9138\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__18431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9114\,
            in3 => \N__9135\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__18431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__9023\,
            in1 => \_gnd_net_\,
            in2 => \N__9126\,
            in3 => \N__9132\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__18431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9101\,
            in1 => \N__9021\,
            in2 => \_gnd_net_\,
            in3 => \N__9129\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18431\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9122\,
            in1 => \N__9110\,
            in2 => \N__9102\,
            in3 => \N__9083\,
            lcout => OPEN,
            ltout => \buart.Z_tx.Z_baudgen.ser_clk_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9074\,
            in1 => \N__9063\,
            in2 => \N__9045\,
            in3 => \N__9037\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_1_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9809\,
            in2 => \_gnd_net_\,
            in3 => \N__16685\,
            lcout => \Lab_UT.cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18490\,
            ce => 'H',
            sr => \N__18693\
        );

    \uu2.w_addr_user_nesr_0_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__12147\,
            in1 => \N__10249\,
            in2 => \N__9416\,
            in3 => \N__9280\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_0C_net\,
            ce => \N__9207\,
            sr => \N__18655\
        );

    \uu2.w_addr_user_nesr_2_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__9281\,
            in1 => \N__12146\,
            in2 => \N__10311\,
            in3 => \N__10149\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_0C_net\,
            ce => \N__9207\,
            sr => \N__18655\
        );

    \uu2.w_addr_user_nesr_6_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__10250\,
            in2 => \N__9417\,
            in3 => \N__9283\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_0C_net\,
            ce => \N__9207\,
            sr => \N__18655\
        );

    \uu2.w_addr_user_nesr_7_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__9284\,
            in1 => \N__9393\,
            in2 => \N__10256\,
            in3 => \N__9377\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_0C_net\,
            ce => \N__9207\,
            sr => \N__18655\
        );

    \uu2.w_addr_user_nesr_4_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011010"
        )
    port map (
            in0 => \N__9235\,
            in1 => \N__9347\,
            in2 => \N__9330\,
            in3 => \N__9282\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_0C_net\,
            ce => \N__9207\,
            sr => \N__18655\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9180\,
            in1 => \N__9507\,
            in2 => \_gnd_net_\,
            in3 => \N__11835\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIARVM2_0_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__15639\,
            in1 => \N__12261\,
            in2 => \_gnd_net_\,
            in3 => \N__15717\,
            lcout => OPEN,
            ltout => \uu2.N_41_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIBTS94_8_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14684\,
            in1 => \N__12075\,
            in2 => \N__9183\,
            in3 => \N__15191\,
            lcout => \uu2.N_132_mux\,
            ltout => \uu2.N_132_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__11836\,
            in1 => \_gnd_net_\,
            in2 => \N__9174\,
            in3 => \N__9483\,
            lcout => \uu2.mem0.N_94_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIREPN6_8_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110100000"
        )
    port map (
            in0 => \N__14685\,
            in1 => \_gnd_net_\,
            in2 => \N__9159\,
            in3 => \N__11834\,
            lcout => \uu2.un21_w_addr_displaying_i\,
            ltout => \uu2.un21_w_addr_displaying_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__15640\,
            in1 => \_gnd_net_\,
            in2 => \N__9459\,
            in3 => \_gnd_net_\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__18653\
        );

    \uu2.w_addr_displaying_fast_1_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__15430\,
            in1 => \N__15641\,
            in2 => \_gnd_net_\,
            in3 => \N__10431\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__18653\
        );

    \uu2.w_addr_displaying_0_rep1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11943\,
            in2 => \_gnd_net_\,
            in3 => \N__15429\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__18653\
        );

    \Lab_UT.bcd2segment1.m68_bm_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100110111"
        )
    port map (
            in0 => \N__10458\,
            in1 => \N__16825\,
            in2 => \N__16722\,
            in3 => \N__19443\,
            lcout => \Lab_UT.bcd2segment1.m68_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011000100"
        )
    port map (
            in0 => \N__16826\,
            in1 => \N__10662\,
            in2 => \N__9456\,
            in3 => \N__16706\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_30_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111110011"
        )
    port map (
            in0 => \N__11176\,
            in1 => \N__12472\,
            in2 => \N__12771\,
            in3 => \N__12324\,
            lcout => \uu2.mem0.N_13_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIDKOL_1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11178\,
            lcout => \uu2.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_32_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__11177\,
            in1 => \N__15642\,
            in2 => \N__10191\,
            in3 => \N__11976\,
            lcout => OPEN,
            ltout => \uu2.mem0.i14_mux_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_18_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__12558\,
            in1 => \N__9441\,
            in2 => \N__9435\,
            in3 => \N__12618\,
            lcout => \uu2.mem0.N_8_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16705\,
            in1 => \N__16827\,
            in2 => \N__9426\,
            in3 => \N__10658\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__10657\,
            in1 => \N__9627\,
            in2 => \_gnd_net_\,
            in3 => \N__9549\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9810\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__10660\,
            in1 => \N__9540\,
            in2 => \_gnd_net_\,
            in3 => \N__10401\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_a2_4_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14414\,
            in1 => \N__11861\,
            in2 => \N__10109\,
            in3 => \N__11041\,
            lcout => \uu2.un28_w_addr_user_i_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__10661\,
            in1 => \N__10596\,
            in2 => \_gnd_net_\,
            in3 => \N__9618\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18458\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_47_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001001"
        )
    port map (
            in0 => \N__12473\,
            in1 => \N__11164\,
            in2 => \N__12754\,
            in3 => \N__12328\,
            lcout => \uu2.mem0.g0_7_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_data_i_o2_4_0_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__9523\,
            in1 => \N__14413\,
            in2 => \N__9506\,
            in3 => \N__9481\,
            lcout => OPEN,
            ltout => \uu2.w_data_i_o2_4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_data_i_o2_0_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__10105\,
            in1 => \N__11860\,
            in2 => \N__9465\,
            in3 => \N__11042\,
            lcout => \N_96\,
            ltout => \N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_data_i_0_tz_0_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9462\,
            in3 => \N__14460\,
            lcout => \uu2.w_data_i_0_tzZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m59_bm_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101011111"
        )
    port map (
            in0 => \N__9612\,
            in1 => \N__18096\,
            in2 => \N__16828\,
            in3 => \N__16695\,
            lcout => \Lab_UT.bcd2segment1.m59_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m52_am_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011111100"
        )
    port map (
            in0 => \N__16811\,
            in1 => \N__10446\,
            in2 => \N__16721\,
            in3 => \N__14166\,
            lcout => \Lab_UT.bcd2segment1.m52_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10584\,
            in2 => \_gnd_net_\,
            in3 => \N__10808\,
            lcout => \Lab_UT.alarmcharZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111110101011"
        )
    port map (
            in0 => \N__10350\,
            in1 => \N__13329\,
            in2 => \N__13314\,
            in3 => \N__13251\,
            lcout => \Lab_UT.dictrl.state_retZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18451\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__9828\,
            in1 => \N__9873\,
            in2 => \N__10854\,
            in3 => \N__10751\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9874\,
            in1 => \N__9827\,
            in2 => \_gnd_net_\,
            in3 => \N__10561\,
            lcout => \Lab_UT.dictrl.next_alarmstateZ0Z_0\,
            ltout => \Lab_UT.dictrl.next_alarmstateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__G_74_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__9829\,
            in1 => \N__9568\,
            in2 => \N__9552\,
            in3 => \N__10349\,
            lcout => \Lab_UT.dictrl.G_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m59_am_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110110000"
        )
    port map (
            in0 => \N__16810\,
            in1 => \N__14255\,
            in2 => \N__16720\,
            in3 => \N__16311\,
            lcout => \Lab_UT.bcd2segment1.m59_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_0_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__10847\,
            in1 => \N__9840\,
            in2 => \N__9888\,
            in3 => \N__10752\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.dictrl.alarmstate_0_0_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9883\,
            in1 => \N__9838\,
            in2 => \_gnd_net_\,
            in3 => \N__10562\,
            lcout => \Lab_UT.dictrl.alarmstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.dictrl.alarmstate_ret_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__10563\,
            in1 => \N__9884\,
            in2 => \_gnd_net_\,
            in3 => \N__9839\,
            lcout => \Lab_UT.dictrl.alarmstate_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.dispString.cnt_3_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__16816\,
            in1 => \N__9797\,
            in2 => \N__16724\,
            in3 => \N__10639\,
            lcout => \Lab_UT.cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.dispString.cnt_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__9795\,
            in1 => \N__16711\,
            in2 => \N__10656\,
            in3 => \N__16817\,
            lcout => \Lab_UT.cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.dispString.cnt_2_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__16710\,
            in1 => \N__10635\,
            in2 => \_gnd_net_\,
            in3 => \N__9796\,
            lcout => \Lab_UT.cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18444\,
            ce => 'H',
            sr => \N__18690\
        );

    \Lab_UT.bcd2segment1.m8_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14102\,
            in1 => \N__14266\,
            in2 => \_gnd_net_\,
            in3 => \N__14177\,
            lcout => \Lab_UT.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_5_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__9777\,
            in1 => \N__10721\,
            in2 => \_gnd_net_\,
            in3 => \N__10740\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu2.l_count_6_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10685\,
            in1 => \N__9753\,
            in2 => \_gnd_net_\,
            in3 => \N__9776\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \Lab_UT.dictrl.state_ret_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13293\,
            in2 => \_gnd_net_\,
            in3 => \N__13272\,
            lcout => \Lab_UT.dictrl.dicRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu0.sec_clk_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9643\,
            in2 => \_gnd_net_\,
            in3 => \N__9726\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu2.vram_rd_clk_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10059\,
            in2 => \_gnd_net_\,
            in3 => \N__10039\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu2.l_count_3_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__9968\,
            in1 => \N__10040\,
            in2 => \N__9984\,
            in3 => \N__10026\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu0.delay_line_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10011\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18437\,
            ce => 'H',
            sr => \N__18691\
        );

    \uu2.l_count_2_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9980\,
            in2 => \_gnd_net_\,
            in3 => \N__9967\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18432\,
            ce => 'H',
            sr => \N__18708\
        );

    \buart.Z_rx.hh_0_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9939\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18432\,
            ce => 'H',
            sr => \N__18708\
        );

    \uu2.l_count_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9907\,
            in2 => \_gnd_net_\,
            in3 => \N__9924\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18432\,
            ce => 'H',
            sr => \N__18708\
        );

    \Lab_UT.dictrl.next_alarmstate_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.next_alarmstate_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18427\,
            ce => \N__9852\,
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13358\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18425\,
            ce => 'H',
            sr => \N__18709\
        );

    \Lab_UT.bcd2segment1.m89_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101110110111"
        )
    port map (
            in0 => \N__19072\,
            in1 => \N__19362\,
            in2 => \N__19180\,
            in3 => \N__19284\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_187_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10179\,
            in3 => \N__14982\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__18659\
        );

    \Lab_UT.bcd2segment1.m92_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111010111111"
        )
    port map (
            in0 => \N__19073\,
            in1 => \N__19363\,
            in2 => \N__19181\,
            in3 => \N__19285\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_221_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10176\,
            in3 => \N__14981\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__18659\
        );

    \uu2.mem0.ram512X8_inst_RNO_78_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001011111"
        )
    port map (
            in0 => \N__15996\,
            in1 => \_gnd_net_\,
            in2 => \N__10164\,
            in3 => \N__10173\,
            lcout => \uu2.mem0.N_107_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_83_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__10172\,
            in1 => \N__10160\,
            in2 => \_gnd_net_\,
            in3 => \N__15995\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_107_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_59_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__11952\,
            in1 => \N__15906\,
            in2 => \N__10152\,
            in3 => \N__10926\,
            lcout => \uu2.mem0.N_74_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__14388\,
            in1 => \N__10148\,
            in2 => \N__14532\,
            in3 => \N__12759\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_23_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12074\,
            in1 => \N__15192\,
            in2 => \N__14670\,
            in3 => \N__15713\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_130_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14526\,
            in1 => \N__10113\,
            in2 => \N__10089\,
            in3 => \N__14389\,
            lcout => \uu2.mem0.N_54_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_33_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000001100"
        )
    port map (
            in0 => \N__11138\,
            in1 => \N__12475\,
            in2 => \N__12770\,
            in3 => \N__12360\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_19_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__11055\,
            in1 => \N__14521\,
            in2 => \N__10263\,
            in3 => \N__14387\,
            lcout => \uu2.mem0.G_13_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__14525\,
            in1 => \N__15329\,
            in2 => \N__10251\,
            in3 => \N__14390\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_50_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12609\,
            in1 => \N__16104\,
            in2 => \N__13919\,
            in3 => \N__11936\,
            lcout => \uu2.mem0.G_13_0_a3_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_55_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__10437\,
            in1 => \N__11939\,
            in2 => \N__10890\,
            in3 => \N__10200\,
            lcout => \uu2.mem0.N_74_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_66_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__11938\,
            in1 => \N__13811\,
            in2 => \N__12477\,
            in3 => \N__16103\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_87_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001001"
        )
    port map (
            in0 => \N__13810\,
            in1 => \N__12608\,
            in2 => \N__16117\,
            in3 => \N__12840\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_7_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_62_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000001111"
        )
    port map (
            in0 => \N__14732\,
            in1 => \N__14277\,
            in2 => \N__10182\,
            in3 => \N__10413\,
            lcout => \uu2.mem0.g0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_91_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__13989\,
            in1 => \N__10430\,
            in2 => \N__11208\,
            in3 => \N__12492\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_85_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100000111"
        )
    port map (
            in0 => \N__15330\,
            in1 => \N__15573\,
            in2 => \N__10440\,
            in3 => \N__10412\,
            lcout => \uu2.mem0.N_57_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_64_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__11937\,
            in1 => \N__12471\,
            in2 => \N__13827\,
            in3 => \N__12341\,
            lcout => \uu2.mem0.g0_i_m2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_77_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__16014\,
            in1 => \N__15994\,
            in2 => \_gnd_net_\,
            in3 => \N__15924\,
            lcout => \uu2.mem0.N_98_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI64LA_1_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000110000001"
        )
    port map (
            in0 => \N__10429\,
            in1 => \N__12839\,
            in2 => \N__11204\,
            in3 => \_gnd_net_\,
            lcout => \uu2.N_1585_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m62_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__16823\,
            in1 => \N__19368\,
            in2 => \_gnd_net_\,
            in3 => \N__12923\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.i6_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m68_am_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001110100"
        )
    port map (
            in0 => \N__16252\,
            in1 => \N__16694\,
            in2 => \N__10404\,
            in3 => \N__16824\,
            lcout => \Lab_UT.bcd2segment1.m68_amZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIV7KP6_8_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10339\,
            in2 => \_gnd_net_\,
            in3 => \N__15428\,
            lcout => \uu2.un21_w_addr_displaying_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_39_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15335\,
            in2 => \_gnd_net_\,
            in3 => \N__15581\,
            lcout => \uu2.mem0.N_126_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10395\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18455\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14352\,
            in1 => \N__10310\,
            in2 => \N__11180\,
            in3 => \N__14487\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__10532\,
            in1 => \N__14486\,
            in2 => \_gnd_net_\,
            in3 => \N__14351\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_36_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__15187\,
            in1 => \N__15332\,
            in2 => \N__14683\,
            in3 => \N__15582\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_20_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__10467\,
            in1 => \N__10473\,
            in2 => \N__10488\,
            in3 => \N__14736\,
            lcout => \uu2.mem0.g1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_35_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__12736\,
            in1 => \N__11168\,
            in2 => \_gnd_net_\,
            in3 => \N__12325\,
            lcout => \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_37_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001001001001"
        )
    port map (
            in0 => \N__12326\,
            in1 => \N__12737\,
            in2 => \N__11179\,
            in3 => \N__12476\,
            lcout => \uu2.mem0.g0_7_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_3_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15678\,
            in1 => \N__11172\,
            in2 => \N__12755\,
            in3 => \N__12327\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_3C_net\,
            ce => \N__14578\,
            sr => \N__18650\
        );

    \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10583\,
            in2 => \_gnd_net_\,
            in3 => \N__10807\,
            lcout => OPEN,
            ltout => \Lab_UT.alarmchar9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_2_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10461\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmcharZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m47_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__19173\,
            in1 => \N__16790\,
            in2 => \_gnd_net_\,
            in3 => \N__13049\,
            lcout => \Lab_UT.bcd2segment1.N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m36_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__16812\,
            in1 => \N__19287\,
            in2 => \_gnd_net_\,
            in3 => \N__12985\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.i5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m42_am_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000011"
        )
    port map (
            in0 => \N__16794\,
            in1 => \N__16719\,
            in2 => \N__10665\,
            in3 => \N__14103\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.m42_amZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10634\,
            in2 => \N__10599\,
            in3 => \N__16626\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18441\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m52_bm_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011100"
        )
    port map (
            in0 => \N__16844\,
            in1 => \N__16718\,
            in2 => \N__16822\,
            in3 => \N__18026\,
            lcout => \Lab_UT.bcd2segment1.m52_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m47_0_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__10590\,
            in1 => \N__13050\,
            in2 => \N__17760\,
            in3 => \N__13628\,
            lcout => \Lab_UT.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m41_0_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12913\,
            in1 => \N__12967\,
            in2 => \_gnd_net_\,
            in3 => \N__16373\,
            lcout => \Lab_UT.bcd2segment1.N_42_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10770\,
            in2 => \_gnd_net_\,
            in3 => \N__10801\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__10582\,
            in1 => \N__10846\,
            in2 => \N__10566\,
            in3 => \N__11330\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10771\,
            in2 => \_gnd_net_\,
            in3 => \N__10803\,
            lcout => \Lab_UT.alarmcharZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18435\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m49_0_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__12912\,
            in1 => \N__12966\,
            in2 => \_gnd_net_\,
            in3 => \N__16374\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m54_0_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13627\,
            in2 => \N__10812\,
            in3 => \N__17709\,
            lcout => \Lab_UT.q_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__10802\,
            in1 => \N__10772\,
            in2 => \_gnd_net_\,
            in3 => \N__11331\,
            lcout => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__11390\,
            in1 => \N__11409\,
            in2 => \_gnd_net_\,
            in3 => \N__16514\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10739\,
            in2 => \_gnd_net_\,
            in3 => \N__10722\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m60_0_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001100110"
        )
    port map (
            in0 => \N__12971\,
            in1 => \N__16378\,
            in2 => \N__11574\,
            in3 => \N__13626\,
            lcout => OPEN,
            ltout => \Lab_UT.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__13194\,
            in1 => \N__13163\,
            in2 => \N__10668\,
            in3 => \N__12972\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11389\,
            in2 => \_gnd_net_\,
            in3 => \N__16513\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18430\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_4_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11667\,
            in1 => \N__11570\,
            in2 => \N__11742\,
            in3 => \N__17752\,
            lcout => \resetGen.escKeyZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI18N1_5_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11495\,
            in2 => \_gnd_net_\,
            in3 => \N__11388\,
            lcout => \buart.Z_rx.ser_clk_2\,
            ltout => \buart.Z_rx.ser_clk_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__11481\,
            in1 => \N__17094\,
            in2 => \N__10860\,
            in3 => \N__16515\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18426\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11361\,
            in1 => \N__11408\,
            in2 => \N__11448\,
            in3 => \N__11466\,
            lcout => \buart.Z_rx.ser_clk_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state16_5_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11731\,
            in1 => \N__11656\,
            in2 => \N__11703\,
            in3 => \N__11528\,
            lcout => \Lab_UT.dictrl.next_state16Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_2_0_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11529\,
            in1 => \N__11733\,
            in2 => \N__11666\,
            in3 => \N__17741\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_alarmstate4_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17703\,
            in1 => \N__10824\,
            in2 => \N__10857\,
            in3 => \N__11561\,
            lcout => \Lab_UT.dictrl.next_alarmstateZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11692\,
            in2 => \_gnd_net_\,
            in3 => \N__11599\,
            lcout => \Lab_UT.dictrl.next_alarmstate4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_sqmuxa_3_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__17702\,
            in1 => \N__11530\,
            in2 => \N__11704\,
            in3 => \N__11562\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__10872\,
            in2 => \N__10818\,
            in3 => \N__17742\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIHE146_2_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__14947\,
            in1 => \N__13427\,
            in2 => \N__10815\,
            in3 => \N__11433\,
            lcout => \Lab_UT.dictrl.next_state_set\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_sqmuxa_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11732\,
            in2 => \_gnd_net_\,
            in3 => \N__11600\,
            lcout => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_sqmuxa_0_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11602\,
            in2 => \_gnd_net_\,
            in3 => \N__17739\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_3_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11665\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18423\,
            ce => \N__17660\,
            sr => \N__18710\
        );

    \buart.Z_rx.shifter_1_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18423\,
            ce => \N__17660\,
            sr => \N__18710\
        );

    \buart.Z_rx.shifter_4_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18423\,
            ce => \N__17660\,
            sr => \N__18710\
        );

    \buart.Z_rx.shifter_5_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11740\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18423\,
            ce => \N__17660\,
            sr => \N__18710\
        );

    \Lab_UT.bcd2segment1.m99_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__19349\,
            in1 => \N__19283\,
            in2 => \N__19179\,
            in3 => \N__19071\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_90_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10863\,
            in3 => \N__14980\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__18663\
        );

    \Lab_UT.bcd2segment1.segmentUQ_1_4_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100010"
        )
    port map (
            in0 => \N__19348\,
            in1 => \N__19282\,
            in2 => \N__19178\,
            in3 => \N__19070\,
            lcout => \Lab_UT.bcd2segment1.segmentUQ_0_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_90_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__10901\,
            in1 => \N__15053\,
            in2 => \_gnd_net_\,
            in3 => \N__10910\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_92_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_84_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011000110111"
        )
    port map (
            in0 => \N__11954\,
            in1 => \N__12220\,
            in2 => \N__10929\,
            in3 => \N__11768\,
            lcout => \uu2.mem0.m73_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_218_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10920\,
            in2 => \_gnd_net_\,
            in3 => \N__14979\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_90C_net\,
            ce => 'H',
            sr => \N__18663\
        );

    \uu2.mem0.ram512X8_inst_RNO_88_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110101111"
        )
    port map (
            in0 => \N__15054\,
            in1 => \_gnd_net_\,
            in2 => \N__10914\,
            in3 => \N__10902\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_92_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_79_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__11769\,
            in1 => \N__12222\,
            in2 => \N__10893\,
            in3 => \N__11955\,
            lcout => \uu2.mem0.m73_ns_1_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m26_0_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14057\,
            in2 => \_gnd_net_\,
            in3 => \N__14243\,
            lcout => \Lab_UT.N_27_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_40_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011010010000"
        )
    port map (
            in0 => \N__15677\,
            in1 => \N__11163\,
            in2 => \N__11972\,
            in3 => \N__10878\,
            lcout => \uu2.mem0.i14_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__16302\,
            in1 => \N__14058\,
            in2 => \N__13113\,
            in3 => \N__14244\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18491\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m106_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011000011"
        )
    port map (
            in0 => \N__14242\,
            in1 => \N__14154\,
            in2 => \N__14083\,
            in3 => \N__16241\,
            lcout => \Lab_UT.bcd2segment1.N_244\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_34_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15328\,
            in2 => \_gnd_net_\,
            in3 => \N__15580\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14386\,
            in1 => \N__14520\,
            in2 => \_gnd_net_\,
            in3 => \N__11049\,
            lcout => \uu2.mem0.N_93_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_60_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12433\,
            in1 => \N__12359\,
            in2 => \N__13920\,
            in3 => \N__13826\,
            lcout => \uu2.mem0.N_67_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_61_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__14519\,
            in1 => \N__14385\,
            in2 => \_gnd_net_\,
            in3 => \N__11019\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_41_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__13932\,
            in1 => \N__11013\,
            in2 => \N__11007\,
            in3 => \N__11004\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_21_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000010000"
        )
    port map (
            in0 => \N__10998\,
            in1 => \N__10992\,
            in2 => \N__10980\,
            in3 => \N__12000\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__10977\,
            in1 => \N__12021\,
            in2 => \N__10971\,
            in3 => \N__14289\,
            lcout => \uu2.mem0.N_66_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_42_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__10956\,
            in1 => \N__15331\,
            in2 => \N__10938\,
            in3 => \N__15577\,
            lcout => \uu2.mem0.g2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_65_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__12331\,
            in1 => \N__13904\,
            in2 => \_gnd_net_\,
            in3 => \N__13816\,
            lcout => \uu2.mem0.bitmap_pmux_u_i_4_0_N_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_RNINBDH1_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11130\,
            in1 => \N__12426\,
            in2 => \N__13917\,
            in3 => \N__12330\,
            lcout => \uu2.N_67_1_0\,
            ltout => \uu2.N_67_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_25_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__15651\,
            in1 => \_gnd_net_\,
            in2 => \N__11076\,
            in3 => \N__11064\,
            lcout => \uu2.mem0.N_55_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_48_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__13900\,
            in1 => \N__12425\,
            in2 => \_gnd_net_\,
            in3 => \N__12329\,
            lcout => \uu2.mem0.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__15652\,
            in1 => \N__11131\,
            in2 => \_gnd_net_\,
            in3 => \N__15451\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__18657\
        );

    \uu2.w_addr_displaying_1_rep1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__15452\,
            in1 => \_gnd_net_\,
            in2 => \N__13828\,
            in3 => \N__15653\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__18657\
        );

    \uu2.w_addr_displaying_1_rep1_RNIKGI51_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12424\,
            in1 => \N__16102\,
            in2 => \N__13918\,
            in3 => \N__13815\,
            lcout => \uu2.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m118_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111001010"
        )
    port map (
            in0 => \N__14245\,
            in1 => \N__14161\,
            in2 => \N__14098\,
            in3 => \N__16242\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_250_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11058\,
            in3 => \N__14935\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__18656\
        );

    \Lab_UT.bcd2segment1.m97_0_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100110000010"
        )
    port map (
            in0 => \N__14246\,
            in1 => \N__14162\,
            in2 => \N__14099\,
            in3 => \N__16243\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11244\,
            in3 => \N__14936\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__18656\
        );

    \uu2.mem0.ram512X8_inst_RNO_74_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__11237\,
            in1 => \_gnd_net_\,
            in2 => \N__11226\,
            in3 => \N__14784\,
            lcout => \uu2.mem0.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIJVK41_40_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111010011"
        )
    port map (
            in0 => \N__11241\,
            in1 => \N__13217\,
            in2 => \N__12221\,
            in3 => \N__11222\,
            lcout => OPEN,
            ltout => \uu2.m95_i_m2_i_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI19S42_34_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110101"
        )
    port map (
            in0 => \N__12525\,
            in1 => \N__12549\,
            in2 => \N__11214\,
            in3 => \N__12213\,
            lcout => \uu2.N_16\,
            ltout => \uu2.N_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_57_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000001"
        )
    port map (
            in0 => \N__15183\,
            in1 => \N__12432\,
            in2 => \N__11211\,
            in3 => \N__11993\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_nesr_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15679\,
            in1 => \N__12731\,
            in2 => \N__11181\,
            in3 => \N__12214\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            ce => \N__14579\,
            sr => \N__18651\
        );

    \uu2.w_addr_displaying_fast_nesr_3_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11151\,
            in1 => \N__15681\,
            in2 => \N__12753\,
            in3 => \N__11203\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            ce => \N__14579\,
            sr => \N__18651\
        );

    \uu2.w_addr_displaying_3_rep2_nesr_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15680\,
            in1 => \N__11152\,
            in2 => \N__16116\,
            in3 => \N__12732\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            ce => \N__14579\,
            sr => \N__18651\
        );

    \uu2.w_addr_displaying_8_rep1_nesr_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15333\,
            in1 => \N__15189\,
            in2 => \N__15399\,
            in3 => \N__14786\,
            lcout => \uu2.w_addr_displaying_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            ce => \N__14579\,
            sr => \N__18651\
        );

    \uu2.w_addr_displaying_fast_nesr_8_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15188\,
            in1 => \N__15334\,
            in2 => \N__13221\,
            in3 => \N__15396\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3_rep1_nesrC_net\,
            ce => \N__14579\,
            sr => \N__18651\
        );

    \CONSTANT_ONE_LUT4_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_0_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__18091\,
            in1 => \N__18025\,
            in2 => \N__18178\,
            in3 => \N__19436\,
            lcout => \Lab_UT.bcd2segment2.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_70_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14793\,
            in1 => \N__12651\,
            in2 => \_gnd_net_\,
            in3 => \N__13233\,
            lcout => \uu2.mem0.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__13102\,
            in1 => \N__11297\,
            in2 => \N__16295\,
            in3 => \N__16254\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__16167\,
            in1 => \N__14160\,
            in2 => \N__11301\,
            in3 => \N__13098\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__16288\,
            in1 => \_gnd_net_\,
            in2 => \N__13106\,
            in3 => \N__14241\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18452\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.un1_num_1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19435\,
            in1 => \N__18090\,
            in2 => \N__18027\,
            in3 => \N__18166\,
            lcout => \Lab_UT.zero\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_71_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14785\,
            in1 => \N__12524\,
            in2 => \_gnd_net_\,
            in3 => \N__12548\,
            lcout => \uu2.mem0.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11757\,
            in1 => \N__11283\,
            in2 => \_gnd_net_\,
            in3 => \N__17058\,
            lcout => \resetGen.escKeyZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_67_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000010001"
        )
    port map (
            in0 => \N__13913\,
            in1 => \N__16108\,
            in2 => \_gnd_net_\,
            in3 => \N__13829\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNIASM81_2_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12959\,
            in1 => \N__16360\,
            in2 => \N__12901\,
            in3 => \N__14216\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.did_alarmMatch_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIUG9D3_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14076\,
            in1 => \N__11322\,
            in2 => \N__11340\,
            in3 => \N__11337\,
            lcout => \Lab_UT.alarmMatch\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNISKK51_3_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__13051\,
            in1 => \N__14136\,
            in2 => \_gnd_net_\,
            in3 => \N__16214\,
            lcout => \Lab_UT.didp.countrce3.did_alarmMatch_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__11316\,
            in1 => \N__13162\,
            in2 => \N__13190\,
            in3 => \N__13052\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m65_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__13629\,
            in1 => \N__16361\,
            in2 => \_gnd_net_\,
            in3 => \N__11532\,
            lcout => OPEN,
            ltout => \Lab_UT.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__16362\,
            in1 => \N__13182\,
            in2 => \N__11310\,
            in3 => \N__13158\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__12883\,
            in1 => \N__13183\,
            in2 => \N__13164\,
            in3 => \N__11307\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18445\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17877\,
            in2 => \_gnd_net_\,
            in3 => \N__18746\,
            lcout => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI72HD1_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11421\,
            in2 => \_gnd_net_\,
            in3 => \N__17948\,
            lcout => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1\,
            ltout => \Lab_UT.dictrl.next_state_RNI72HD1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__17949\,
            in1 => \N__17547\,
            in2 => \N__11424\,
            in3 => \N__17804\,
            lcout => \Lab_UT.dictrl.next_state_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18438\,
            ce => \N__17494\,
            sr => \N__13647\
        );

    \Lab_UT.dictrl.state_0_RNITK4F_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__16907\,
            in1 => \N__13776\,
            in2 => \_gnd_net_\,
            in3 => \N__13507\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_RNIS90D1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__18908\,
            in1 => \N__16908\,
            in2 => \N__11415\,
            in3 => \N__18953\,
            lcout => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1\,
            ltout => \Lab_UT.dictrl.state_ret_3_RNIS90DZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIR0FR1_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11412\,
            in3 => \N__16551\,
            lcout => \Lab_UT.dictrl.next_state_RNIR0FR1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18983\,
            in1 => \N__18952\,
            in2 => \_gnd_net_\,
            in3 => \N__18877\,
            lcout => \Lab_UT.Run\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11407\,
            in2 => \N__11391\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11465\,
            in2 => \_gnd_net_\,
            in3 => \N__11364\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16487\,
            in1 => \N__11357\,
            in2 => \_gnd_net_\,
            in3 => \N__11346\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__18433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11447\,
            in2 => \_gnd_net_\,
            in3 => \N__11343\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11496\,
            in2 => \_gnd_net_\,
            in3 => \N__11484\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__16485\,
            in1 => \N__17087\,
            in2 => \N__11475\,
            in3 => \N__17121\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIPU6T9_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__17945\,
            in1 => \N__17911\,
            in2 => \N__17870\,
            in3 => \N__17796\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__16486\,
            in1 => \N__17122\,
            in2 => \N__17100\,
            in3 => \N__11454\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18433\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_7_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18428\,
            ce => \N__17653\,
            sr => \N__18711\
        );

    \buart.Z_rx.shifter_6_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11702\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18428\,
            ce => \N__17653\,
            sr => \N__18711\
        );

    \Lab_UT.dictrl.state_0_RNILGF17_3_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__13640\,
            in1 => \N__11748\,
            in2 => \N__14934\,
            in3 => \N__11621\,
            lcout => \Lab_UT.dictrl.next_state_set_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__13586\,
            in1 => \N__13770\,
            in2 => \_gnd_net_\,
            in3 => \N__13565\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxa_1\,
            ltout => \Lab_UT.dictrl.next_state_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIJ9317_2_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__11622\,
            in1 => \N__14886\,
            in2 => \N__11427\,
            in3 => \N__17465\,
            lcout => \Lab_UT.dictrl.next_state_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_5_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__17704\,
            in1 => \N__11531\,
            in2 => \N__11706\,
            in3 => \N__11610\,
            lcout => \resetGen.escKeyZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNICJTA2_3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__13548\,
            in1 => \N__13585\,
            in2 => \_gnd_net_\,
            in3 => \N__13564\,
            lcout => \Lab_UT.dictrl.next_state_set_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_sqmuxa_4_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__11741\,
            in1 => \N__11524\,
            in2 => \N__11705\,
            in3 => \N__11560\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_sqmuxa_5_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11661\,
            in1 => \N__11631\,
            in2 => \N__11625\,
            in3 => \N__17686\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNI0MRT_1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__18969\,
            in1 => \N__16905\,
            in2 => \_gnd_net_\,
            in3 => \N__13516\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_state_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIS90D1_2_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__13771\,
            in1 => \N__16906\,
            in2 => \N__11613\,
            in3 => \N__18904\,
            lcout => \Lab_UT.dictrl.state_0_RNIS90D1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state16_4_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11601\,
            in1 => \N__11559\,
            in2 => \N__17701\,
            in3 => \N__17740\,
            lcout => \Lab_UT.dictrl.next_state16Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11569\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18424\,
            ce => \N__17661\,
            sr => \N__18712\
        );

    \Lab_UT.bcd2segment1.m84_0_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101100110"
        )
    port map (
            in0 => \N__13063\,
            in1 => \N__12920\,
            in2 => \N__16408\,
            in3 => \N__13000\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_127_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11790\,
            in3 => \N__14989\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_162C_net\,
            ce => 'H',
            sr => \N__18666\
        );

    \Lab_UT.bcd2segment1.m87_0_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001100111"
        )
    port map (
            in0 => \N__13064\,
            in1 => \N__12921\,
            in2 => \N__16409\,
            in3 => \N__13001\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_235_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_66_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11787\,
            in3 => \N__14991\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_162C_net\,
            ce => 'H',
            sr => \N__18666\
        );

    \Lab_UT.bcd2segment1.m90_0_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__13065\,
            in1 => \N__12922\,
            in2 => \N__16410\,
            in3 => \N__13002\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_194_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11784\,
            in3 => \N__14990\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_162C_net\,
            ce => 'H',
            sr => \N__18666\
        );

    \uu2.bitmap_RNIIGUI_66_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__11781\,
            in1 => \N__15044\,
            in2 => \_gnd_net_\,
            in3 => \N__11775\,
            lcout => \uu2.N_101_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m93_0_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101101011"
        )
    port map (
            in0 => \N__12999\,
            in1 => \N__16398\,
            in2 => \N__12924\,
            in3 => \N__13062\,
            lcout => \Lab_UT.bcd2segment1.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m101_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__14259\,
            in1 => \N__14180\,
            in2 => \N__14084\,
            in3 => \N__16255\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11760\,
            in3 => \N__14985\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_75C_net\,
            ce => 'H',
            sr => \N__18664\
        );

    \Lab_UT.bcd2segment3.segment_0_2_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__14260\,
            in1 => \N__14181\,
            in2 => \N__14085\,
            in3 => \N__16256\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segment_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_203_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11982\,
            in3 => \N__14983\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_75C_net\,
            ce => 'H',
            sr => \N__18664\
        );

    \uu2.bitmap_RNIC6T81_212_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000011"
        )
    port map (
            in0 => \N__11874\,
            in1 => \N__15992\,
            in2 => \N__12663\,
            in3 => \N__13701\,
            lcout => OPEN,
            ltout => \uu2.N_1580_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIL4F73_3_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12368\,
            in2 => \N__11979\,
            in3 => \N__11880\,
            lcout => \uu2.N_77_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIPIHG1_75_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100100010"
        )
    port map (
            in0 => \N__11953\,
            in1 => \N__11895\,
            in2 => \N__11889\,
            in3 => \N__13995\,
            lcout => \uu2.N_1581_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_212_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18195\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14984\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_75C_net\,
            ce => 'H',
            sr => \N__18664\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15157\,
            in1 => \N__12064\,
            in2 => \N__14669\,
            in3 => \N__11796\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_134_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11868\,
            in2 => \N__11847\,
            in3 => \N__11843\,
            lcout => \uu2.mem0.N_60_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_28_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__15675\,
            in1 => \N__12257\,
            in2 => \_gnd_net_\,
            in3 => \N__15711\,
            lcout => \uu2.mem0.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIF00Q_5_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15550\,
            lcout => \uu2.N_126\,
            ltout => \uu2.N_126_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_46_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110110"
        )
    port map (
            in0 => \N__15156\,
            in1 => \N__14652\,
            in2 => \N__12153\,
            in3 => \N__15712\,
            lcout => \uu2.mem0.bitmap_pmux_u_i_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__14531\,
            in1 => \N__15676\,
            in2 => \N__14397\,
            in3 => \N__12150\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_44_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12099\,
            in1 => \N__12087\,
            in2 => \_gnd_net_\,
            in3 => \N__12063\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_24_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__14697\,
            in1 => \N__12045\,
            in2 => \N__12030\,
            in3 => \N__12027\,
            lcout => \uu2.mem0.g0_7_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_58_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011101111"
        )
    port map (
            in0 => \N__12428\,
            in1 => \N__11994\,
            in2 => \N__15190\,
            in3 => \N__12015\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_38_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__16047\,
            in1 => \_gnd_net_\,
            in2 => \N__12009\,
            in3 => \N__12006\,
            lcout => \uu2.mem0.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI43641_162_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12216\,
            in1 => \N__13676\,
            in2 => \_gnd_net_\,
            in3 => \N__12245\,
            lcout => \uu2.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_73_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12594\,
            in2 => \_gnd_net_\,
            in3 => \N__12215\,
            lcout => \uu2.mem0.m317_0_a6_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_rep1_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__12595\,
            in1 => \N__12772\,
            in2 => \N__12367\,
            in3 => \N__12512\,
            lcout => \uu2.w_addr_displaying_4_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__18660\
        );

    \uu2.w_addr_displaying_4_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__12447\,
            in1 => \N__12354\,
            in2 => \N__12777\,
            in3 => \N__12511\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__18660\
        );

    \uu2.w_addr_displaying_fast_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12358\,
            in1 => \N__12776\,
            in2 => \N__12513\,
            in3 => \N__12491\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4_rep1C_net\,
            ce => 'H',
            sr => \N__18660\
        );

    \uu2.w_addr_displaying_2_rep1_RNI01H61_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13912\,
            in1 => \N__12427\,
            in2 => \_gnd_net_\,
            in3 => \N__12353\,
            lcout => \uu2.N_9_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_75_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12208\,
            in1 => \N__13677\,
            in2 => \_gnd_net_\,
            in3 => \N__12246\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_54_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__15124\,
            in1 => \N__12228\,
            in2 => \N__12231\,
            in3 => \N__12601\,
            lcout => \uu2.mem0.m317_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_76_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12207\,
            in1 => \N__15973\,
            in2 => \N__12607\,
            in3 => \N__16041\,
            lcout => \uu2.mem0.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_72_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15966\,
            in2 => \_gnd_net_\,
            in3 => \N__12209\,
            lcout => OPEN,
            ltout => \uu2.mem0.m317_0_a6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_51_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__12599\,
            in1 => \N__12162\,
            in2 => \N__12639\,
            in3 => \N__12636\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_11_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_29_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12627\,
            in1 => \N__15003\,
            in2 => \N__12621\,
            in3 => \N__12564\,
            lcout => \uu2.mem0.N_6_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_53_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__12600\,
            in1 => \N__16115\,
            in2 => \N__15158\,
            in3 => \N__12570\,
            lcout => \uu2.mem0.N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_31_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15313\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15560\,
            lcout => \uu2.mem0.g1_2_2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_34_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13083\,
            in2 => \_gnd_net_\,
            in3 => \N__14951\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.bitmap_69_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14952\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13074\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.bitmap_197_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12849\,
            in2 => \_gnd_net_\,
            in3 => \N__14948\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.bitmap_290_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14949\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12537\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.bitmap_308_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17574\,
            in2 => \_gnd_net_\,
            in3 => \N__14950\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.w_addr_displaying_2_rep1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12808\,
            in1 => \N__13887\,
            in2 => \_gnd_net_\,
            in3 => \N__15472\,
            lcout => \uu2.w_addr_displaying_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.w_addr_displaying_fast_2_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__15473\,
            in1 => \N__12809\,
            in2 => \_gnd_net_\,
            in3 => \N__12832\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \uu2.w_addr_displaying_2_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__12807\,
            in1 => \N__12727\,
            in2 => \_gnd_net_\,
            in3 => \N__15471\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_34C_net\,
            ce => 'H',
            sr => \N__18654\
        );

    \Lab_UT.bcd2segment2.segmentUQ_6_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100111100001"
        )
    port map (
            in0 => \N__19432\,
            in1 => \N__18171\,
            in2 => \N__18021\,
            in3 => \N__18089\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment2.segmentUQ_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_180_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12675\,
            in3 => \N__14900\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_180C_net\,
            ce => 'H',
            sr => \N__18658\
        );

    \uu2.bitmap_52_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12672\,
            in2 => \_gnd_net_\,
            in3 => \N__14902\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_180C_net\,
            ce => 'H',
            sr => \N__18658\
        );

    \Lab_UT.bcd2segment2.segment_0_1_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__19431\,
            in1 => \N__18170\,
            in2 => \N__18020\,
            in3 => \N__18087\,
            lcout => \Lab_UT.bcd2segment2.segment_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_0_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111101111"
        )
    port map (
            in0 => \N__18088\,
            in1 => \N__18003\,
            in2 => \N__18179\,
            in3 => \N__19433\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment2.segment_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14901\,
            in1 => \_gnd_net_\,
            in2 => \N__12666\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_180C_net\,
            ce => 'H',
            sr => \N__18658\
        );

    \uu2.mem0.ram512X8_inst_RNO_89_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12650\,
            in1 => \N__13232\,
            in2 => \_gnd_net_\,
            in3 => \N__13216\,
            lcout => \uu2.mem0.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m39_e_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13048\,
            in1 => \N__16229\,
            in2 => \N__16387\,
            in3 => \N__18743\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.m39_eZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m39_e_3_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12889\,
            in2 => \N__13200\,
            in3 => \N__12989\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.m39_eZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__13130\,
            in1 => \N__18777\,
            in2 => \N__13197\,
            in3 => \N__18745\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18453\,
            ce => 'H',
            sr => \N__18223\
        );

    \Lab_UT.didp.ce_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__16230\,
            in1 => \N__13126\,
            in2 => \_gnd_net_\,
            in3 => \N__18776\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18453\,
            ce => 'H',
            sr => \N__18223\
        );

    \Lab_UT.didp.reset_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__18775\,
            in1 => \N__16231\,
            in2 => \N__13131\,
            in3 => \N__18744\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18453\,
            ce => 'H',
            sr => \N__18223\
        );

    \Lab_UT.bcd2segment1.m76_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000110010000"
        )
    port map (
            in0 => \N__13043\,
            in1 => \N__12987\,
            in2 => \N__16382\,
            in3 => \N__12887\,
            lcout => \Lab_UT.bcd2segment1.N_181\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m76_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011110011111"
        )
    port map (
            in0 => \N__12986\,
            in1 => \N__16363\,
            in2 => \N__12902\,
            in3 => \N__13042\,
            lcout => \Lab_UT.bcd2segment1.N_229\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m81_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111111011"
        )
    port map (
            in0 => \N__13044\,
            in1 => \N__12988\,
            in2 => \N__16383\,
            in3 => \N__12888\,
            lcout => \Lab_UT.bcd2segment1.N_233\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13239\,
            in2 => \_gnd_net_\,
            in3 => \N__13408\,
            lcout => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\,
            ltout => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIQ35U8_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__13409\,
            in1 => \N__17874\,
            in2 => \N__13332\,
            in3 => \N__13456\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_0\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIFPRO41_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__13265\,
            in1 => \N__13292\,
            in2 => \N__13317\,
            in3 => \N__13304\,
            lcout => \Lab_UT.dictrl.un1_state_21_reti_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIQCSRA_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__17340\,
            in1 => \N__17875\,
            in2 => \N__17305\,
            in3 => \N__17525\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNI2AJ17_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__16998\,
            in1 => \N__16959\,
            in2 => \N__17886\,
            in3 => \N__16936\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_3\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIR8QUG_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13275\,
            in3 => \N__13264\,
            lcout => \Lab_UT.dictrl.dicRun_2_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__13457\,
            in1 => \N__17548\,
            in2 => \N__13475\,
            in3 => \N__13410\,
            lcout => \Lab_UT.dictrl.next_state_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18446\,
            ce => \N__17493\,
            sr => \N__13428\
        );

    \Lab_UT.dictrl.state_0_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__17946\,
            in1 => \N__17912\,
            in2 => \N__17876\,
            in3 => \N__17803\,
            lcout => \Lab_UT.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18439\,
            ce => 'H',
            sr => \N__18694\
        );

    \Lab_UT.dictrl.state_0_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__17002\,
            in1 => \N__16937\,
            in2 => \N__16977\,
            in3 => \N__17861\,
            lcout => \Lab_UT.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18439\,
            ce => 'H',
            sr => \N__18694\
        );

    \Lab_UT.dictrl.state_ret_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__17521\,
            in1 => \N__17859\,
            in2 => \N__17306\,
            in3 => \N__17339\,
            lcout => \Lab_UT.state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18439\,
            ce => 'H',
            sr => \N__18694\
        );

    \Lab_UT.dictrl.state_0_0_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__17860\,
            in1 => \N__13407\,
            in2 => \N__13476\,
            in3 => \N__13458\,
            lcout => \Lab_UT.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18439\,
            ce => 'H',
            sr => \N__18694\
        );

    \buart.Z_rx.bitcount_RNO_0_3_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001011011110"
        )
    port map (
            in0 => \N__17410\,
            in1 => \N__17368\,
            in2 => \N__16149\,
            in3 => \N__16483\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__16484\,
            in1 => \N__17021\,
            in2 => \N__13431\,
            in3 => \N__17411\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18439\,
            ce => 'H',
            sr => \N__18694\
        );

    \Lab_UT.bcd2segment1.m72_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__18894\,
            in1 => \N__13505\,
            in2 => \N__13389\,
            in3 => \N__16878\,
            lcout => \Lab_UT.m72_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIDH8U_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__13506\,
            in1 => \N__18955\,
            in2 => \N__16893\,
            in3 => \N__18896\,
            lcout => \Lab_UT.dictrl.state_0_RNIDH8UZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m29_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13531\,
            in2 => \_gnd_net_\,
            in3 => \N__13766\,
            lcout => \Lab_UT.un1_state_13\,
            ltout => \Lab_UT.un1_state_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_RNIAD2V_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__17773\,
            in1 => \N__18893\,
            in2 => \N__13380\,
            in3 => \N__13338\,
            lcout => \Lab_UT.dictrl.state_ret_1_RNIAD2VZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNI065O1_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__13376\,
            in1 => \N__13359\,
            in2 => \_gnd_net_\,
            in3 => \N__17139\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIENNE_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13504\,
            in2 => \_gnd_net_\,
            in3 => \N__16877\,
            lcout => \Lab_UT.dictrl.un1_state_11\,
            ltout => \Lab_UT.dictrl.un1_state_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_RNITFCD1_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__17774\,
            in1 => \N__18954\,
            in2 => \N__13650\,
            in3 => \N__18895\,
            lcout => \Lab_UT.dictrl.state_ret_1_RNITFCDZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m47_e_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18903\,
            in1 => \N__17775\,
            in2 => \N__13772\,
            in3 => \N__16884\,
            lcout => \Lab_UT.bcd2segment1.N_264\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m68_0_ns_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__16883\,
            in1 => \N__13761\,
            in2 => \_gnd_net_\,
            in3 => \N__18902\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.m68_0_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m68_0_ns_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__18960\,
            in1 => \N__13543\,
            in2 => \N__13596\,
            in3 => \N__13517\,
            lcout => \Lab_UT.m68_0_ns\,
            ltout => \Lab_UT.m68_0_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIO00A3_3_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111010"
        )
    port map (
            in0 => \N__13544\,
            in1 => \N__13593\,
            in2 => \N__13569\,
            in3 => \N__13566\,
            lcout => \Lab_UT.dictrl.next_state_set_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIFOTF_3_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__18901\,
            in1 => \N__18959\,
            in2 => \_gnd_net_\,
            in3 => \N__13542\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_RNIFOTFZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIB7JE1_1_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13518\,
            in1 => \_gnd_net_\,
            in2 => \N__13482\,
            in3 => \N__13731\,
            lcout => \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1\,
            ltout => \Lab_UT.dictrl.state_0_RNIB7JE1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__17887\,
            in1 => \N__17307\,
            in2 => \N__13479\,
            in3 => \N__17520\,
            lcout => \Lab_UT.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18429\,
            ce => 'H',
            sr => \N__18695\
        );

    \Lab_UT.dictrl.state_0_RNIEI8U_2_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__16882\,
            in1 => \N__13762\,
            in2 => \N__18967\,
            in3 => \N__18900\,
            lcout => \Lab_UT.dictrl.state_0_RNIEI8UZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_3_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111100010"
        )
    port map (
            in0 => \N__19350\,
            in1 => \N__19286\,
            in2 => \N__19182\,
            in3 => \N__19074\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_314_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13725\,
            in3 => \N__14976\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__18668\
        );

    \uu2.bitmap_87_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14978\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13722\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__18668\
        );

    \uu2.bitmap_RNI672H_84_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110011101"
        )
    port map (
            in0 => \N__13981\,
            in1 => \N__15050\,
            in2 => \N__13695\,
            in3 => \N__13707\,
            lcout => \uu2.m76_am_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_84_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14977\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17589\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__18668\
        );

    \uu2.w_addr_displaying_fast_7_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15310\,
            in1 => \N__15477\,
            in2 => \N__15397\,
            in3 => \N__15051\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__18668\
        );

    \uu2.bitmap_168_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13686\,
            in2 => \_gnd_net_\,
            in3 => \N__14986\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__18667\
        );

    \Lab_UT.bcd2segment1.m109_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011110010"
        )
    port map (
            in0 => \N__14267\,
            in1 => \N__14178\,
            in2 => \N__14100\,
            in3 => \N__16262\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_246_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_72_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13653\,
            in3 => \N__14988\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__18667\
        );

    \Lab_UT.bcd2segment1.m113_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111101010"
        )
    port map (
            in0 => \N__14268\,
            in1 => \N__14179\,
            in2 => \N__14101\,
            in3 => \N__16263\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.N_248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_200_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14010\,
            in3 => \N__14987\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__18667\
        );

    \uu2.bitmap_RNI65TM_72_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100111101"
        )
    port map (
            in0 => \N__14007\,
            in1 => \N__15043\,
            in2 => \N__13985\,
            in3 => \N__14001\,
            lcout => \uu2.m76_bm_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_0_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13980\,
            in2 => \_gnd_net_\,
            in3 => \N__15470\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__18667\
        );

    \uu2.mem0.ram512X8_inst_RNO_26_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15542\,
            in1 => \N__14621\,
            in2 => \N__15312\,
            in3 => \N__15112\,
            lcout => \uu2.mem0.g1_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_43_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111001011010"
        )
    port map (
            in0 => \N__15113\,
            in1 => \N__15281\,
            in2 => \N__14650\,
            in3 => \N__15543\,
            lcout => \uu2.mem0.g2_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_63_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111101100"
        )
    port map (
            in0 => \N__15541\,
            in1 => \N__14620\,
            in2 => \N__15311\,
            in3 => \N__15111\,
            lcout => \uu2.mem0.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_68_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111101110"
        )
    port map (
            in0 => \N__13908\,
            in1 => \N__16119\,
            in2 => \_gnd_net_\,
            in3 => \N__13833\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_68_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_45_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__14731\,
            in1 => \_gnd_net_\,
            in2 => \N__14700\,
            in3 => \N__14691\,
            lcout => \uu2.mem0.bitmap_pmux_u_i_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_69_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__15110\,
            in1 => \N__15274\,
            in2 => \N__14649\,
            in3 => \N__15540\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_ness_6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110101010"
        )
    port map (
            in0 => \N__15283\,
            in1 => \N__14625\,
            in2 => \N__15196\,
            in3 => \N__15374\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_ness_6C_net\,
            ce => \N__14580\,
            sr => \N__18665\
        );

    \uu2.w_addr_displaying_nesr_8_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15373\,
            in1 => \N__15179\,
            in2 => \N__14651\,
            in3 => \N__15282\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_ness_6C_net\,
            ce => \N__14580\,
            sr => \N__18665\
        );

    \uu2.mem0.ram512X8_inst_RNO_49_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14802\,
            in1 => \N__15309\,
            in2 => \N__15993\,
            in3 => \N__15538\,
            lcout => OPEN,
            ltout => \uu2.mem0.G_13_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_27_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001000000"
        )
    port map (
            in0 => \N__15672\,
            in1 => \N__15714\,
            in2 => \N__14544\,
            in3 => \N__14541\,
            lcout => OPEN,
            ltout => \uu2.mem0.G_13_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__14530\,
            in1 => \N__14421\,
            in2 => \N__14400\,
            in3 => \N__14384\,
            lcout => \uu2.mem0.G_13_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_86_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000101"
        )
    port map (
            in0 => \N__15537\,
            in1 => \N__15977\,
            in2 => \N__14805\,
            in3 => \N__15259\,
            lcout => \uu2.mem0.bitmap_pmux_u_i_4_0_N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI59BR1_5_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15715\,
            in1 => \N__15673\,
            in2 => \_gnd_net_\,
            in3 => \N__15539\,
            lcout => \uu2.N_12_i\,
            ltout => \uu2.N_12_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15476\,
            in1 => \N__15261\,
            in2 => \N__15720\,
            in3 => \N__15981\,
            lcout => \uu2.w_addr_displaying_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7_rep1C_net\,
            ce => 'H',
            sr => \N__18662\
        );

    \uu2.w_addr_displaying_5_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__15716\,
            in1 => \N__15674\,
            in2 => \N__15579\,
            in3 => \N__15474\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7_rep1C_net\,
            ce => 'H',
            sr => \N__18662\
        );

    \uu2.w_addr_displaying_7_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__15475\,
            in1 => \N__15149\,
            in2 => \N__15386\,
            in3 => \N__15260\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_7_rep1C_net\,
            ce => 'H',
            sr => \N__18662\
        );

    \uu2.bitmap_RNIKGSI_58_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14997\,
            in1 => \N__15052\,
            in2 => \_gnd_net_\,
            in3 => \N__14823\,
            lcout => \uu2.N_272\,
            ltout => \uu2.N_272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_52_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__14817\,
            in1 => \N__14804\,
            in2 => \N__15012\,
            in3 => \N__15009\,
            lcout => \uu2.mem0.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_58_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17607\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14975\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_58C_net\,
            ce => 'H',
            sr => \N__18661\
        );

    \uu2.bitmap_186_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17598\,
            in2 => \_gnd_net_\,
            in3 => \N__14974\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_58C_net\,
            ce => 'H',
            sr => \N__18661\
        );

    \uu2.mem0.ram512X8_inst_RNO_81_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14816\,
            in1 => \N__14803\,
            in2 => \_gnd_net_\,
            in3 => \N__14742\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_56_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16118\,
            in2 => \N__16050\,
            in3 => \N__16020\,
            lcout => \uu2.mem0.N_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__17227\,
            in1 => \N__16563\,
            in2 => \N__17039\,
            in3 => \N__16511\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \buart.Z_rx.bitcount_4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__16510\,
            in1 => \N__17038\,
            in2 => \N__17273\,
            in3 => \N__16128\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \buart.Z_rx.bitcount_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__16524\,
            in1 => \N__17449\,
            in2 => \N__17040\,
            in3 => \N__16512\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \buart.Z_rx.bitcount_2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__16509\,
            in1 => \N__17037\,
            in2 => \N__17182\,
            in3 => \N__16419\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \uu2.mem0.ram512X8_inst_RNO_80_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15982\,
            in1 => \N__16037\,
            in2 => \_gnd_net_\,
            in3 => \N__16026\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_82_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__16007\,
            in1 => \N__15983\,
            in2 => \_gnd_net_\,
            in3 => \N__15917\,
            lcout => \uu2.mem0.N_98_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_2_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__15795\,
            in1 => \N__15868\,
            in2 => \N__15849\,
            in3 => \N__15737\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \uu2.r_addr_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__15736\,
            in1 => \N__15844\,
            in2 => \_gnd_net_\,
            in3 => \N__15794\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18476\,
            ce => 'H',
            sr => \N__18692\
        );

    \Lab_UT.didp.ce_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__19069\,
            in1 => \N__19367\,
            in2 => \N__19177\,
            in3 => \N__19281\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18468\,
            ce => 'H',
            sr => \N__18235\
        );

    \Lab_UT.bcd2segment1.m53_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__16832\,
            in1 => \N__19068\,
            in2 => \_gnd_net_\,
            in3 => \N__16397\,
            lcout => \Lab_UT.bcd2segment1.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18822\,
            in1 => \N__19434\,
            in2 => \N__18111\,
            in3 => \N__18095\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18468\,
            ce => 'H',
            sr => \N__18235\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16279\,
            in2 => \_gnd_net_\,
            in3 => \N__16253\,
            lcout => \Lab_UT.didp.countrce3.q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17230\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_10_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17453\,
            in2 => \_gnd_net_\,
            in3 => \N__16155\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17197\,
            in3 => \N__16152\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17415\,
            in3 => \N__16134\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_4_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011101110010"
        )
    port map (
            in0 => \N__17366\,
            in1 => \N__16491\,
            in2 => \N__17274\,
            in3 => \N__16131\,
            lcout => \buart.Z_rx.bitcount_lm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m42_bm_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001011"
        )
    port map (
            in0 => \N__16848\,
            in1 => \N__16821\,
            in2 => \N__16728\,
            in3 => \N__18180\,
            lcout => \Lab_UT.bcd2segment1.m42_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__16490\,
            in1 => \N__16599\,
            in2 => \N__17235\,
            in3 => \N__17367\,
            lcout => \buart.Z_rx.bitcount_lm_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIMK771_4_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17451\,
            in1 => \N__17269\,
            in2 => \N__17198\,
            in3 => \N__17409\,
            lcout => OPEN,
            ltout => \buart.Z_rx.un1_sample_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIC77M1_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17098\,
            in1 => \N__17127\,
            in2 => \N__16554\,
            in3 => \N__17234\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__16972\,
            in1 => \N__17006\,
            in2 => \N__17561\,
            in3 => \N__16938\,
            lcout => \Lab_UT.dictrl.next_state_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18454\,
            ce => \N__17495\,
            sr => \N__16542\
        );

    \buart.Z_rx.bitcount_RNIAPJJ_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17404\,
            in2 => \_gnd_net_\,
            in3 => \N__17450\,
            lcout => \buart.Z_rx.idle_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011011110110"
        )
    port map (
            in0 => \N__17452\,
            in1 => \N__16530\,
            in2 => \N__17373\,
            in3 => \N__16488\,
            lcout => \buart.Z_rx.bitcount_lm_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__16489\,
            in1 => \N__16425\,
            in2 => \N__17199\,
            in3 => \N__17372\,
            lcout => \buart.Z_rx.bitcount_lm_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_2_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__17298\,
            in1 => \N__17338\,
            in2 => \N__17565\,
            in3 => \N__17529\,
            lcout => \Lab_UT.dictrl.next_state_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18447\,
            ce => \N__17496\,
            sr => \N__17472\
        );

    \buart.Z_rx.bitcount_RNIBQJJ_4_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17454\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17268\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_0_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__17186\,
            in1 => \N__17229\,
            in2 => \N__17418\,
            in3 => \N__17405\,
            lcout => bu_rx_data_rdy,
            ltout => \bu_rx_data_rdy_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIIU223_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17376\,
            in3 => \N__17138\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI9T1T1_2_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17313\,
            lcout => \Lab_UT.dictrl.next_state_RNI9T1T1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_4_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17267\,
            in1 => \N__17228\,
            in2 => \N__17196\,
            in3 => \N__17145\,
            lcout => \buart.Z_rx.idle\,
            ltout => \buart.Z_rx.idle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNILM873_0_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__17123\,
            in1 => \N__17099\,
            in2 => \N__17061\,
            in3 => \N__17054\,
            lcout => \buart.Z_rx.bitcountlde_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001111110011"
        )
    port map (
            in0 => \N__17010\,
            in1 => \N__16976\,
            in2 => \N__17895\,
            in3 => \N__16935\,
            lcout => \Lab_UT.state_i_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18440\,
            ce => 'H',
            sr => \N__18696\
        );

    \Lab_UT.dictrl.state_ret_1_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001111110011"
        )
    port map (
            in0 => \N__17947\,
            in1 => \N__17919\,
            in2 => \N__17894\,
            in3 => \N__17805\,
            lcout => \Lab_UT.state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18440\,
            ce => 'H',
            sr => \N__18696\
        );

    \buart.Z_rx.shifter_2_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17756\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18434\,
            ce => \N__17652\,
            sr => \N__18713\
        );

    \Lab_UT.bcd2segment1.segment_0_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__19313\,
            in1 => \N__19226\,
            in2 => \N__19141\,
            in3 => \N__19024\,
            lcout => \Lab_UT.bcd2segment1.segment_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m96_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__19312\,
            in1 => \N__19227\,
            in2 => \N__19140\,
            in3 => \N__19025\,
            lcout => \Lab_UT.bcd2segment1.N_192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__18796\,
            in1 => \N__18844\,
            in2 => \_gnd_net_\,
            in3 => \N__19038\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_5_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111000010"
        )
    port map (
            in0 => \N__18080\,
            in1 => \N__19422\,
            in2 => \N__18017\,
            in3 => \N__18159\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010001010000"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__19039\,
            in2 => \N__19264\,
            in3 => \N__18845\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.un1_num_5_2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18083\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18160\,
            lcout => \Lab_UT.three_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100111100010"
        )
    port map (
            in0 => \N__19424\,
            in1 => \N__18157\,
            in2 => \N__18019\,
            in3 => \N__18082\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segmentUQ_4_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101110"
        )
    port map (
            in0 => \N__18081\,
            in1 => \N__19423\,
            in2 => \N__18018\,
            in3 => \N__18158\,
            lcout => \Lab_UT.bcd2segment2.segmentUQ_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m1_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19243\,
            in2 => \_gnd_net_\,
            in3 => \N__19037\,
            lcout => OPEN,
            ltout => \Lab_UT.three_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__18846\,
            in1 => \N__18798\,
            in2 => \N__18183\,
            in3 => \N__19329\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18485\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__18085\,
            in1 => \N__18522\,
            in2 => \_gnd_net_\,
            in3 => \N__19467\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__18162\,
            in1 => \N__18526\,
            in2 => \N__19473\,
            in3 => \N__18086\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI4V78_3_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18015\,
            in2 => \_gnd_net_\,
            in3 => \N__18161\,
            lcout => \Lab_UT.didp.countrce2.un15_ce_2\,
            ltout => \Lab_UT.didp.countrce2.un15_ce_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI84NN1_2_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18814\,
            in1 => \N__19428\,
            in2 => \N__18099\,
            in3 => \N__18084\,
            lcout => \Lab_UT.q_RNI84NN1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19451\,
            in2 => \_gnd_net_\,
            in3 => \N__19429\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__18527\,
            in1 => \N__19468\,
            in2 => \N__18030\,
            in3 => \N__18016\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__19472\,
            in1 => \N__19452\,
            in2 => \N__18528\,
            in3 => \N__19430\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__19054\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__19260\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__19115\,
            in1 => \N__18795\,
            in2 => \N__19371\,
            in3 => \N__18843\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.m5_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19338\,
            in1 => \N__19256\,
            in2 => \N__19136\,
            in3 => \N__19053\,
            lcout => \Lab_UT.nine\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_0_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__18968\,
            in2 => \_gnd_net_\,
            in3 => \N__18909\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18461\,
            ce => 'H',
            sr => \N__18246\
        );

    \Lab_UT.didp.reset_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18815\,
            in2 => \_gnd_net_\,
            in3 => \N__18750\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18461\,
            ce => 'H',
            sr => \N__18246\
        );

    \Lab_UT.didp.reset_1_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18766\,
            in2 => \_gnd_net_\,
            in3 => \N__18749\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18486\,
            ce => 'H',
            sr => \N__18242\
        );
end \INTERFACE\;
