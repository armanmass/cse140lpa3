-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 19 2019 07:46:31

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18318\ : std_logic;
signal \N__18317\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18305\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18245\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18119\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18095\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18092\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18089\ : std_logic;
signal \N__18088\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18085\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18065\ : std_logic;
signal \N__18064\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18062\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18059\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18041\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18038\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18035\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17844\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17833\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17826\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17811\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17787\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17784\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17781\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17645\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17642\ : std_logic;
signal \N__17639\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17603\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17550\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17547\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17544\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17520\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17348\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17336\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17303\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17249\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17240\ : std_logic;
signal \N__17231\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17153\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17123\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17043\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17009\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16874\ : std_logic;
signal \N__16871\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16820\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16805\ : std_logic;
signal \N__16802\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16574\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16568\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16553\ : std_logic;
signal \N__16550\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16520\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16499\ : std_logic;
signal \N__16496\ : std_logic;
signal \N__16493\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16399\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16387\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16313\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16310\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16292\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16262\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16247\ : std_logic;
signal \N__16244\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16220\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16160\ : std_logic;
signal \N__16157\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16079\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16027\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15947\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15820\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15788\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15753\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15728\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15672\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15526\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15265\ : std_logic;
signal \N__15262\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15122\ : std_logic;
signal \N__15121\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15112\ : std_logic;
signal \N__15109\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15091\ : std_logic;
signal \N__15088\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15056\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14915\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14909\ : std_logic;
signal \N__14906\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14888\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14734\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14664\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14311\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14236\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14093\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13934\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13751\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13712\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13706\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13398\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12649\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10241\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7730\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7533\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal \uu2.un284_ci_cascade_\ : std_logic;
signal \uu2.un306_ci_cascade_\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_11_cascade_\ : std_logic;
signal \uu0.un4_l_count_16_cascade_\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un55_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \uu0.un4_l_count_0_8_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \bfn_2_3_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0_cascade_\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.un1_l_count_2_2_cascade_\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.un1_l_count_1_2_0_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \uu0.sec_clkDZ0\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu0.un88_ci_3_cascade_\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \resetGen.escKeyZ0_cascade_\ : std_logic;
signal \resetGen.un252_ci_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen.reset_countZ0Z_0\ : std_logic;
signal \resetGen.reset_countZ0Z_1\ : std_logic;
signal \resetGen.reset_countZ0Z_2\ : std_logic;
signal \resetGen.un241_ci\ : std_logic;
signal \resetGen.reset_count_2_0_4\ : std_logic;
signal \resetGen.escKeyZ0\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.un220_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.trig_rd_is_det_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.mem0.N_77_i\ : std_logic;
signal \uu2.mem0.w_data_i_a3_1_0_cascade_\ : std_logic;
signal \uu2.mem0.N_79_i_0\ : std_logic;
signal clk : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.N_75_i\ : std_logic;
signal \uu2.N_361\ : std_logic;
signal \uu2.N_361_cascade_\ : std_logic;
signal \uu2.mem0.w_data_4\ : std_logic;
signal \uu2.mem0.N_69_i\ : std_logic;
signal \uu2.mem0.w_data_0_a3_0_4\ : std_logic;
signal \uu2.N_61_cascade_\ : std_logic;
signal \uu2.mem0.un51_w_data_displaying_cascade_\ : std_logic;
signal \uu2.mem0.w_data_5\ : std_logic;
signal \uu2.mem0.w_data_6\ : std_logic;
signal \uu2.mem0.N_71_i\ : std_logic;
signal \uu2.mem0.w_data_1\ : std_logic;
signal \uu2.mem0.N_76_i_0\ : std_logic;
signal \uu2.mem0.N_2166_0_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_3\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_42\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_43\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_\ : std_logic;
signal \uu2.bitmap_RNIMQ601Z0Z_58_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \INVuu2.bitmap_186C_net\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \uu2.bitmap_RNI8LB51Z0Z_186\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \INVuu2.bitmap_308C_net\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.mem0.N_70_i\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.bitmap_pmux_20_ns_1_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_0Z0Z_2\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \Lab_UT.bcd2segment4.N_217\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_i_1Z0Z_5\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \INVuu2.bitmap_197C_net\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_\ : std_logic;
signal \uu2.mem0.g1_2_0\ : std_logic;
signal \uu2.N_40_0\ : std_logic;
signal \uu2.N_48_i_0\ : std_logic;
signal \uu2.N_404\ : std_logic;
signal \uu2.mem0.g1_1_1_0\ : std_logic;
signal \uu2.N_404_cascade_\ : std_logic;
signal \uu2.mem0.bitmap_pmux_1_0_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_42_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_46\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_\ : std_logic;
signal \uu2.g2_0_0\ : std_logic;
signal \uu2.mem0.g1_6_cascade_\ : std_logic;
signal \uu2.mem0.N_1201_0_0_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20_0\ : std_logic;
signal \uu2.bitmap_pmux_19_i_m2_ns_1\ : std_logic;
signal \uu2.N_55_0\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_20_1_0_1\ : std_logic;
signal \uu2.mem0.N_2166_1_0_1\ : std_logic;
signal \uu2.mem0.N_247_0_cascade_\ : std_logic;
signal \uu2.mem0.N_2171_1_0_1_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7\ : std_logic;
signal \uu2.mem0.N_397_1_0_1\ : std_logic;
signal \uu2.mem0.g1_3_0\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.N_247_cascade_\ : std_logic;
signal \uu2.N_2171_0\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_44\ : std_logic;
signal \Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.N_383\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \INVuu2.bitmap_290C_net\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmap_pmux_15_i_m2_ns_1\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_54_mux_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_15\ : std_logic;
signal \uu2.N_395_cascade_\ : std_logic;
signal \uu2.N_56\ : std_logic;
signal \uu2.N_401\ : std_logic;
signal \buart.Z_rx.idle_1_cascade_\ : std_logic;
signal \buart.Z_rx.valid_1_cascade_\ : std_logic;
signal \buart.Z_rx.hhZ0Z_1\ : std_logic;
signal \buart.Z_rx.hhZ0Z_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \uu2.N_150_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \INVuu2.w_addr_user_nesr_6C_net\ : std_logic;
signal \uu2.mem0.N_78_i_0\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.N_93\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_0Z0Z_2\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \INVuu2.w_addr_displaying_4C_net\ : std_logic;
signal \uu2.mem0.g0_7_3_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_27_ns_1_0\ : std_logic;
signal \uu2.mem0.g0_6_4\ : std_logic;
signal \uu2.mem0.g0_6_5_cascade_\ : std_logic;
signal \uu2.un426_ci\ : std_logic;
signal \INVuu2.w_addr_displaying_2_rep1C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \uu2.N_46_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_fast_nesr_8C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_\ : std_logic;
signal \uu2.N_4_cascade_\ : std_logic;
signal \uu2.g0_17_1\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \uu2.N_5\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \INVuu2.bitmap_200C_net\ : std_logic;
signal \Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.bitmap_RNISSSNZ0Z_162\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \INVuu2.bitmap_168C_net\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_i_0Z0Z_1\ : std_logic;
signal \Lab_UT.bcd2segment3.segment_i_0Z0Z_2\ : std_logic;
signal \resetGen.escKeyZ0Z_3\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \buart.Z_rx.N_27_0_i_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_lm_0_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_lm_1_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_lm_2_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_rx.bitcount_lm_4\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_4\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.N_27_0_i\ : std_logic;
signal \buart.Z_rx.bitcount_lm_3_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_3\ : std_logic;
signal \uu2.N_153\ : std_logic;
signal \uu2.N_90_cascade_\ : std_logic;
signal \uu2.N_105\ : std_logic;
signal \uu2.N_90\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \INVuu2.w_addr_user_nesr_3C_net\ : std_logic;
signal \uu2.mem0.N_111\ : std_logic;
signal \uu2.un28_w_addr_user_i_0_0\ : std_logic;
signal \uu2.mem0.N_73_i\ : std_logic;
signal \uu2.un31_w_data_displaying_0_a2_1_cascade_\ : std_logic;
signal \uu2.un31_w_data_displaying\ : std_logic;
signal \uu2.un15_w_data_displaying_6\ : std_logic;
signal \uu2.un15_w_data_displaying_6_cascade_\ : std_logic;
signal \uu2.un49_w_data_displaying_1\ : std_logic;
signal \uu2.un49_w_data_displaying\ : std_logic;
signal \uu2.un15_w_data_displaying_i_i_o2_0\ : std_logic;
signal \uu2.un15_w_data_displaying_i_i_o2_0_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_8C_net\ : std_logic;
signal \uu2.mem0.un49_w_data_displaying_0\ : std_logic;
signal \uu2.mem0.g0_5_5\ : std_logic;
signal \uu2.mem0.un31_w_data_displaying_0\ : std_logic;
signal \uu2.mem0.g1_1_1\ : std_logic;
signal \uu2.w_addr_displaying_7_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_8_repZ0Z1\ : std_logic;
signal \uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_45\ : std_logic;
signal \uu2.w_addr_displaying_2_repZ0Z1\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z1\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_31_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_31_0_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_48\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_\ : std_logic;
signal \uu2.mem0.ram512X8_inst_RNOZ0Z_47\ : std_logic;
signal \uu2.mem0.bitmap_pmux_u_ns_1\ : std_logic;
signal \uu2.mem0.g0_5_3_cascade_\ : std_logic;
signal \uu2.mem0.g0_5_6\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.w_addr_displaying_1_repZ0Z1\ : std_logic;
signal \uu2.N_7_cascade_\ : std_logic;
signal \uu2.N_10\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.N_8\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \INVuu2.bitmap_215C_net\ : std_logic;
signal \Lab_UT.didp.countrce2.N_178\ : std_logic;
signal \Lab_UT.didp.countrce2.N_175\ : std_logic;
signal \Lab_UT.didp.countrce2.N_170\ : std_logic;
signal \Lab_UT.didp.countrce2.N_183\ : std_logic;
signal \Lab_UT.didp.countrce2.N_180\ : std_logic;
signal \Lab_UT.didp.countrce4.N_80_i_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_RNO_0Z0Z_3\ : std_logic;
signal \Lab_UT.bcd2segment4.segment_i_0Z0Z_6\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4_1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_\ : std_logic;
signal \resetGen_escKey_4_cascade_\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\ : std_logic;
signal \resetGen_escKey_2_0\ : std_logic;
signal bu_rx_data_6 : std_logic;
signal bu_rx_data_3 : std_logic;
signal bu_rx_data_7 : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa_cascade_\ : std_logic;
signal \Lab_UT.m37_ns_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_2\ : std_logic;
signal \Lab_UT.m45\ : std_logic;
signal \Lab_UT.m40_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.dicRun_2_reti\ : std_logic;
signal \buart.Z_rx.idle\ : std_logic;
signal bu_rx_data_rdy : std_logic;
signal \buart.Z_rx.bitcountlde_0\ : std_logic;
signal \buart.Z_rx.un1_sample_0\ : std_logic;
signal \buart.Z_rx.ser_clk_2_cascade_\ : std_logic;
signal \buart.Z_rx.bitcountZ0Z_0\ : std_logic;
signal \buart.Z_rx.sample\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.ser_clk_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\ : std_logic;
signal \buart.Z_rx.ser_clk_3\ : std_logic;
signal \buart.Z_rx.startbit\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \Lab_UT.didp.countrce4.q_RNO_0Z0Z_2\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.w_addr_user_3_i_a2_2_6\ : std_logic;
signal \uu2.mem0.N_72_i\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.mem0.N_74_i\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_3_0\ : std_logic;
signal \uu2.N_84_cascade_\ : std_logic;
signal \uu2.N_97\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \uu2.N_97_cascade_\ : std_logic;
signal \uu2.N_159\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \uu2.N_86\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.N_86_cascade_\ : std_logic;
signal \uu2.N_84\ : std_logic;
signal \uu2.w_addr_i_0_tzZ0Z_0\ : std_logic;
signal \uu2.w_addr_i_0_tzZ0Z_0_cascade_\ : std_logic;
signal \uu2.N_61\ : std_logic;
signal \uu2.un21_w_addr_displaying_i\ : std_logic;
signal \uu2.N_49\ : std_logic;
signal \uu2.mem0.g0_7_5_0_cascade_\ : std_logic;
signal \uu2.mem0.un31_w_data_displaying_1_0_0_cascade_\ : std_logic;
signal \uu2.mem0.g1_0_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.mem0.g1_0_1_1\ : std_logic;
signal \uu2.mem0.g1_5_5\ : std_logic;
signal \uu2.w_addr_displaying_3_repZ0Z2\ : std_logic;
signal \uu2.mem0.g0_7_4_0\ : std_logic;
signal \uu2.N_46\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_4\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_3\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_5C_net\ : std_logic;
signal \uu2.un21_w_addr_displaying_i_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.mem0.g0_16_1\ : std_logic;
signal \Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \Lab_UT.nine_cascade_\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_i_0Z0Z_1\ : std_logic;
signal \Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \Lab_UT.three_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_1_sqmuxa\ : std_logic;
signal \Lab_UT.didp.m34_nsZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.next_state16Z0Z_4\ : std_logic;
signal \Lab_UT.m34_ns_cascade_\ : std_logic;
signal \resetGen_escKey_4\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \resetGen.reset_countZ0Z_4\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_3\ : std_logic;
signal \Lab_UT.m34_ns\ : std_logic;
signal \Lab_UT.didp.N_164_cascade_\ : std_logic;
signal \Lab_UT.m42\ : std_logic;
signal \Lab_UT.didp.countrce4.N_88_i\ : std_logic;
signal \Lab_UT.N_68_0\ : std_logic;
signal \Lab_UT.didp.un31_reset_i_a4_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2\ : std_logic;
signal \Lab_UT.m37_ns\ : std_logic;
signal \Lab_UT.Run\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.un1_state_12_cascade_\ : std_logic;
signal \Lab_UT.didp.m37_nsZ0Z_1\ : std_logic;
signal \Lab_UT.state_i_3_1\ : std_logic;
signal \Lab_UT.state_2\ : std_logic;
signal \Lab_UT.state_3\ : std_logic;
signal \Lab_UT.dictrl.un1_state_24_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_out_1\ : std_logic;
signal \Lab_UT.dictrl.un1_state_21_reti_i\ : std_logic;
signal \Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_3_2_cascade_\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_0_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_0\ : std_logic;
signal \Lab_UT.un29_dOutP\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_1\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_1_cascade_\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_3_1\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0\ : std_logic;
signal \Lab_UT.m24\ : std_logic;
signal \Lab_UT.dispString.un22_dOutP\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_3\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_3_3_cascade_\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_0\ : std_logic;
signal \Lab_UT.alarmchar9_cascade_\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_1\ : std_logic;
signal \Lab_UT.zero\ : std_logic;
signal \Lab_UT.didp.countrce3.qPone_3_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.N_79_i_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_3\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.N_207_cascade_\ : std_logic;
signal \Lab_UT.didp.q_RNIIKFH3_3\ : std_logic;
signal \Lab_UT.m40\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI970UZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_set_2\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_2_cascade_\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_2\ : std_logic;
signal \Lab_UT.un3_dOutP\ : std_logic;
signal \Lab_UT.cnt_3\ : std_logic;
signal \Lab_UT.cnt_0\ : std_logic;
signal \Lab_UT.cnt_1\ : std_logic;
signal \Lab_UT.cnt_2\ : std_logic;
signal \Lab_UT.N_204\ : std_logic;
signal \Lab_UT.N_204_cascade_\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.nine\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.three_2\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.didp.countrce2.three_2_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.N_207\ : std_logic;
signal \Lab_UT.didp.q_RNI84NN1_3\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.bcd2segment4.G_64_a0Z0Z_1\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.dictrl.dicRun_2\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \oneSecStrb_i\ : std_logic;
signal \Lab_UT.state_1\ : std_logic;
signal \Lab_UT.dictrl.state_i_3Z0Z_2\ : std_logic;
signal \Lab_UT.state_i_3_3\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.state_ret_3_RNIDH8UZ0\ : std_logic;
signal \Lab_UT.dictrl.state_retZ0Z_4\ : std_logic;
signal \Lab_UT.dictrl.next_state_set\ : std_logic;
signal \Lab_UT.state_0\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_4\ : std_logic;
signal \Lab_UT.alarmchar_2_1_1_cascade_\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_6\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_cascade_\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.G_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstateZ0Z_0\ : std_logic;
signal \Lab_UT.alarmMatch\ : std_logic;
signal \Lab_UT.dictrl.idle\ : std_logic;
signal \Lab_UT.alarmchar10\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1\ : std_logic;
signal \Lab_UT.next_alarmstate4\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\ : std_logic;
signal \Lab_UT.alarmstate_1\ : std_logic;
signal \Lab_UT.alarmchar10_i_2\ : std_logic;
signal \Lab_UT.alarmcharZ0Z_5\ : std_logic;
signal \Lab_UT.alarmstate_0\ : std_logic;
signal \Lab_UT.bcd2segment4.GZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_0_0\ : std_logic;
signal \Lab_UT.un1_next_alarmstate21_0\ : std_logic;
signal \Lab_UT.dictrl.next_alarmstate_1_0\ : std_logic;
signal \Lab_UT.dictrl.alarmstate_i_3_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_g : std_logic;
signal rst_g : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal sd_wire : std_logic;
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    sd <= sd_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__9037\&\N__9412\&\N__9442\&\N__9499\&\N__9532\&\N__9301\&\N__9375\&\N__9339\&\N__9267\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__9457\&\N__8941\&\N__11848\&\N__10600\&\N__12622\&\N__8890\&\N__8926\&\N__8734\&\N__10060\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__8836\&'0'&\N__8842\&'0'&\N__8869\&'0'&\N__8908\&'0'&\N__8863\&'0'&\N__8932\&'0'&\N__8722\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__6901\,
            RESETB => \N__10413\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__18081\,
            RE => \N__10414\,
            WCLKE => \N__8679\,
            WCLK => \N__18080\,
            WE => \N__8689\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18473\,
            DIN => \N__18472\,
            DOUT => \N__18471\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__18473\,
            PADOUT => \N__18472\,
            PADIN => \N__18471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18464\,
            DIN => \N__18463\,
            DOUT => \N__18462\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18464\,
            PADOUT => \N__18463\,
            PADIN => \N__18462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18455\,
            DIN => \N__18454\,
            DOUT => \N__18453\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__18455\,
            PADOUT => \N__18454\,
            PADIN => \N__18453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18446\,
            DIN => \N__18445\,
            DOUT => \N__18444\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__18446\,
            PADOUT => \N__18445\,
            PADIN => \N__18444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18437\,
            DIN => \N__18436\,
            DOUT => \N__18435\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__18437\,
            PADOUT => \N__18436\,
            PADIN => \N__18435\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__18076\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18428\,
            DIN => \N__18427\,
            DOUT => \N__18426\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__18428\,
            PADOUT => \N__18427\,
            PADIN => \N__18426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18419\,
            DIN => \N__18418\,
            DOUT => \N__18417\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__18419\,
            PADOUT => \N__18418\,
            PADIN => \N__18417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18410\,
            DIN => \N__18409\,
            DOUT => \N__18408\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__18410\,
            PADOUT => \N__18409\,
            PADIN => \N__18408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18401\,
            DIN => \N__18400\,
            DOUT => \N__18399\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18401\,
            PADOUT => \N__18400\,
            PADIN => \N__18399\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__18392\,
            DIN => \N__18391\,
            DOUT => \N__18390\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__18392\,
            PADOUT => \N__18391\,
            PADIN => \N__18390\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6913\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4412\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__18370\,
            I => \N__18367\
        );

    \I__4410\ : Odrv4
    port map (
            O => \N__18367\,
            I => \Lab_UT.alarmchar10\
        );

    \I__4409\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18358\
        );

    \I__4408\ : InMux
    port map (
            O => \N__18363\,
            I => \N__18358\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__18358\,
            I => \Lab_UT.dictrl.next_alarmstate_1\
        );

    \I__4406\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18349\
        );

    \I__4405\ : InMux
    port map (
            O => \N__18354\,
            I => \N__18342\
        );

    \I__4404\ : InMux
    port map (
            O => \N__18353\,
            I => \N__18342\
        );

    \I__4403\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18342\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__18349\,
            I => \N__18337\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18337\
        );

    \I__4400\ : Span12Mux_s10_v
    port map (
            O => \N__18337\,
            I => \N__18334\
        );

    \I__4399\ : Odrv12
    port map (
            O => \N__18334\,
            I => \Lab_UT.next_alarmstate4\
        );

    \I__4398\ : InMux
    port map (
            O => \N__18331\,
            I => \N__18327\
        );

    \I__4397\ : InMux
    port map (
            O => \N__18330\,
            I => \N__18324\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__18327\,
            I => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__18324\,
            I => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\
        );

    \I__4394\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18309\
        );

    \I__4393\ : InMux
    port map (
            O => \N__18318\,
            I => \N__18309\
        );

    \I__4392\ : InMux
    port map (
            O => \N__18317\,
            I => \N__18309\
        );

    \I__4391\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18306\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__18309\,
            I => \N__18300\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__18306\,
            I => \N__18297\
        );

    \I__4388\ : InMux
    port map (
            O => \N__18305\,
            I => \N__18290\
        );

    \I__4387\ : InMux
    port map (
            O => \N__18304\,
            I => \N__18290\
        );

    \I__4386\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18290\
        );

    \I__4385\ : Odrv4
    port map (
            O => \N__18300\,
            I => \Lab_UT.alarmstate_1\
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__18297\,
            I => \Lab_UT.alarmstate_1\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__18290\,
            I => \Lab_UT.alarmstate_1\
        );

    \I__4382\ : InMux
    port map (
            O => \N__18283\,
            I => \N__18280\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__18280\,
            I => \Lab_UT.alarmchar10_i_2\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__18277\,
            I => \N__18274\
        );

    \I__4379\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18271\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18268\
        );

    \I__4377\ : Span4Mux_v
    port map (
            O => \N__18268\,
            I => \N__18265\
        );

    \I__4376\ : Odrv4
    port map (
            O => \N__18265\,
            I => \Lab_UT.alarmcharZ0Z_5\
        );

    \I__4375\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18257\
        );

    \I__4374\ : InMux
    port map (
            O => \N__18261\,
            I => \N__18254\
        );

    \I__4373\ : CascadeMux
    port map (
            O => \N__18260\,
            I => \N__18250\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__18257\,
            I => \N__18245\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__18254\,
            I => \N__18245\
        );

    \I__4370\ : InMux
    port map (
            O => \N__18253\,
            I => \N__18242\
        );

    \I__4369\ : InMux
    port map (
            O => \N__18250\,
            I => \N__18239\
        );

    \I__4368\ : Odrv4
    port map (
            O => \N__18245\,
            I => \Lab_UT.alarmstate_0\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__18242\,
            I => \Lab_UT.alarmstate_0\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__18239\,
            I => \Lab_UT.alarmstate_0\
        );

    \I__4365\ : CascadeMux
    port map (
            O => \N__18232\,
            I => \N__18229\
        );

    \I__4364\ : InMux
    port map (
            O => \N__18229\,
            I => \N__18226\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__18226\,
            I => \Lab_UT.bcd2segment4.GZ0Z_1\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__18223\,
            I => \N__18219\
        );

    \I__4361\ : InMux
    port map (
            O => \N__18222\,
            I => \N__18212\
        );

    \I__4360\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18207\
        );

    \I__4359\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18207\
        );

    \I__4358\ : InMux
    port map (
            O => \N__18217\,
            I => \N__18204\
        );

    \I__4357\ : InMux
    port map (
            O => \N__18216\,
            I => \N__18199\
        );

    \I__4356\ : InMux
    port map (
            O => \N__18215\,
            I => \N__18199\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__18212\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__18207\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__18204\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__4352\ : LocalMux
    port map (
            O => \N__18199\,
            I => \Lab_UT.dictrl.next_alarmstate_0_0\
        );

    \I__4351\ : CascadeMux
    port map (
            O => \N__18190\,
            I => \N__18182\
        );

    \I__4350\ : InMux
    port map (
            O => \N__18189\,
            I => \N__18173\
        );

    \I__4349\ : InMux
    port map (
            O => \N__18188\,
            I => \N__18173\
        );

    \I__4348\ : InMux
    port map (
            O => \N__18187\,
            I => \N__18173\
        );

    \I__4347\ : InMux
    port map (
            O => \N__18186\,
            I => \N__18170\
        );

    \I__4346\ : InMux
    port map (
            O => \N__18185\,
            I => \N__18167\
        );

    \I__4345\ : InMux
    port map (
            O => \N__18182\,
            I => \N__18162\
        );

    \I__4344\ : InMux
    port map (
            O => \N__18181\,
            I => \N__18162\
        );

    \I__4343\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18159\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__18173\,
            I => \Lab_UT.un1_next_alarmstate21_0\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__18170\,
            I => \Lab_UT.un1_next_alarmstate21_0\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__18167\,
            I => \Lab_UT.un1_next_alarmstate21_0\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__18162\,
            I => \Lab_UT.un1_next_alarmstate21_0\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__18159\,
            I => \Lab_UT.un1_next_alarmstate21_0\
        );

    \I__4337\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18142\
        );

    \I__4336\ : InMux
    port map (
            O => \N__18147\,
            I => \N__18139\
        );

    \I__4335\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18134\
        );

    \I__4334\ : InMux
    port map (
            O => \N__18145\,
            I => \N__18134\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__18142\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__18139\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__18134\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0\
        );

    \I__4330\ : InMux
    port map (
            O => \N__18127\,
            I => \N__18123\
        );

    \I__4329\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18120\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__18123\,
            I => \N__18115\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__18120\,
            I => \N__18112\
        );

    \I__4326\ : InMux
    port map (
            O => \N__18119\,
            I => \N__18109\
        );

    \I__4325\ : InMux
    port map (
            O => \N__18118\,
            I => \N__18106\
        );

    \I__4324\ : Odrv4
    port map (
            O => \N__18115\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__18112\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__18109\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__18106\,
            I => \Lab_UT.dictrl.alarmstate_i_3_0\
        );

    \I__4320\ : ClkMux
    port map (
            O => \N__18097\,
            I => \N__17863\
        );

    \I__4319\ : ClkMux
    port map (
            O => \N__18096\,
            I => \N__17863\
        );

    \I__4318\ : ClkMux
    port map (
            O => \N__18095\,
            I => \N__17863\
        );

    \I__4317\ : ClkMux
    port map (
            O => \N__18094\,
            I => \N__17863\
        );

    \I__4316\ : ClkMux
    port map (
            O => \N__18093\,
            I => \N__17863\
        );

    \I__4315\ : ClkMux
    port map (
            O => \N__18092\,
            I => \N__17863\
        );

    \I__4314\ : ClkMux
    port map (
            O => \N__18091\,
            I => \N__17863\
        );

    \I__4313\ : ClkMux
    port map (
            O => \N__18090\,
            I => \N__17863\
        );

    \I__4312\ : ClkMux
    port map (
            O => \N__18089\,
            I => \N__17863\
        );

    \I__4311\ : ClkMux
    port map (
            O => \N__18088\,
            I => \N__17863\
        );

    \I__4310\ : ClkMux
    port map (
            O => \N__18087\,
            I => \N__17863\
        );

    \I__4309\ : ClkMux
    port map (
            O => \N__18086\,
            I => \N__17863\
        );

    \I__4308\ : ClkMux
    port map (
            O => \N__18085\,
            I => \N__17863\
        );

    \I__4307\ : ClkMux
    port map (
            O => \N__18084\,
            I => \N__17863\
        );

    \I__4306\ : ClkMux
    port map (
            O => \N__18083\,
            I => \N__17863\
        );

    \I__4305\ : ClkMux
    port map (
            O => \N__18082\,
            I => \N__17863\
        );

    \I__4304\ : ClkMux
    port map (
            O => \N__18081\,
            I => \N__17863\
        );

    \I__4303\ : ClkMux
    port map (
            O => \N__18080\,
            I => \N__17863\
        );

    \I__4302\ : ClkMux
    port map (
            O => \N__18079\,
            I => \N__17863\
        );

    \I__4301\ : ClkMux
    port map (
            O => \N__18078\,
            I => \N__17863\
        );

    \I__4300\ : ClkMux
    port map (
            O => \N__18077\,
            I => \N__17863\
        );

    \I__4299\ : ClkMux
    port map (
            O => \N__18076\,
            I => \N__17863\
        );

    \I__4298\ : ClkMux
    port map (
            O => \N__18075\,
            I => \N__17863\
        );

    \I__4297\ : ClkMux
    port map (
            O => \N__18074\,
            I => \N__17863\
        );

    \I__4296\ : ClkMux
    port map (
            O => \N__18073\,
            I => \N__17863\
        );

    \I__4295\ : ClkMux
    port map (
            O => \N__18072\,
            I => \N__17863\
        );

    \I__4294\ : ClkMux
    port map (
            O => \N__18071\,
            I => \N__17863\
        );

    \I__4293\ : ClkMux
    port map (
            O => \N__18070\,
            I => \N__17863\
        );

    \I__4292\ : ClkMux
    port map (
            O => \N__18069\,
            I => \N__17863\
        );

    \I__4291\ : ClkMux
    port map (
            O => \N__18068\,
            I => \N__17863\
        );

    \I__4290\ : ClkMux
    port map (
            O => \N__18067\,
            I => \N__17863\
        );

    \I__4289\ : ClkMux
    port map (
            O => \N__18066\,
            I => \N__17863\
        );

    \I__4288\ : ClkMux
    port map (
            O => \N__18065\,
            I => \N__17863\
        );

    \I__4287\ : ClkMux
    port map (
            O => \N__18064\,
            I => \N__17863\
        );

    \I__4286\ : ClkMux
    port map (
            O => \N__18063\,
            I => \N__17863\
        );

    \I__4285\ : ClkMux
    port map (
            O => \N__18062\,
            I => \N__17863\
        );

    \I__4284\ : ClkMux
    port map (
            O => \N__18061\,
            I => \N__17863\
        );

    \I__4283\ : ClkMux
    port map (
            O => \N__18060\,
            I => \N__17863\
        );

    \I__4282\ : ClkMux
    port map (
            O => \N__18059\,
            I => \N__17863\
        );

    \I__4281\ : ClkMux
    port map (
            O => \N__18058\,
            I => \N__17863\
        );

    \I__4280\ : ClkMux
    port map (
            O => \N__18057\,
            I => \N__17863\
        );

    \I__4279\ : ClkMux
    port map (
            O => \N__18056\,
            I => \N__17863\
        );

    \I__4278\ : ClkMux
    port map (
            O => \N__18055\,
            I => \N__17863\
        );

    \I__4277\ : ClkMux
    port map (
            O => \N__18054\,
            I => \N__17863\
        );

    \I__4276\ : ClkMux
    port map (
            O => \N__18053\,
            I => \N__17863\
        );

    \I__4275\ : ClkMux
    port map (
            O => \N__18052\,
            I => \N__17863\
        );

    \I__4274\ : ClkMux
    port map (
            O => \N__18051\,
            I => \N__17863\
        );

    \I__4273\ : ClkMux
    port map (
            O => \N__18050\,
            I => \N__17863\
        );

    \I__4272\ : ClkMux
    port map (
            O => \N__18049\,
            I => \N__17863\
        );

    \I__4271\ : ClkMux
    port map (
            O => \N__18048\,
            I => \N__17863\
        );

    \I__4270\ : ClkMux
    port map (
            O => \N__18047\,
            I => \N__17863\
        );

    \I__4269\ : ClkMux
    port map (
            O => \N__18046\,
            I => \N__17863\
        );

    \I__4268\ : ClkMux
    port map (
            O => \N__18045\,
            I => \N__17863\
        );

    \I__4267\ : ClkMux
    port map (
            O => \N__18044\,
            I => \N__17863\
        );

    \I__4266\ : ClkMux
    port map (
            O => \N__18043\,
            I => \N__17863\
        );

    \I__4265\ : ClkMux
    port map (
            O => \N__18042\,
            I => \N__17863\
        );

    \I__4264\ : ClkMux
    port map (
            O => \N__18041\,
            I => \N__17863\
        );

    \I__4263\ : ClkMux
    port map (
            O => \N__18040\,
            I => \N__17863\
        );

    \I__4262\ : ClkMux
    port map (
            O => \N__18039\,
            I => \N__17863\
        );

    \I__4261\ : ClkMux
    port map (
            O => \N__18038\,
            I => \N__17863\
        );

    \I__4260\ : ClkMux
    port map (
            O => \N__18037\,
            I => \N__17863\
        );

    \I__4259\ : ClkMux
    port map (
            O => \N__18036\,
            I => \N__17863\
        );

    \I__4258\ : ClkMux
    port map (
            O => \N__18035\,
            I => \N__17863\
        );

    \I__4257\ : ClkMux
    port map (
            O => \N__18034\,
            I => \N__17863\
        );

    \I__4256\ : ClkMux
    port map (
            O => \N__18033\,
            I => \N__17863\
        );

    \I__4255\ : ClkMux
    port map (
            O => \N__18032\,
            I => \N__17863\
        );

    \I__4254\ : ClkMux
    port map (
            O => \N__18031\,
            I => \N__17863\
        );

    \I__4253\ : ClkMux
    port map (
            O => \N__18030\,
            I => \N__17863\
        );

    \I__4252\ : ClkMux
    port map (
            O => \N__18029\,
            I => \N__17863\
        );

    \I__4251\ : ClkMux
    port map (
            O => \N__18028\,
            I => \N__17863\
        );

    \I__4250\ : ClkMux
    port map (
            O => \N__18027\,
            I => \N__17863\
        );

    \I__4249\ : ClkMux
    port map (
            O => \N__18026\,
            I => \N__17863\
        );

    \I__4248\ : ClkMux
    port map (
            O => \N__18025\,
            I => \N__17863\
        );

    \I__4247\ : ClkMux
    port map (
            O => \N__18024\,
            I => \N__17863\
        );

    \I__4246\ : ClkMux
    port map (
            O => \N__18023\,
            I => \N__17863\
        );

    \I__4245\ : ClkMux
    port map (
            O => \N__18022\,
            I => \N__17863\
        );

    \I__4244\ : ClkMux
    port map (
            O => \N__18021\,
            I => \N__17863\
        );

    \I__4243\ : ClkMux
    port map (
            O => \N__18020\,
            I => \N__17863\
        );

    \I__4242\ : GlobalMux
    port map (
            O => \N__17863\,
            I => \N__17860\
        );

    \I__4241\ : gio2CtrlBuf
    port map (
            O => \N__17860\,
            I => clk_g
        );

    \I__4240\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17847\
        );

    \I__4239\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17847\
        );

    \I__4238\ : InMux
    port map (
            O => \N__17855\,
            I => \N__17844\
        );

    \I__4237\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17841\
        );

    \I__4236\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17838\
        );

    \I__4235\ : InMux
    port map (
            O => \N__17852\,
            I => \N__17835\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17802\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__17844\,
            I => \N__17799\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__17841\,
            I => \N__17796\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__17838\,
            I => \N__17793\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17773\
        );

    \I__4229\ : SRMux
    port map (
            O => \N__17834\,
            I => \N__17668\
        );

    \I__4228\ : SRMux
    port map (
            O => \N__17833\,
            I => \N__17668\
        );

    \I__4227\ : SRMux
    port map (
            O => \N__17832\,
            I => \N__17668\
        );

    \I__4226\ : SRMux
    port map (
            O => \N__17831\,
            I => \N__17668\
        );

    \I__4225\ : SRMux
    port map (
            O => \N__17830\,
            I => \N__17668\
        );

    \I__4224\ : SRMux
    port map (
            O => \N__17829\,
            I => \N__17668\
        );

    \I__4223\ : SRMux
    port map (
            O => \N__17828\,
            I => \N__17668\
        );

    \I__4222\ : SRMux
    port map (
            O => \N__17827\,
            I => \N__17668\
        );

    \I__4221\ : SRMux
    port map (
            O => \N__17826\,
            I => \N__17668\
        );

    \I__4220\ : SRMux
    port map (
            O => \N__17825\,
            I => \N__17668\
        );

    \I__4219\ : SRMux
    port map (
            O => \N__17824\,
            I => \N__17668\
        );

    \I__4218\ : SRMux
    port map (
            O => \N__17823\,
            I => \N__17668\
        );

    \I__4217\ : SRMux
    port map (
            O => \N__17822\,
            I => \N__17668\
        );

    \I__4216\ : SRMux
    port map (
            O => \N__17821\,
            I => \N__17668\
        );

    \I__4215\ : SRMux
    port map (
            O => \N__17820\,
            I => \N__17668\
        );

    \I__4214\ : SRMux
    port map (
            O => \N__17819\,
            I => \N__17668\
        );

    \I__4213\ : SRMux
    port map (
            O => \N__17818\,
            I => \N__17668\
        );

    \I__4212\ : SRMux
    port map (
            O => \N__17817\,
            I => \N__17668\
        );

    \I__4211\ : SRMux
    port map (
            O => \N__17816\,
            I => \N__17668\
        );

    \I__4210\ : SRMux
    port map (
            O => \N__17815\,
            I => \N__17668\
        );

    \I__4209\ : SRMux
    port map (
            O => \N__17814\,
            I => \N__17668\
        );

    \I__4208\ : SRMux
    port map (
            O => \N__17813\,
            I => \N__17668\
        );

    \I__4207\ : SRMux
    port map (
            O => \N__17812\,
            I => \N__17668\
        );

    \I__4206\ : SRMux
    port map (
            O => \N__17811\,
            I => \N__17668\
        );

    \I__4205\ : SRMux
    port map (
            O => \N__17810\,
            I => \N__17668\
        );

    \I__4204\ : SRMux
    port map (
            O => \N__17809\,
            I => \N__17668\
        );

    \I__4203\ : SRMux
    port map (
            O => \N__17808\,
            I => \N__17668\
        );

    \I__4202\ : SRMux
    port map (
            O => \N__17807\,
            I => \N__17668\
        );

    \I__4201\ : SRMux
    port map (
            O => \N__17806\,
            I => \N__17668\
        );

    \I__4200\ : SRMux
    port map (
            O => \N__17805\,
            I => \N__17668\
        );

    \I__4199\ : Glb2LocalMux
    port map (
            O => \N__17802\,
            I => \N__17668\
        );

    \I__4198\ : Glb2LocalMux
    port map (
            O => \N__17799\,
            I => \N__17668\
        );

    \I__4197\ : Glb2LocalMux
    port map (
            O => \N__17796\,
            I => \N__17668\
        );

    \I__4196\ : Glb2LocalMux
    port map (
            O => \N__17793\,
            I => \N__17668\
        );

    \I__4195\ : SRMux
    port map (
            O => \N__17792\,
            I => \N__17668\
        );

    \I__4194\ : SRMux
    port map (
            O => \N__17791\,
            I => \N__17668\
        );

    \I__4193\ : SRMux
    port map (
            O => \N__17790\,
            I => \N__17668\
        );

    \I__4192\ : SRMux
    port map (
            O => \N__17789\,
            I => \N__17668\
        );

    \I__4191\ : SRMux
    port map (
            O => \N__17788\,
            I => \N__17668\
        );

    \I__4190\ : SRMux
    port map (
            O => \N__17787\,
            I => \N__17668\
        );

    \I__4189\ : SRMux
    port map (
            O => \N__17786\,
            I => \N__17668\
        );

    \I__4188\ : SRMux
    port map (
            O => \N__17785\,
            I => \N__17668\
        );

    \I__4187\ : SRMux
    port map (
            O => \N__17784\,
            I => \N__17668\
        );

    \I__4186\ : SRMux
    port map (
            O => \N__17783\,
            I => \N__17668\
        );

    \I__4185\ : SRMux
    port map (
            O => \N__17782\,
            I => \N__17668\
        );

    \I__4184\ : SRMux
    port map (
            O => \N__17781\,
            I => \N__17668\
        );

    \I__4183\ : SRMux
    port map (
            O => \N__17780\,
            I => \N__17668\
        );

    \I__4182\ : SRMux
    port map (
            O => \N__17779\,
            I => \N__17668\
        );

    \I__4181\ : SRMux
    port map (
            O => \N__17778\,
            I => \N__17668\
        );

    \I__4180\ : SRMux
    port map (
            O => \N__17777\,
            I => \N__17668\
        );

    \I__4179\ : SRMux
    port map (
            O => \N__17776\,
            I => \N__17668\
        );

    \I__4178\ : Glb2LocalMux
    port map (
            O => \N__17773\,
            I => \N__17668\
        );

    \I__4177\ : GlobalMux
    port map (
            O => \N__17668\,
            I => \N__17665\
        );

    \I__4176\ : gio2CtrlBuf
    port map (
            O => \N__17665\,
            I => rst_g
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__17662\,
            I => \Lab_UT.alarmchar_2_1_1_cascade_\
        );

    \I__4174\ : InMux
    port map (
            O => \N__17659\,
            I => \N__17656\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__17656\,
            I => \N__17653\
        );

    \I__4172\ : Odrv4
    port map (
            O => \N__17653\,
            I => \Lab_UT.alarmcharZ0Z_6\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \Lab_UT.dictrl.next_alarmstate_1_cascade_\
        );

    \I__4170\ : IoInMux
    port map (
            O => \N__17647\,
            I => \N__17639\
        );

    \I__4169\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17632\
        );

    \I__4168\ : InMux
    port map (
            O => \N__17645\,
            I => \N__17632\
        );

    \I__4167\ : InMux
    port map (
            O => \N__17644\,
            I => \N__17625\
        );

    \I__4166\ : InMux
    port map (
            O => \N__17643\,
            I => \N__17625\
        );

    \I__4165\ : InMux
    port map (
            O => \N__17642\,
            I => \N__17625\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__17639\,
            I => \N__17622\
        );

    \I__4163\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17617\
        );

    \I__4162\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17617\
        );

    \I__4161\ : LocalMux
    port map (
            O => \N__17632\,
            I => \N__17614\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17611\
        );

    \I__4159\ : Span4Mux_s3_h
    port map (
            O => \N__17622\,
            I => \N__17608\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__17617\,
            I => \N__17603\
        );

    \I__4157\ : Span12Mux_s4_h
    port map (
            O => \N__17614\,
            I => \N__17603\
        );

    \I__4156\ : Span4Mux_v
    port map (
            O => \N__17611\,
            I => \N__17598\
        );

    \I__4155\ : Span4Mux_h
    port map (
            O => \N__17608\,
            I => \N__17598\
        );

    \I__4154\ : Odrv12
    port map (
            O => \N__17603\,
            I => rst
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__17598\,
            I => rst
        );

    \I__4152\ : CascadeMux
    port map (
            O => \N__17593\,
            I => \Lab_UT.G_3_cascade_\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__17590\,
            I => \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\
        );

    \I__4150\ : InMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__17584\,
            I => \Lab_UT.dictrl.next_alarmstateZ0Z_0\
        );

    \I__4148\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17572\
        );

    \I__4147\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17572\
        );

    \I__4146\ : InMux
    port map (
            O => \N__17579\,
            I => \N__17572\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__17569\,
            I => \Lab_UT.alarmMatch\
        );

    \I__4143\ : InMux
    port map (
            O => \N__17566\,
            I => \N__17563\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__17563\,
            I => \Lab_UT.dictrl.idle\
        );

    \I__4141\ : CascadeMux
    port map (
            O => \N__17560\,
            I => \N__17555\
        );

    \I__4140\ : InMux
    port map (
            O => \N__17559\,
            I => \N__17552\
        );

    \I__4139\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17539\
        );

    \I__4138\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17536\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__17552\,
            I => \N__17533\
        );

    \I__4136\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17528\
        );

    \I__4135\ : InMux
    port map (
            O => \N__17550\,
            I => \N__17528\
        );

    \I__4134\ : InMux
    port map (
            O => \N__17549\,
            I => \N__17523\
        );

    \I__4133\ : InMux
    port map (
            O => \N__17548\,
            I => \N__17523\
        );

    \I__4132\ : InMux
    port map (
            O => \N__17547\,
            I => \N__17520\
        );

    \I__4131\ : InMux
    port map (
            O => \N__17546\,
            I => \N__17509\
        );

    \I__4130\ : InMux
    port map (
            O => \N__17545\,
            I => \N__17509\
        );

    \I__4129\ : InMux
    port map (
            O => \N__17544\,
            I => \N__17509\
        );

    \I__4128\ : InMux
    port map (
            O => \N__17543\,
            I => \N__17509\
        );

    \I__4127\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17509\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__17539\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__17536\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4124\ : Odrv4
    port map (
            O => \N__17533\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__17528\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__17523\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__17520\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__17509\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__17494\,
            I => \N__17489\
        );

    \I__4118\ : InMux
    port map (
            O => \N__17493\,
            I => \N__17483\
        );

    \I__4117\ : InMux
    port map (
            O => \N__17492\,
            I => \N__17480\
        );

    \I__4116\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17475\
        );

    \I__4115\ : InMux
    port map (
            O => \N__17488\,
            I => \N__17475\
        );

    \I__4114\ : InMux
    port map (
            O => \N__17487\,
            I => \N__17466\
        );

    \I__4113\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17466\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__17483\,
            I => \N__17463\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__17480\,
            I => \N__17460\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__17475\,
            I => \N__17457\
        );

    \I__4109\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17454\
        );

    \I__4108\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17447\
        );

    \I__4107\ : InMux
    port map (
            O => \N__17472\,
            I => \N__17447\
        );

    \I__4106\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17444\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__17466\,
            I => \N__17441\
        );

    \I__4104\ : Span4Mux_h
    port map (
            O => \N__17463\,
            I => \N__17434\
        );

    \I__4103\ : Span4Mux_v
    port map (
            O => \N__17460\,
            I => \N__17434\
        );

    \I__4102\ : Span4Mux_h
    port map (
            O => \N__17457\,
            I => \N__17434\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17431\
        );

    \I__4100\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17426\
        );

    \I__4099\ : InMux
    port map (
            O => \N__17452\,
            I => \N__17426\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__17447\,
            I => \N__17421\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17444\,
            I => \N__17421\
        );

    \I__4096\ : Span4Mux_h
    port map (
            O => \N__17441\,
            I => \N__17416\
        );

    \I__4095\ : Span4Mux_v
    port map (
            O => \N__17434\,
            I => \N__17416\
        );

    \I__4094\ : Span4Mux_h
    port map (
            O => \N__17431\,
            I => \N__17409\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__17426\,
            I => \N__17409\
        );

    \I__4092\ : Span4Mux_h
    port map (
            O => \N__17421\,
            I => \N__17409\
        );

    \I__4091\ : Odrv4
    port map (
            O => \N__17416\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__4090\ : Odrv4
    port map (
            O => \N__17409\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__4089\ : InMux
    port map (
            O => \N__17404\,
            I => \N__17401\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__4087\ : Odrv12
    port map (
            O => \N__17398\,
            I => \Lab_UT.bcd2segment4.G_64_a0Z0Z_1\
        );

    \I__4086\ : InMux
    port map (
            O => \N__17395\,
            I => \N__17392\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__17392\,
            I => \N__17389\
        );

    \I__4084\ : Span4Mux_h
    port map (
            O => \N__17389\,
            I => \N__17382\
        );

    \I__4083\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17377\
        );

    \I__4082\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17377\
        );

    \I__4081\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17372\
        );

    \I__4080\ : InMux
    port map (
            O => \N__17385\,
            I => \N__17372\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__17382\,
            I => bu_rx_data_0
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17377\,
            I => bu_rx_data_0
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__17372\,
            I => bu_rx_data_0
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__4075\ : InMux
    port map (
            O => \N__17364\,
            I => \N__17356\
        );

    \I__4074\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17351\
        );

    \I__4073\ : InMux
    port map (
            O => \N__17362\,
            I => \N__17351\
        );

    \I__4072\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17348\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__17356\,
            I => \Lab_UT.LdMtens\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__17351\,
            I => \Lab_UT.LdMtens\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__17348\,
            I => \Lab_UT.LdMtens\
        );

    \I__4068\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17337\
        );

    \I__4067\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17332\
        );

    \I__4066\ : InMux
    port map (
            O => \N__17337\,
            I => \N__17329\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__17336\,
            I => \N__17326\
        );

    \I__4064\ : InMux
    port map (
            O => \N__17335\,
            I => \N__17323\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__17332\,
            I => \N__17320\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__17329\,
            I => \N__17317\
        );

    \I__4061\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17314\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__17323\,
            I => \N__17311\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__17320\,
            I => \N__17308\
        );

    \I__4058\ : Span4Mux_v
    port map (
            O => \N__17317\,
            I => \N__17303\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17303\
        );

    \I__4056\ : Odrv12
    port map (
            O => \N__17311\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__17308\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__17303\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__4053\ : CascadeMux
    port map (
            O => \N__17296\,
            I => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_\
        );

    \I__4052\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17289\
        );

    \I__4051\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17286\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17282\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__17286\,
            I => \N__17279\
        );

    \I__4048\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17276\
        );

    \I__4047\ : Span4Mux_v
    port map (
            O => \N__17282\,
            I => \N__17272\
        );

    \I__4046\ : Span4Mux_v
    port map (
            O => \N__17279\,
            I => \N__17269\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__17276\,
            I => \N__17266\
        );

    \I__4044\ : InMux
    port map (
            O => \N__17275\,
            I => \N__17263\
        );

    \I__4043\ : Odrv4
    port map (
            O => \N__17272\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__4042\ : Odrv4
    port map (
            O => \N__17269\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__17266\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__17263\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__4039\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17243\
        );

    \I__4038\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17243\
        );

    \I__4037\ : InMux
    port map (
            O => \N__17252\,
            I => \N__17240\
        );

    \I__4036\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17231\
        );

    \I__4035\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17231\
        );

    \I__4034\ : InMux
    port map (
            O => \N__17249\,
            I => \N__17231\
        );

    \I__4033\ : InMux
    port map (
            O => \N__17248\,
            I => \N__17231\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__17243\,
            I => \N__17227\
        );

    \I__4031\ : LocalMux
    port map (
            O => \N__17240\,
            I => \N__17222\
        );

    \I__4030\ : LocalMux
    port map (
            O => \N__17231\,
            I => \N__17222\
        );

    \I__4029\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17216\
        );

    \I__4028\ : Span4Mux_v
    port map (
            O => \N__17227\,
            I => \N__17209\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__17222\,
            I => \N__17209\
        );

    \I__4026\ : InMux
    port map (
            O => \N__17221\,
            I => \N__17204\
        );

    \I__4025\ : InMux
    port map (
            O => \N__17220\,
            I => \N__17204\
        );

    \I__4024\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17198\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__17216\,
            I => \N__17195\
        );

    \I__4022\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17190\
        );

    \I__4021\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17190\
        );

    \I__4020\ : Span4Mux_h
    port map (
            O => \N__17209\,
            I => \N__17187\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__17204\,
            I => \N__17184\
        );

    \I__4018\ : InMux
    port map (
            O => \N__17203\,
            I => \N__17177\
        );

    \I__4017\ : InMux
    port map (
            O => \N__17202\,
            I => \N__17177\
        );

    \I__4016\ : InMux
    port map (
            O => \N__17201\,
            I => \N__17177\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__17198\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4014\ : Odrv12
    port map (
            O => \N__17195\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__17190\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__17187\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4011\ : Odrv12
    port map (
            O => \N__17184\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4010\ : LocalMux
    port map (
            O => \N__17177\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4009\ : InMux
    port map (
            O => \N__17164\,
            I => \N__17159\
        );

    \I__4008\ : InMux
    port map (
            O => \N__17163\,
            I => \N__17156\
        );

    \I__4007\ : InMux
    port map (
            O => \N__17162\,
            I => \N__17153\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__17159\,
            I => \Lab_UT.dictrl.dicRun_2\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__17156\,
            I => \Lab_UT.dictrl.dicRun_2\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__17153\,
            I => \Lab_UT.dictrl.dicRun_2\
        );

    \I__4003\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17134\
        );

    \I__4002\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17134\
        );

    \I__4001\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17134\
        );

    \I__4000\ : InMux
    port map (
            O => \N__17143\,
            I => \N__17134\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__17134\,
            I => \N__17131\
        );

    \I__3998\ : Odrv4
    port map (
            O => \N__17131\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__3997\ : SRMux
    port map (
            O => \N__17128\,
            I => \N__17123\
        );

    \I__3996\ : SRMux
    port map (
            O => \N__17127\,
            I => \N__17120\
        );

    \I__3995\ : SRMux
    port map (
            O => \N__17126\,
            I => \N__17117\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__17123\,
            I => \N__17114\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__17120\,
            I => \N__17111\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__17117\,
            I => \N__17108\
        );

    \I__3991\ : Span4Mux_h
    port map (
            O => \N__17114\,
            I => \N__17105\
        );

    \I__3990\ : Span4Mux_h
    port map (
            O => \N__17111\,
            I => \N__17102\
        );

    \I__3989\ : Span4Mux_h
    port map (
            O => \N__17108\,
            I => \N__17099\
        );

    \I__3988\ : Span4Mux_h
    port map (
            O => \N__17105\,
            I => \N__17096\
        );

    \I__3987\ : Span4Mux_h
    port map (
            O => \N__17102\,
            I => \N__17093\
        );

    \I__3986\ : Span4Mux_h
    port map (
            O => \N__17099\,
            I => \N__17090\
        );

    \I__3985\ : Span4Mux_v
    port map (
            O => \N__17096\,
            I => \N__17087\
        );

    \I__3984\ : Odrv4
    port map (
            O => \N__17093\,
            I => \oneSecStrb_i\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__17090\,
            I => \oneSecStrb_i\
        );

    \I__3982\ : Odrv4
    port map (
            O => \N__17087\,
            I => \oneSecStrb_i\
        );

    \I__3981\ : InMux
    port map (
            O => \N__17080\,
            I => \N__17075\
        );

    \I__3980\ : InMux
    port map (
            O => \N__17079\,
            I => \N__17068\
        );

    \I__3979\ : InMux
    port map (
            O => \N__17078\,
            I => \N__17065\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17062\
        );

    \I__3977\ : InMux
    port map (
            O => \N__17074\,
            I => \N__17053\
        );

    \I__3976\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17053\
        );

    \I__3975\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17053\
        );

    \I__3974\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17053\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__17068\,
            I => \Lab_UT.state_1\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__17065\,
            I => \Lab_UT.state_1\
        );

    \I__3971\ : Odrv12
    port map (
            O => \N__17062\,
            I => \Lab_UT.state_1\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__17053\,
            I => \Lab_UT.state_1\
        );

    \I__3969\ : InMux
    port map (
            O => \N__17044\,
            I => \N__17038\
        );

    \I__3968\ : InMux
    port map (
            O => \N__17043\,
            I => \N__17035\
        );

    \I__3967\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17032\
        );

    \I__3966\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17029\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__17038\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_2\
        );

    \I__3964\ : LocalMux
    port map (
            O => \N__17035\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_2\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__17032\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_2\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__17029\,
            I => \Lab_UT.dictrl.state_i_3Z0Z_2\
        );

    \I__3961\ : InMux
    port map (
            O => \N__17020\,
            I => \N__17010\
        );

    \I__3960\ : InMux
    port map (
            O => \N__17019\,
            I => \N__17010\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__17018\,
            I => \N__17005\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__17017\,
            I => \N__17001\
        );

    \I__3957\ : InMux
    port map (
            O => \N__17016\,
            I => \N__16996\
        );

    \I__3956\ : InMux
    port map (
            O => \N__17015\,
            I => \N__16996\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__17010\,
            I => \N__16993\
        );

    \I__3954\ : InMux
    port map (
            O => \N__17009\,
            I => \N__16984\
        );

    \I__3953\ : InMux
    port map (
            O => \N__17008\,
            I => \N__16984\
        );

    \I__3952\ : InMux
    port map (
            O => \N__17005\,
            I => \N__16984\
        );

    \I__3951\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16984\
        );

    \I__3950\ : InMux
    port map (
            O => \N__17001\,
            I => \N__16981\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__16996\,
            I => \N__16974\
        );

    \I__3948\ : Span4Mux_s3_v
    port map (
            O => \N__16993\,
            I => \N__16974\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__16984\,
            I => \N__16974\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__16981\,
            I => \N__16971\
        );

    \I__3945\ : Span4Mux_v
    port map (
            O => \N__16974\,
            I => \N__16968\
        );

    \I__3944\ : Odrv12
    port map (
            O => \N__16971\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3943\ : Odrv4
    port map (
            O => \N__16968\,
            I => \Lab_UT.state_i_3_3\
        );

    \I__3942\ : InMux
    port map (
            O => \N__16963\,
            I => \N__16958\
        );

    \I__3941\ : InMux
    port map (
            O => \N__16962\,
            I => \N__16953\
        );

    \I__3940\ : InMux
    port map (
            O => \N__16961\,
            I => \N__16953\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__16958\,
            I => \N__16950\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__16953\,
            I => \N__16947\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__16950\,
            I => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\
        );

    \I__3936\ : Odrv4
    port map (
            O => \N__16947\,
            I => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\
        );

    \I__3935\ : InMux
    port map (
            O => \N__16942\,
            I => \N__16933\
        );

    \I__3934\ : InMux
    port map (
            O => \N__16941\,
            I => \N__16933\
        );

    \I__3933\ : InMux
    port map (
            O => \N__16940\,
            I => \N__16933\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__16933\,
            I => \N__16929\
        );

    \I__3931\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16926\
        );

    \I__3930\ : Span4Mux_h
    port map (
            O => \N__16929\,
            I => \N__16923\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__16926\,
            I => \Lab_UT.dictrl.state_ret_3_RNIDH8UZ0\
        );

    \I__3928\ : Odrv4
    port map (
            O => \N__16923\,
            I => \Lab_UT.dictrl.state_ret_3_RNIDH8UZ0\
        );

    \I__3927\ : CascadeMux
    port map (
            O => \N__16918\,
            I => \N__16915\
        );

    \I__3926\ : InMux
    port map (
            O => \N__16915\,
            I => \N__16908\
        );

    \I__3925\ : InMux
    port map (
            O => \N__16914\,
            I => \N__16905\
        );

    \I__3924\ : CascadeMux
    port map (
            O => \N__16913\,
            I => \N__16902\
        );

    \I__3923\ : CascadeMux
    port map (
            O => \N__16912\,
            I => \N__16898\
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__16911\,
            I => \N__16893\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__16908\,
            I => \N__16888\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__16905\,
            I => \N__16888\
        );

    \I__3919\ : InMux
    port map (
            O => \N__16902\,
            I => \N__16881\
        );

    \I__3918\ : InMux
    port map (
            O => \N__16901\,
            I => \N__16881\
        );

    \I__3917\ : InMux
    port map (
            O => \N__16898\,
            I => \N__16874\
        );

    \I__3916\ : InMux
    port map (
            O => \N__16897\,
            I => \N__16874\
        );

    \I__3915\ : InMux
    port map (
            O => \N__16896\,
            I => \N__16874\
        );

    \I__3914\ : InMux
    port map (
            O => \N__16893\,
            I => \N__16871\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__16888\,
            I => \N__16868\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__16887\,
            I => \N__16864\
        );

    \I__3911\ : InMux
    port map (
            O => \N__16886\,
            I => \N__16860\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__16881\,
            I => \N__16855\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__16874\,
            I => \N__16855\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__16871\,
            I => \N__16852\
        );

    \I__3907\ : Span4Mux_s2_v
    port map (
            O => \N__16868\,
            I => \N__16849\
        );

    \I__3906\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16844\
        );

    \I__3905\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16844\
        );

    \I__3904\ : InMux
    port map (
            O => \N__16863\,
            I => \N__16841\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__16860\,
            I => \N__16838\
        );

    \I__3902\ : Span4Mux_v
    port map (
            O => \N__16855\,
            I => \N__16835\
        );

    \I__3901\ : Sp12to4
    port map (
            O => \N__16852\,
            I => \N__16826\
        );

    \I__3900\ : Sp12to4
    port map (
            O => \N__16849\,
            I => \N__16826\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__16844\,
            I => \N__16826\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__16841\,
            I => \N__16826\
        );

    \I__3897\ : Span4Mux_v
    port map (
            O => \N__16838\,
            I => \N__16823\
        );

    \I__3896\ : Span4Mux_v
    port map (
            O => \N__16835\,
            I => \N__16820\
        );

    \I__3895\ : Span12Mux_s10_v
    port map (
            O => \N__16826\,
            I => \N__16817\
        );

    \I__3894\ : Odrv4
    port map (
            O => \N__16823\,
            I => \Lab_UT.dictrl.state_retZ0Z_4\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__16820\,
            I => \Lab_UT.dictrl.state_retZ0Z_4\
        );

    \I__3892\ : Odrv12
    port map (
            O => \N__16817\,
            I => \Lab_UT.dictrl.state_retZ0Z_4\
        );

    \I__3891\ : InMux
    port map (
            O => \N__16810\,
            I => \N__16807\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__16807\,
            I => \N__16802\
        );

    \I__3889\ : InMux
    port map (
            O => \N__16806\,
            I => \N__16797\
        );

    \I__3888\ : InMux
    port map (
            O => \N__16805\,
            I => \N__16797\
        );

    \I__3887\ : Span4Mux_v
    port map (
            O => \N__16802\,
            I => \N__16794\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__16797\,
            I => \N__16791\
        );

    \I__3885\ : Odrv4
    port map (
            O => \N__16794\,
            I => \Lab_UT.dictrl.next_state_set\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__16791\,
            I => \Lab_UT.dictrl.next_state_set\
        );

    \I__3883\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16773\
        );

    \I__3882\ : InMux
    port map (
            O => \N__16785\,
            I => \N__16773\
        );

    \I__3881\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16773\
        );

    \I__3880\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16769\
        );

    \I__3879\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16762\
        );

    \I__3878\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16762\
        );

    \I__3877\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16762\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__16773\,
            I => \N__16756\
        );

    \I__3875\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16752\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__16769\,
            I => \N__16747\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__16762\,
            I => \N__16747\
        );

    \I__3872\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16740\
        );

    \I__3871\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16740\
        );

    \I__3870\ : InMux
    port map (
            O => \N__16759\,
            I => \N__16740\
        );

    \I__3869\ : Span4Mux_h
    port map (
            O => \N__16756\,
            I => \N__16737\
        );

    \I__3868\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16734\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__16752\,
            I => \Lab_UT.state_0\
        );

    \I__3866\ : Odrv4
    port map (
            O => \N__16747\,
            I => \Lab_UT.state_0\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__16740\,
            I => \Lab_UT.state_0\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__16737\,
            I => \Lab_UT.state_0\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__16734\,
            I => \Lab_UT.state_0\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__3861\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__16717\,
            I => \N__16714\
        );

    \I__3859\ : Odrv4
    port map (
            O => \N__16714\,
            I => \Lab_UT.alarmcharZ0Z_4\
        );

    \I__3858\ : InMux
    port map (
            O => \N__16711\,
            I => \N__16705\
        );

    \I__3857\ : InMux
    port map (
            O => \N__16710\,
            I => \N__16705\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__16705\,
            I => \Lab_UT.N_204\
        );

    \I__3855\ : CascadeMux
    port map (
            O => \N__16702\,
            I => \Lab_UT.N_204_cascade_\
        );

    \I__3854\ : InMux
    port map (
            O => \N__16699\,
            I => \N__16687\
        );

    \I__3853\ : InMux
    port map (
            O => \N__16698\,
            I => \N__16687\
        );

    \I__3852\ : InMux
    port map (
            O => \N__16697\,
            I => \N__16687\
        );

    \I__3851\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16687\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__16687\,
            I => \N__16684\
        );

    \I__3849\ : Odrv4
    port map (
            O => \N__16684\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__3848\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16675\
        );

    \I__3847\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16675\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__16675\,
            I => \Lab_UT.nine\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__16672\,
            I => \N__16668\
        );

    \I__3844\ : CascadeMux
    port map (
            O => \N__16671\,
            I => \N__16664\
        );

    \I__3843\ : InMux
    port map (
            O => \N__16668\,
            I => \N__16658\
        );

    \I__3842\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16658\
        );

    \I__3841\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16653\
        );

    \I__3840\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16653\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__16658\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__16653\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__16648\,
            I => \N__16640\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__16647\,
            I => \N__16637\
        );

    \I__3835\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16633\
        );

    \I__3834\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16626\
        );

    \I__3833\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16626\
        );

    \I__3832\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16626\
        );

    \I__3831\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16619\
        );

    \I__3830\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16619\
        );

    \I__3829\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16619\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16614\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__16626\,
            I => \N__16606\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__16619\,
            I => \N__16606\
        );

    \I__3825\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16603\
        );

    \I__3824\ : InMux
    port map (
            O => \N__16617\,
            I => \N__16600\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__16614\,
            I => \N__16597\
        );

    \I__3822\ : InMux
    port map (
            O => \N__16613\,
            I => \N__16590\
        );

    \I__3821\ : InMux
    port map (
            O => \N__16612\,
            I => \N__16590\
        );

    \I__3820\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16590\
        );

    \I__3819\ : Span4Mux_v
    port map (
            O => \N__16606\,
            I => \N__16587\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__16603\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__16600\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3816\ : Odrv4
    port map (
            O => \N__16597\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__16590\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3814\ : Odrv4
    port map (
            O => \N__16587\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3813\ : InMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__3812\ : InMux
    port map (
            O => \N__16575\,
            I => \N__16559\
        );

    \I__3811\ : InMux
    port map (
            O => \N__16574\,
            I => \N__16559\
        );

    \I__3810\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16559\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__16570\,
            I => \N__16555\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__16569\,
            I => \N__16550\
        );

    \I__3807\ : InMux
    port map (
            O => \N__16568\,
            I => \N__16541\
        );

    \I__3806\ : InMux
    port map (
            O => \N__16567\,
            I => \N__16541\
        );

    \I__3805\ : InMux
    port map (
            O => \N__16566\,
            I => \N__16541\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__16559\,
            I => \N__16538\
        );

    \I__3803\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16535\
        );

    \I__3802\ : Span4Mux_s3_h
    port map (
            O => \N__16555\,
            I => \N__16532\
        );

    \I__3801\ : InMux
    port map (
            O => \N__16554\,
            I => \N__16527\
        );

    \I__3800\ : InMux
    port map (
            O => \N__16553\,
            I => \N__16527\
        );

    \I__3799\ : InMux
    port map (
            O => \N__16550\,
            I => \N__16520\
        );

    \I__3798\ : InMux
    port map (
            O => \N__16549\,
            I => \N__16520\
        );

    \I__3797\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16520\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__16541\,
            I => \N__16515\
        );

    \I__3795\ : Span12Mux_s9_v
    port map (
            O => \N__16538\,
            I => \N__16515\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__16535\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__16532\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__16527\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__16520\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3790\ : Odrv12
    port map (
            O => \N__16515\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__3789\ : CascadeMux
    port map (
            O => \N__16504\,
            I => \N__16496\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__16503\,
            I => \N__16493\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__16502\,
            I => \N__16490\
        );

    \I__3786\ : InMux
    port map (
            O => \N__16501\,
            I => \N__16483\
        );

    \I__3785\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16483\
        );

    \I__3784\ : InMux
    port map (
            O => \N__16499\,
            I => \N__16483\
        );

    \I__3783\ : InMux
    port map (
            O => \N__16496\,
            I => \N__16474\
        );

    \I__3782\ : InMux
    port map (
            O => \N__16493\,
            I => \N__16474\
        );

    \I__3781\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16474\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16471\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__16482\,
            I => \N__16468\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16481\,
            I => \N__16462\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__16474\,
            I => \N__16454\
        );

    \I__3776\ : Span4Mux_v
    port map (
            O => \N__16471\,
            I => \N__16454\
        );

    \I__3775\ : InMux
    port map (
            O => \N__16468\,
            I => \N__16451\
        );

    \I__3774\ : InMux
    port map (
            O => \N__16467\,
            I => \N__16444\
        );

    \I__3773\ : InMux
    port map (
            O => \N__16466\,
            I => \N__16444\
        );

    \I__3772\ : InMux
    port map (
            O => \N__16465\,
            I => \N__16444\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__16462\,
            I => \N__16441\
        );

    \I__3770\ : InMux
    port map (
            O => \N__16461\,
            I => \N__16434\
        );

    \I__3769\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16434\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16434\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__16454\,
            I => \N__16431\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__16451\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__16444\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3764\ : Odrv12
    port map (
            O => \N__16441\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__16434\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3762\ : Odrv4
    port map (
            O => \N__16431\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__16420\,
            I => \N__16414\
        );

    \I__3760\ : InMux
    port map (
            O => \N__16419\,
            I => \N__16411\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16399\
        );

    \I__3758\ : InMux
    port map (
            O => \N__16417\,
            I => \N__16399\
        );

    \I__3757\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16399\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16394\
        );

    \I__3755\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16387\
        );

    \I__3754\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16387\
        );

    \I__3753\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16387\
        );

    \I__3752\ : CascadeMux
    port map (
            O => \N__16407\,
            I => \N__16384\
        );

    \I__3751\ : CascadeMux
    port map (
            O => \N__16406\,
            I => \N__16381\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__16399\,
            I => \N__16378\
        );

    \I__3749\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16375\
        );

    \I__3748\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16372\
        );

    \I__3747\ : Span12Mux_s9_v
    port map (
            O => \N__16394\,
            I => \N__16367\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__16387\,
            I => \N__16367\
        );

    \I__3745\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16362\
        );

    \I__3744\ : InMux
    port map (
            O => \N__16381\,
            I => \N__16362\
        );

    \I__3743\ : Span4Mux_h
    port map (
            O => \N__16378\,
            I => \N__16359\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__16375\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__16372\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3740\ : Odrv12
    port map (
            O => \N__16367\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16362\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__16359\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3737\ : InMux
    port map (
            O => \N__16348\,
            I => \N__16345\
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__16345\,
            I => \N__16342\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__16342\,
            I => \N__16336\
        );

    \I__3734\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16333\
        );

    \I__3733\ : InMux
    port map (
            O => \N__16340\,
            I => \N__16328\
        );

    \I__3732\ : InMux
    port map (
            O => \N__16339\,
            I => \N__16328\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__16336\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__16333\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__16328\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__3728\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16314\
        );

    \I__3727\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__3726\ : CascadeMux
    port map (
            O => \N__16319\,
            I => \N__16305\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__16314\,
            I => \N__16302\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16313\,
            I => \N__16297\
        );

    \I__3723\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16297\
        );

    \I__3722\ : CascadeMux
    port map (
            O => \N__16311\,
            I => \N__16293\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__16310\,
            I => \N__16288\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16285\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16280\
        );

    \I__3718\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16280\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__16302\,
            I => \N__16275\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__16297\,
            I => \N__16275\
        );

    \I__3715\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16262\
        );

    \I__3714\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16262\
        );

    \I__3713\ : InMux
    port map (
            O => \N__16292\,
            I => \N__16262\
        );

    \I__3712\ : InMux
    port map (
            O => \N__16291\,
            I => \N__16262\
        );

    \I__3711\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16262\
        );

    \I__3710\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16262\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__16280\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__16275\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__16262\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__16255\,
            I => \N__16252\
        );

    \I__3705\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16247\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__16251\,
            I => \N__16244\
        );

    \I__3703\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16240\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__16247\,
            I => \N__16236\
        );

    \I__3701\ : InMux
    port map (
            O => \N__16244\,
            I => \N__16231\
        );

    \I__3700\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16231\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16226\
        );

    \I__3698\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16217\
        );

    \I__3697\ : Span4Mux_v
    port map (
            O => \N__16236\,
            I => \N__16212\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__16231\,
            I => \N__16212\
        );

    \I__3695\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16207\
        );

    \I__3694\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16207\
        );

    \I__3693\ : Span4Mux_s3_h
    port map (
            O => \N__16226\,
            I => \N__16204\
        );

    \I__3692\ : InMux
    port map (
            O => \N__16225\,
            I => \N__16191\
        );

    \I__3691\ : InMux
    port map (
            O => \N__16224\,
            I => \N__16191\
        );

    \I__3690\ : InMux
    port map (
            O => \N__16223\,
            I => \N__16191\
        );

    \I__3689\ : InMux
    port map (
            O => \N__16222\,
            I => \N__16191\
        );

    \I__3688\ : InMux
    port map (
            O => \N__16221\,
            I => \N__16191\
        );

    \I__3687\ : InMux
    port map (
            O => \N__16220\,
            I => \N__16191\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__16217\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__3685\ : Odrv4
    port map (
            O => \N__16212\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__16207\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__16204\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__16191\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__3681\ : InMux
    port map (
            O => \N__16180\,
            I => \N__16177\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__16177\,
            I => \Lab_UT.didp.countrce2.three_2\
        );

    \I__3679\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16168\
        );

    \I__3678\ : CascadeMux
    port map (
            O => \N__16173\,
            I => \N__16165\
        );

    \I__3677\ : CascadeMux
    port map (
            O => \N__16172\,
            I => \N__16157\
        );

    \I__3676\ : InMux
    port map (
            O => \N__16171\,
            I => \N__16152\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__16168\,
            I => \N__16149\
        );

    \I__3674\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16146\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__16164\,
            I => \N__16142\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__16163\,
            I => \N__16139\
        );

    \I__3671\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16134\
        );

    \I__3670\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16131\
        );

    \I__3669\ : InMux
    port map (
            O => \N__16160\,
            I => \N__16126\
        );

    \I__3668\ : InMux
    port map (
            O => \N__16157\,
            I => \N__16126\
        );

    \I__3667\ : InMux
    port map (
            O => \N__16156\,
            I => \N__16121\
        );

    \I__3666\ : InMux
    port map (
            O => \N__16155\,
            I => \N__16121\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__16152\,
            I => \N__16114\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__16149\,
            I => \N__16114\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__16146\,
            I => \N__16114\
        );

    \I__3662\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16103\
        );

    \I__3661\ : InMux
    port map (
            O => \N__16142\,
            I => \N__16103\
        );

    \I__3660\ : InMux
    port map (
            O => \N__16139\,
            I => \N__16103\
        );

    \I__3659\ : InMux
    port map (
            O => \N__16138\,
            I => \N__16103\
        );

    \I__3658\ : InMux
    port map (
            O => \N__16137\,
            I => \N__16103\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__16134\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__16131\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__16126\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__16121\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__16114\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__16103\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__3651\ : CascadeMux
    port map (
            O => \N__16090\,
            I => \Lab_UT.didp.countrce2.three_2_cascade_\
        );

    \I__3650\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__16084\,
            I => \Lab_UT.didp.countrce2.un20_qPone\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__16080\,
            I => \N__16072\
        );

    \I__3646\ : InMux
    port map (
            O => \N__16079\,
            I => \N__16064\
        );

    \I__3645\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16064\
        );

    \I__3644\ : InMux
    port map (
            O => \N__16075\,
            I => \N__16059\
        );

    \I__3643\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16059\
        );

    \I__3642\ : CascadeMux
    port map (
            O => \N__16071\,
            I => \N__16056\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__16070\,
            I => \N__16053\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__16069\,
            I => \N__16050\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__16064\,
            I => \N__16044\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__16059\,
            I => \N__16041\
        );

    \I__3637\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16032\
        );

    \I__3636\ : InMux
    port map (
            O => \N__16053\,
            I => \N__16032\
        );

    \I__3635\ : InMux
    port map (
            O => \N__16050\,
            I => \N__16032\
        );

    \I__3634\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16032\
        );

    \I__3633\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16028\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__16047\,
            I => \N__16022\
        );

    \I__3631\ : Span4Mux_v
    port map (
            O => \N__16044\,
            I => \N__16015\
        );

    \I__3630\ : Span4Mux_h
    port map (
            O => \N__16041\,
            I => \N__16015\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__16032\,
            I => \N__16015\
        );

    \I__3628\ : InMux
    port map (
            O => \N__16031\,
            I => \N__16012\
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__16028\,
            I => \N__16009\
        );

    \I__3626\ : InMux
    port map (
            O => \N__16027\,
            I => \N__16006\
        );

    \I__3625\ : InMux
    port map (
            O => \N__16026\,
            I => \N__15999\
        );

    \I__3624\ : InMux
    port map (
            O => \N__16025\,
            I => \N__15999\
        );

    \I__3623\ : InMux
    port map (
            O => \N__16022\,
            I => \N__15999\
        );

    \I__3622\ : Span4Mux_h
    port map (
            O => \N__16015\,
            I => \N__15996\
        );

    \I__3621\ : LocalMux
    port map (
            O => \N__16012\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3620\ : Odrv4
    port map (
            O => \N__16009\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__16006\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__15999\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3617\ : Odrv4
    port map (
            O => \N__15996\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__15985\,
            I => \N__15974\
        );

    \I__3615\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15969\
        );

    \I__3614\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15969\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15982\,
            I => \N__15963\
        );

    \I__3612\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15963\
        );

    \I__3611\ : InMux
    port map (
            O => \N__15980\,
            I => \N__15954\
        );

    \I__3610\ : InMux
    port map (
            O => \N__15979\,
            I => \N__15954\
        );

    \I__3609\ : InMux
    port map (
            O => \N__15978\,
            I => \N__15954\
        );

    \I__3608\ : InMux
    port map (
            O => \N__15977\,
            I => \N__15954\
        );

    \I__3607\ : InMux
    port map (
            O => \N__15974\,
            I => \N__15950\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__15969\,
            I => \N__15947\
        );

    \I__3605\ : InMux
    port map (
            O => \N__15968\,
            I => \N__15940\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__15963\,
            I => \N__15937\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__15954\,
            I => \N__15934\
        );

    \I__3602\ : InMux
    port map (
            O => \N__15953\,
            I => \N__15931\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__15950\,
            I => \N__15928\
        );

    \I__3600\ : Span4Mux_v
    port map (
            O => \N__15947\,
            I => \N__15925\
        );

    \I__3599\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15916\
        );

    \I__3598\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15916\
        );

    \I__3597\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15916\
        );

    \I__3596\ : InMux
    port map (
            O => \N__15943\,
            I => \N__15916\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__15940\,
            I => \N__15909\
        );

    \I__3594\ : Span4Mux_h
    port map (
            O => \N__15937\,
            I => \N__15909\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__15934\,
            I => \N__15909\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__15931\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__15928\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__15925\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__15916\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__15909\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__3587\ : InMux
    port map (
            O => \N__15898\,
            I => \N__15895\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__15895\,
            I => \N__15891\
        );

    \I__3585\ : InMux
    port map (
            O => \N__15894\,
            I => \N__15888\
        );

    \I__3584\ : Span4Mux_h
    port map (
            O => \N__15891\,
            I => \N__15885\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__15888\,
            I => \Lab_UT.N_207\
        );

    \I__3582\ : Odrv4
    port map (
            O => \N__15885\,
            I => \Lab_UT.N_207\
        );

    \I__3581\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \N__15876\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15879\,
            I => \N__15872\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15876\,
            I => \N__15867\
        );

    \I__3578\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15867\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__15872\,
            I => \N__15864\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__15867\,
            I => \Lab_UT.didp.q_RNI84NN1_3\
        );

    \I__3575\ : Odrv4
    port map (
            O => \N__15864\,
            I => \Lab_UT.didp.q_RNI84NN1_3\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__15859\,
            I => \N__15856\
        );

    \I__3573\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15852\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__15855\,
            I => \N__15848\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15852\,
            I => \N__15844\
        );

    \I__3570\ : InMux
    port map (
            O => \N__15851\,
            I => \N__15837\
        );

    \I__3569\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15837\
        );

    \I__3568\ : InMux
    port map (
            O => \N__15847\,
            I => \N__15837\
        );

    \I__3567\ : Odrv4
    port map (
            O => \N__15844\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__15837\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__3565\ : InMux
    port map (
            O => \N__15832\,
            I => \N__15829\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__15829\,
            I => \N__15826\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__15826\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_3\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__15823\,
            I => \N__15815\
        );

    \I__3561\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15808\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15808\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15820\,
            I => \N__15803\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15819\,
            I => \N__15803\
        );

    \I__3557\ : InMux
    port map (
            O => \N__15818\,
            I => \N__15796\
        );

    \I__3556\ : InMux
    port map (
            O => \N__15815\,
            I => \N__15796\
        );

    \I__3555\ : InMux
    port map (
            O => \N__15814\,
            I => \N__15796\
        );

    \I__3554\ : InMux
    port map (
            O => \N__15813\,
            I => \N__15791\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__15808\,
            I => \N__15788\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__15803\,
            I => \N__15785\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__15796\,
            I => \N__15782\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__15795\,
            I => \N__15779\
        );

    \I__3549\ : CascadeMux
    port map (
            O => \N__15794\,
            I => \N__15775\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__15791\,
            I => \N__15770\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__15788\,
            I => \N__15767\
        );

    \I__3546\ : Span4Mux_h
    port map (
            O => \N__15785\,
            I => \N__15762\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__15782\,
            I => \N__15762\
        );

    \I__3544\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15753\
        );

    \I__3543\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15753\
        );

    \I__3542\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15753\
        );

    \I__3541\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15753\
        );

    \I__3540\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15750\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__15770\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3538\ : Odrv4
    port map (
            O => \N__15767\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3537\ : Odrv4
    port map (
            O => \N__15762\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__15753\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__15750\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__15739\,
            I => \N__15735\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__15738\,
            I => \N__15732\
        );

    \I__3532\ : InMux
    port map (
            O => \N__15735\,
            I => \N__15721\
        );

    \I__3531\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15721\
        );

    \I__3530\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15716\
        );

    \I__3529\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15716\
        );

    \I__3528\ : InMux
    port map (
            O => \N__15729\,
            I => \N__15709\
        );

    \I__3527\ : InMux
    port map (
            O => \N__15728\,
            I => \N__15709\
        );

    \I__3526\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15709\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15706\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__15721\,
            I => \N__15703\
        );

    \I__3523\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15693\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__15709\,
            I => \N__15693\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__15706\,
            I => \N__15689\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__15703\,
            I => \N__15686\
        );

    \I__3519\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15675\
        );

    \I__3518\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15675\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15675\
        );

    \I__3516\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15675\
        );

    \I__3515\ : InMux
    port map (
            O => \N__15698\,
            I => \N__15675\
        );

    \I__3514\ : Span4Mux_h
    port map (
            O => \N__15693\,
            I => \N__15672\
        );

    \I__3513\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15669\
        );

    \I__3512\ : Odrv4
    port map (
            O => \N__15689\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__15686\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__15675\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__15672\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__15669\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__15658\,
            I => \Lab_UT.N_207_cascade_\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__15655\,
            I => \N__15652\
        );

    \I__3505\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__3504\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15646\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__15646\,
            I => \N__15643\
        );

    \I__3502\ : Odrv4
    port map (
            O => \N__15643\,
            I => \Lab_UT.didp.q_RNIIKFH3_3\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__15640\,
            I => \N__15635\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15639\,
            I => \N__15632\
        );

    \I__3499\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15629\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15635\,
            I => \N__15626\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__15632\,
            I => \N__15623\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__15629\,
            I => \N__15619\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__15626\,
            I => \N__15614\
        );

    \I__3494\ : Span4Mux_h
    port map (
            O => \N__15623\,
            I => \N__15614\
        );

    \I__3493\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15611\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__15619\,
            I => \Lab_UT.m40\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__15614\,
            I => \Lab_UT.m40\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15611\,
            I => \Lab_UT.m40\
        );

    \I__3489\ : CascadeMux
    port map (
            O => \N__15604\,
            I => \N__15601\
        );

    \I__3488\ : InMux
    port map (
            O => \N__15601\,
            I => \N__15597\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__15600\,
            I => \N__15594\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__15597\,
            I => \N__15590\
        );

    \I__3485\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15587\
        );

    \I__3484\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15584\
        );

    \I__3483\ : Span4Mux_h
    port map (
            O => \N__15590\,
            I => \N__15581\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__15587\,
            I => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__15584\,
            I => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3\
        );

    \I__3480\ : Odrv4
    port map (
            O => \N__15581\,
            I => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3\
        );

    \I__3479\ : InMux
    port map (
            O => \N__15574\,
            I => \N__15571\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__15571\,
            I => \N__15566\
        );

    \I__3477\ : InMux
    port map (
            O => \N__15570\,
            I => \N__15562\
        );

    \I__3476\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15559\
        );

    \I__3475\ : Span4Mux_h
    port map (
            O => \N__15566\,
            I => \N__15556\
        );

    \I__3474\ : InMux
    port map (
            O => \N__15565\,
            I => \N__15553\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__15562\,
            I => \N__15548\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__15559\,
            I => \N__15548\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__15556\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__15553\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__15548\,
            I => \Lab_UT.dictrl.next_state_set_2\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15541\,
            I => \N__15538\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__15538\,
            I => \N__15535\
        );

    \I__3466\ : Odrv4
    port map (
            O => \N__15535\,
            I => \Lab_UT.alarmcharZ0Z_2\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__15532\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_2_cascade_\
        );

    \I__3464\ : CascadeMux
    port map (
            O => \N__15529\,
            I => \N__15522\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15519\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__15527\,
            I => \N__15516\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__15526\,
            I => \N__15513\
        );

    \I__3460\ : InMux
    port map (
            O => \N__15525\,
            I => \N__15508\
        );

    \I__3459\ : InMux
    port map (
            O => \N__15522\,
            I => \N__15503\
        );

    \I__3458\ : InMux
    port map (
            O => \N__15519\,
            I => \N__15503\
        );

    \I__3457\ : InMux
    port map (
            O => \N__15516\,
            I => \N__15498\
        );

    \I__3456\ : InMux
    port map (
            O => \N__15513\,
            I => \N__15498\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15495\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__15511\,
            I => \N__15491\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__15508\,
            I => \N__15483\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__15503\,
            I => \N__15480\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__15498\,
            I => \N__15477\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15474\
        );

    \I__3449\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15469\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15469\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__15490\,
            I => \N__15466\
        );

    \I__3446\ : InMux
    port map (
            O => \N__15489\,
            I => \N__15461\
        );

    \I__3445\ : InMux
    port map (
            O => \N__15488\,
            I => \N__15461\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__15487\,
            I => \N__15458\
        );

    \I__3443\ : InMux
    port map (
            O => \N__15486\,
            I => \N__15455\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__15483\,
            I => \N__15450\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__15480\,
            I => \N__15450\
        );

    \I__3440\ : Span4Mux_v
    port map (
            O => \N__15477\,
            I => \N__15443\
        );

    \I__3439\ : Span4Mux_v
    port map (
            O => \N__15474\,
            I => \N__15443\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__15469\,
            I => \N__15443\
        );

    \I__3437\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15440\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__15461\,
            I => \N__15437\
        );

    \I__3435\ : InMux
    port map (
            O => \N__15458\,
            I => \N__15434\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__15455\,
            I => \N__15429\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__15450\,
            I => \N__15429\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__15443\,
            I => \N__15426\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__15440\,
            I => \N__15423\
        );

    \I__3430\ : Odrv12
    port map (
            O => \N__15437\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__15434\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__15429\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__15426\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3426\ : Odrv12
    port map (
            O => \N__15423\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__3425\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__15409\,
            I => \N__15406\
        );

    \I__3423\ : Odrv12
    port map (
            O => \N__15406\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_2\
        );

    \I__3422\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15394\
        );

    \I__3421\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15394\
        );

    \I__3420\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15394\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__15394\,
            I => \N__15390\
        );

    \I__3418\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__3417\ : Odrv4
    port map (
            O => \N__15390\,
            I => \Lab_UT.un3_dOutP\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__15387\,
            I => \Lab_UT.un3_dOutP\
        );

    \I__3415\ : InMux
    port map (
            O => \N__15382\,
            I => \N__15378\
        );

    \I__3414\ : InMux
    port map (
            O => \N__15381\,
            I => \N__15368\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15365\
        );

    \I__3412\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15362\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__15376\,
            I => \N__15359\
        );

    \I__3410\ : InMux
    port map (
            O => \N__15375\,
            I => \N__15348\
        );

    \I__3409\ : InMux
    port map (
            O => \N__15374\,
            I => \N__15348\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15373\,
            I => \N__15348\
        );

    \I__3407\ : InMux
    port map (
            O => \N__15372\,
            I => \N__15348\
        );

    \I__3406\ : InMux
    port map (
            O => \N__15371\,
            I => \N__15348\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__15368\,
            I => \N__15341\
        );

    \I__3404\ : Span4Mux_h
    port map (
            O => \N__15365\,
            I => \N__15341\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__15362\,
            I => \N__15341\
        );

    \I__3402\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15336\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__15348\,
            I => \N__15333\
        );

    \I__3400\ : Span4Mux_v
    port map (
            O => \N__15341\,
            I => \N__15330\
        );

    \I__3399\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15325\
        );

    \I__3398\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15325\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__15336\,
            I => \Lab_UT.cnt_3\
        );

    \I__3396\ : Odrv12
    port map (
            O => \N__15333\,
            I => \Lab_UT.cnt_3\
        );

    \I__3395\ : Odrv4
    port map (
            O => \N__15330\,
            I => \Lab_UT.cnt_3\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__15325\,
            I => \Lab_UT.cnt_3\
        );

    \I__3393\ : InMux
    port map (
            O => \N__15316\,
            I => \N__15313\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__15313\,
            I => \N__15308\
        );

    \I__3391\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15303\
        );

    \I__3390\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15303\
        );

    \I__3389\ : Span4Mux_v
    port map (
            O => \N__15308\,
            I => \N__15300\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__15303\,
            I => \N__15297\
        );

    \I__3387\ : Sp12to4
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__15297\,
            I => \N__15291\
        );

    \I__3385\ : Span12Mux_s6_h
    port map (
            O => \N__15294\,
            I => \N__15286\
        );

    \I__3384\ : Span4Mux_h
    port map (
            O => \N__15291\,
            I => \N__15283\
        );

    \I__3383\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15278\
        );

    \I__3382\ : InMux
    port map (
            O => \N__15289\,
            I => \N__15278\
        );

    \I__3381\ : Odrv12
    port map (
            O => \N__15286\,
            I => \Lab_UT.cnt_0\
        );

    \I__3380\ : Odrv4
    port map (
            O => \N__15283\,
            I => \Lab_UT.cnt_0\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__15278\,
            I => \Lab_UT.cnt_0\
        );

    \I__3378\ : InMux
    port map (
            O => \N__15271\,
            I => \N__15262\
        );

    \I__3377\ : InMux
    port map (
            O => \N__15270\,
            I => \N__15251\
        );

    \I__3376\ : InMux
    port map (
            O => \N__15269\,
            I => \N__15251\
        );

    \I__3375\ : InMux
    port map (
            O => \N__15268\,
            I => \N__15251\
        );

    \I__3374\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15251\
        );

    \I__3373\ : InMux
    port map (
            O => \N__15266\,
            I => \N__15251\
        );

    \I__3372\ : InMux
    port map (
            O => \N__15265\,
            I => \N__15248\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__15262\,
            I => \N__15236\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__15251\,
            I => \N__15236\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__15248\,
            I => \N__15233\
        );

    \I__3368\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15224\
        );

    \I__3367\ : InMux
    port map (
            O => \N__15246\,
            I => \N__15224\
        );

    \I__3366\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15224\
        );

    \I__3365\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15224\
        );

    \I__3364\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15221\
        );

    \I__3363\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15218\
        );

    \I__3362\ : InMux
    port map (
            O => \N__15241\,
            I => \N__15215\
        );

    \I__3361\ : Span4Mux_h
    port map (
            O => \N__15236\,
            I => \N__15212\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__15233\,
            I => \N__15207\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__15224\,
            I => \N__15207\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__15221\,
            I => \N__15199\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__15218\,
            I => \N__15199\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__15215\,
            I => \N__15199\
        );

    \I__3355\ : Span4Mux_v
    port map (
            O => \N__15212\,
            I => \N__15194\
        );

    \I__3354\ : Span4Mux_h
    port map (
            O => \N__15207\,
            I => \N__15194\
        );

    \I__3353\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15191\
        );

    \I__3352\ : Span12Mux_s11_h
    port map (
            O => \N__15199\,
            I => \N__15188\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__15194\,
            I => \N__15185\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__15191\,
            I => \Lab_UT.cnt_1\
        );

    \I__3349\ : Odrv12
    port map (
            O => \N__15188\,
            I => \Lab_UT.cnt_1\
        );

    \I__3348\ : Odrv4
    port map (
            O => \N__15185\,
            I => \Lab_UT.cnt_1\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__15178\,
            I => \N__15175\
        );

    \I__3346\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15167\
        );

    \I__3345\ : InMux
    port map (
            O => \N__15174\,
            I => \N__15164\
        );

    \I__3344\ : CascadeMux
    port map (
            O => \N__15173\,
            I => \N__15159\
        );

    \I__3343\ : CascadeMux
    port map (
            O => \N__15172\,
            I => \N__15156\
        );

    \I__3342\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15152\
        );

    \I__3341\ : InMux
    port map (
            O => \N__15170\,
            I => \N__15149\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15142\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__15164\,
            I => \N__15142\
        );

    \I__3338\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15131\
        );

    \I__3337\ : InMux
    port map (
            O => \N__15162\,
            I => \N__15131\
        );

    \I__3336\ : InMux
    port map (
            O => \N__15159\,
            I => \N__15131\
        );

    \I__3335\ : InMux
    port map (
            O => \N__15156\,
            I => \N__15131\
        );

    \I__3334\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15131\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__15152\,
            I => \N__15126\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__15149\,
            I => \N__15126\
        );

    \I__3331\ : CascadeMux
    port map (
            O => \N__15148\,
            I => \N__15123\
        );

    \I__3330\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15117\
        );

    \I__3329\ : Sp12to4
    port map (
            O => \N__15142\,
            I => \N__15112\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__15131\,
            I => \N__15112\
        );

    \I__3327\ : Span4Mux_h
    port map (
            O => \N__15126\,
            I => \N__15109\
        );

    \I__3326\ : InMux
    port map (
            O => \N__15123\,
            I => \N__15100\
        );

    \I__3325\ : InMux
    port map (
            O => \N__15122\,
            I => \N__15100\
        );

    \I__3324\ : InMux
    port map (
            O => \N__15121\,
            I => \N__15100\
        );

    \I__3323\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15100\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__15117\,
            I => \Lab_UT.cnt_2\
        );

    \I__3321\ : Odrv12
    port map (
            O => \N__15112\,
            I => \Lab_UT.cnt_2\
        );

    \I__3320\ : Odrv4
    port map (
            O => \N__15109\,
            I => \Lab_UT.cnt_2\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__15100\,
            I => \Lab_UT.cnt_2\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__15091\,
            I => \Lab_UT.alarmchar9_cascade_\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__15088\,
            I => \N__15084\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__15087\,
            I => \N__15081\
        );

    \I__3315\ : InMux
    port map (
            O => \N__15084\,
            I => \N__15076\
        );

    \I__3314\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15076\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__15076\,
            I => \Lab_UT.alarmcharZ0Z_1\
        );

    \I__3312\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15070\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__15070\,
            I => \N__15067\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__15067\,
            I => \Lab_UT.zero\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__15064\,
            I => \Lab_UT.didp.countrce3.qPone_3_cascade_\
        );

    \I__3308\ : CascadeMux
    port map (
            O => \N__15061\,
            I => \Lab_UT.didp.countrce3.N_79_i_cascade_\
        );

    \I__3307\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15052\
        );

    \I__3306\ : InMux
    port map (
            O => \N__15057\,
            I => \N__15045\
        );

    \I__3305\ : InMux
    port map (
            O => \N__15056\,
            I => \N__15045\
        );

    \I__3304\ : InMux
    port map (
            O => \N__15055\,
            I => \N__15045\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__15052\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__15045\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__15040\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_0_cascade_\
        );

    \I__3300\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__15034\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_0\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__15031\,
            I => \N__15025\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__15030\,
            I => \N__15022\
        );

    \I__3296\ : InMux
    port map (
            O => \N__15029\,
            I => \N__15019\
        );

    \I__3295\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15016\
        );

    \I__3294\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15011\
        );

    \I__3293\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15011\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__15019\,
            I => \Lab_UT.un29_dOutP\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__15016\,
            I => \Lab_UT.un29_dOutP\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__15011\,
            I => \Lab_UT.un29_dOutP\
        );

    \I__3289\ : InMux
    port map (
            O => \N__15004\,
            I => \N__15001\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__15001\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_1\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__14998\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_1_cascade_\
        );

    \I__3286\ : InMux
    port map (
            O => \N__14995\,
            I => \N__14992\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__14992\,
            I => \N__14988\
        );

    \I__3284\ : InMux
    port map (
            O => \N__14991\,
            I => \N__14984\
        );

    \I__3283\ : Span4Mux_h
    port map (
            O => \N__14988\,
            I => \N__14981\
        );

    \I__3282\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14978\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14973\
        );

    \I__3280\ : Span4Mux_h
    port map (
            O => \N__14981\,
            I => \N__14970\
        );

    \I__3279\ : LocalMux
    port map (
            O => \N__14978\,
            I => \N__14967\
        );

    \I__3278\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14962\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14962\
        );

    \I__3276\ : Odrv12
    port map (
            O => \N__14973\,
            I => \L3_tx_data_1\
        );

    \I__3275\ : Odrv4
    port map (
            O => \N__14970\,
            I => \L3_tx_data_1\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__14967\,
            I => \L3_tx_data_1\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__14962\,
            I => \L3_tx_data_1\
        );

    \I__3272\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14950\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__14950\,
            I => \N__14947\
        );

    \I__3270\ : Odrv4
    port map (
            O => \N__14947\,
            I => \Lab_UT.dispString.dOutP_0_iv_3_1\
        );

    \I__3269\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14938\
        );

    \I__3268\ : InMux
    port map (
            O => \N__14943\,
            I => \N__14932\
        );

    \I__3267\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14929\
        );

    \I__3266\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14926\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__14938\,
            I => \N__14923\
        );

    \I__3264\ : InMux
    port map (
            O => \N__14937\,
            I => \N__14920\
        );

    \I__3263\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14909\
        );

    \I__3262\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14909\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__14932\,
            I => \N__14906\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__14929\,
            I => \N__14903\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__14926\,
            I => \N__14896\
        );

    \I__3258\ : Span4Mux_v
    port map (
            O => \N__14923\,
            I => \N__14896\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__14920\,
            I => \N__14896\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14919\,
            I => \N__14893\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14888\
        );

    \I__3254\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14888\
        );

    \I__3253\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14883\
        );

    \I__3252\ : InMux
    port map (
            O => \N__14915\,
            I => \N__14883\
        );

    \I__3251\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14879\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__14909\,
            I => \N__14874\
        );

    \I__3249\ : Span4Mux_v
    port map (
            O => \N__14906\,
            I => \N__14874\
        );

    \I__3248\ : Span4Mux_s3_h
    port map (
            O => \N__14903\,
            I => \N__14867\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__14896\,
            I => \N__14867\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__14893\,
            I => \N__14867\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__14888\,
            I => \N__14862\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14883\,
            I => \N__14862\
        );

    \I__3243\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14859\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__14879\,
            I => \N__14852\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__14874\,
            I => \N__14852\
        );

    \I__3240\ : Span4Mux_v
    port map (
            O => \N__14867\,
            I => \N__14852\
        );

    \I__3239\ : Odrv4
    port map (
            O => \N__14862\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__14859\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3237\ : Odrv4
    port map (
            O => \N__14852\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__3236\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14842\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__14842\,
            I => \Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0\
        );

    \I__3234\ : InMux
    port map (
            O => \N__14839\,
            I => \N__14835\
        );

    \I__3233\ : InMux
    port map (
            O => \N__14838\,
            I => \N__14832\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__14835\,
            I => \N__14826\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__14832\,
            I => \N__14826\
        );

    \I__3230\ : InMux
    port map (
            O => \N__14831\,
            I => \N__14823\
        );

    \I__3229\ : Span4Mux_h
    port map (
            O => \N__14826\,
            I => \N__14820\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__14823\,
            I => \Lab_UT.m24\
        );

    \I__3227\ : Odrv4
    port map (
            O => \N__14820\,
            I => \Lab_UT.m24\
        );

    \I__3226\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14809\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14809\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__14809\,
            I => \Lab_UT.dispString.un22_dOutP\
        );

    \I__3223\ : InMux
    port map (
            O => \N__14806\,
            I => \N__14803\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__14803\,
            I => \N__14800\
        );

    \I__3221\ : Odrv4
    port map (
            O => \N__14800\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_3\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__14797\,
            I => \Lab_UT.dispString.dOutP_0_iv_3_3_cascade_\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14794\,
            I => \N__14791\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__14791\,
            I => \N__14787\
        );

    \I__3217\ : InMux
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__14787\,
            I => \N__14781\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__14784\,
            I => \N__14778\
        );

    \I__3214\ : Span4Mux_h
    port map (
            O => \N__14781\,
            I => \N__14774\
        );

    \I__3213\ : Span12Mux_s8_h
    port map (
            O => \N__14778\,
            I => \N__14771\
        );

    \I__3212\ : InMux
    port map (
            O => \N__14777\,
            I => \N__14768\
        );

    \I__3211\ : Odrv4
    port map (
            O => \N__14774\,
            I => \L3_tx_data_3\
        );

    \I__3210\ : Odrv12
    port map (
            O => \N__14771\,
            I => \L3_tx_data_3\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__14768\,
            I => \L3_tx_data_3\
        );

    \I__3208\ : InMux
    port map (
            O => \N__14761\,
            I => \N__14758\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__14758\,
            I => \Lab_UT.alarmcharZ0Z_0\
        );

    \I__3206\ : SRMux
    port map (
            O => \N__14755\,
            I => \N__14752\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__14752\,
            I => \N__14748\
        );

    \I__3204\ : InMux
    port map (
            O => \N__14751\,
            I => \N__14745\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__14745\,
            I => \N__14739\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__14742\,
            I => \Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1\
        );

    \I__3200\ : Odrv12
    port map (
            O => \N__14739\,
            I => \Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14734\,
            I => \N__14728\
        );

    \I__3198\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14728\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__14728\,
            I => \N__14725\
        );

    \I__3196\ : Span4Mux_h
    port map (
            O => \N__14725\,
            I => \N__14722\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__14722\,
            I => \N__14718\
        );

    \I__3194\ : InMux
    port map (
            O => \N__14721\,
            I => \N__14715\
        );

    \I__3193\ : Odrv4
    port map (
            O => \N__14718\,
            I => \L3_tx_data_5\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__14715\,
            I => \L3_tx_data_5\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__14710\,
            I => \Lab_UT.dispString.dOutP_0_iv_3_2_cascade_\
        );

    \I__3190\ : InMux
    port map (
            O => \N__14707\,
            I => \N__14701\
        );

    \I__3189\ : InMux
    port map (
            O => \N__14706\,
            I => \N__14701\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__14701\,
            I => \N__14696\
        );

    \I__3187\ : InMux
    port map (
            O => \N__14700\,
            I => \N__14691\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14691\
        );

    \I__3185\ : Odrv12
    port map (
            O => \N__14696\,
            I => \L3_tx_data_2\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__14691\,
            I => \L3_tx_data_2\
        );

    \I__3183\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14680\
        );

    \I__3182\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14680\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__14680\,
            I => \N__14677\
        );

    \I__3180\ : Span4Mux_v
    port map (
            O => \N__14677\,
            I => \N__14673\
        );

    \I__3179\ : CascadeMux
    port map (
            O => \N__14676\,
            I => \N__14670\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__14673\,
            I => \N__14667\
        );

    \I__3177\ : InMux
    port map (
            O => \N__14670\,
            I => \N__14664\
        );

    \I__3176\ : Odrv4
    port map (
            O => \N__14667\,
            I => \L3_tx_data_6\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__14664\,
            I => \L3_tx_data_6\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__14656\,
            I => \N__14652\
        );

    \I__3172\ : InMux
    port map (
            O => \N__14655\,
            I => \N__14649\
        );

    \I__3171\ : Odrv12
    port map (
            O => \N__14652\,
            I => \L3_tx_data_4\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__14649\,
            I => \L3_tx_data_4\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__14644\,
            I => \Lab_UT.dictrl.un1_state_12_cascade_\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14641\,
            I => \N__14638\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14638\,
            I => \Lab_UT.didp.m37_nsZ0Z_1\
        );

    \I__3166\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__14632\,
            I => \N__14624\
        );

    \I__3164\ : InMux
    port map (
            O => \N__14631\,
            I => \N__14619\
        );

    \I__3163\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14619\
        );

    \I__3162\ : InMux
    port map (
            O => \N__14629\,
            I => \N__14612\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14612\
        );

    \I__3160\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14612\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__14624\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__14619\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__14612\,
            I => \Lab_UT.state_i_3_1\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__14605\,
            I => \N__14598\
        );

    \I__3155\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14594\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__14603\,
            I => \N__14591\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__14602\,
            I => \N__14588\
        );

    \I__3152\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14584\
        );

    \I__3151\ : InMux
    port map (
            O => \N__14598\,
            I => \N__14577\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14577\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__14594\,
            I => \N__14574\
        );

    \I__3148\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14567\
        );

    \I__3147\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14567\
        );

    \I__3146\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14567\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14564\
        );

    \I__3144\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14559\
        );

    \I__3143\ : InMux
    port map (
            O => \N__14582\,
            I => \N__14559\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__14577\,
            I => \Lab_UT.state_2\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__14574\,
            I => \Lab_UT.state_2\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__14567\,
            I => \Lab_UT.state_2\
        );

    \I__3139\ : Odrv4
    port map (
            O => \N__14564\,
            I => \Lab_UT.state_2\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__14559\,
            I => \Lab_UT.state_2\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__14548\,
            I => \N__14543\
        );

    \I__3136\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14538\
        );

    \I__3135\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14533\
        );

    \I__3134\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14533\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__14542\,
            I => \N__14530\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \N__14526\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14538\,
            I => \N__14523\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14520\
        );

    \I__3129\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14517\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14514\
        );

    \I__3127\ : InMux
    port map (
            O => \N__14526\,
            I => \N__14511\
        );

    \I__3126\ : Odrv12
    port map (
            O => \N__14523\,
            I => \Lab_UT.state_3\
        );

    \I__3125\ : Odrv4
    port map (
            O => \N__14520\,
            I => \Lab_UT.state_3\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__14517\,
            I => \Lab_UT.state_3\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__14514\,
            I => \Lab_UT.state_3\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__14511\,
            I => \Lab_UT.state_3\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__14500\,
            I => \Lab_UT.dictrl.un1_state_24_ns_1_cascade_\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__14497\,
            I => \N__14493\
        );

    \I__3119\ : InMux
    port map (
            O => \N__14496\,
            I => \N__14489\
        );

    \I__3118\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14486\
        );

    \I__3117\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14483\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14489\,
            I => \N__14480\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14477\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__14483\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__14480\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__14477\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__14470\,
            I => \N__14466\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14469\,
            I => \N__14462\
        );

    \I__3109\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14457\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14457\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14454\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__14457\,
            I => \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1\
        );

    \I__3105\ : Odrv4
    port map (
            O => \N__14454\,
            I => \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1\
        );

    \I__3104\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14440\
        );

    \I__3103\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14440\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14447\,
            I => \N__14437\
        );

    \I__3101\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14434\
        );

    \I__3100\ : InMux
    port map (
            O => \N__14445\,
            I => \N__14431\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__14440\,
            I => \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__14437\,
            I => \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__14434\,
            I => \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__14431\,
            I => \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__14422\,
            I => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_\
        );

    \I__3094\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14413\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14408\
        );

    \I__3092\ : InMux
    port map (
            O => \N__14417\,
            I => \N__14408\
        );

    \I__3091\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14405\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__14413\,
            I => \N__14398\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14398\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__14405\,
            I => \N__14398\
        );

    \I__3087\ : Odrv4
    port map (
            O => \N__14398\,
            I => \Lab_UT.dictrl.next_state_set_0\
        );

    \I__3086\ : InMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__14392\,
            I => \Lab_UT.dictrl.next_state_out_1\
        );

    \I__3084\ : CEMux
    port map (
            O => \N__14389\,
            I => \N__14384\
        );

    \I__3083\ : CEMux
    port map (
            O => \N__14388\,
            I => \N__14380\
        );

    \I__3082\ : CEMux
    port map (
            O => \N__14387\,
            I => \N__14377\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__14384\,
            I => \N__14374\
        );

    \I__3080\ : CEMux
    port map (
            O => \N__14383\,
            I => \N__14371\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14380\,
            I => \N__14368\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14365\
        );

    \I__3077\ : Span4Mux_v
    port map (
            O => \N__14374\,
            I => \N__14362\
        );

    \I__3076\ : LocalMux
    port map (
            O => \N__14371\,
            I => \N__14359\
        );

    \I__3075\ : Odrv4
    port map (
            O => \N__14368\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__3074\ : Odrv4
    port map (
            O => \N__14365\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__3073\ : Odrv4
    port map (
            O => \N__14362\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__14359\,
            I => \Lab_UT.dictrl.un1_state_21_reti_i\
        );

    \I__3071\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14347\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__14347\,
            I => \Lab_UT.didp.countrce4.N_88_i\
        );

    \I__3069\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14340\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14343\,
            I => \N__14337\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__14340\,
            I => \N__14334\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__14337\,
            I => \N__14331\
        );

    \I__3065\ : Span4Mux_h
    port map (
            O => \N__14334\,
            I => \N__14328\
        );

    \I__3064\ : Odrv4
    port map (
            O => \N__14331\,
            I => \Lab_UT.N_68_0\
        );

    \I__3063\ : Odrv4
    port map (
            O => \N__14328\,
            I => \Lab_UT.N_68_0\
        );

    \I__3062\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14320\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__14320\,
            I => \N__14317\
        );

    \I__3060\ : Span4Mux_v
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__14314\,
            I => \Lab_UT.didp.un31_reset_i_a4_1\
        );

    \I__3058\ : InMux
    port map (
            O => \N__14311\,
            I => \N__14305\
        );

    \I__3057\ : InMux
    port map (
            O => \N__14310\,
            I => \N__14300\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14309\,
            I => \N__14300\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14297\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__14305\,
            I => \N__14294\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__14300\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__14297\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__3051\ : Odrv4
    port map (
            O => \N__14294\,
            I => \Lab_UT.dictrl.next_state_set_1\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__14287\,
            I => \N__14283\
        );

    \I__3049\ : InMux
    port map (
            O => \N__14286\,
            I => \N__14276\
        );

    \I__3048\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14276\
        );

    \I__3047\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14273\
        );

    \I__3046\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14270\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__14276\,
            I => \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14273\,
            I => \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__14270\,
            I => \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2\
        );

    \I__3042\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14255\
        );

    \I__3041\ : InMux
    port map (
            O => \N__14262\,
            I => \N__14255\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14261\,
            I => \N__14252\
        );

    \I__3039\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14249\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__14255\,
            I => \Lab_UT.m37_ns\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__14252\,
            I => \Lab_UT.m37_ns\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__14249\,
            I => \Lab_UT.m37_ns\
        );

    \I__3035\ : InMux
    port map (
            O => \N__14242\,
            I => \N__14218\
        );

    \I__3034\ : InMux
    port map (
            O => \N__14241\,
            I => \N__14218\
        );

    \I__3033\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14212\
        );

    \I__3032\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14204\
        );

    \I__3031\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14199\
        );

    \I__3030\ : InMux
    port map (
            O => \N__14237\,
            I => \N__14199\
        );

    \I__3029\ : InMux
    port map (
            O => \N__14236\,
            I => \N__14192\
        );

    \I__3028\ : InMux
    port map (
            O => \N__14235\,
            I => \N__14192\
        );

    \I__3027\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14192\
        );

    \I__3026\ : InMux
    port map (
            O => \N__14233\,
            I => \N__14187\
        );

    \I__3025\ : InMux
    port map (
            O => \N__14232\,
            I => \N__14187\
        );

    \I__3024\ : InMux
    port map (
            O => \N__14231\,
            I => \N__14180\
        );

    \I__3023\ : InMux
    port map (
            O => \N__14230\,
            I => \N__14180\
        );

    \I__3022\ : InMux
    port map (
            O => \N__14229\,
            I => \N__14180\
        );

    \I__3021\ : InMux
    port map (
            O => \N__14228\,
            I => \N__14173\
        );

    \I__3020\ : InMux
    port map (
            O => \N__14227\,
            I => \N__14173\
        );

    \I__3019\ : InMux
    port map (
            O => \N__14226\,
            I => \N__14173\
        );

    \I__3018\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14166\
        );

    \I__3017\ : InMux
    port map (
            O => \N__14224\,
            I => \N__14166\
        );

    \I__3016\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14166\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__14218\,
            I => \N__14163\
        );

    \I__3014\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14156\
        );

    \I__3013\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14156\
        );

    \I__3012\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14156\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__14212\,
            I => \N__14153\
        );

    \I__3010\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14146\
        );

    \I__3009\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14146\
        );

    \I__3008\ : InMux
    port map (
            O => \N__14209\,
            I => \N__14146\
        );

    \I__3007\ : InMux
    port map (
            O => \N__14208\,
            I => \N__14141\
        );

    \I__3006\ : InMux
    port map (
            O => \N__14207\,
            I => \N__14141\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14138\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__14199\,
            I => \N__14129\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__14192\,
            I => \N__14129\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__14187\,
            I => \N__14129\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__14180\,
            I => \N__14129\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__14173\,
            I => \N__14126\
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__14166\,
            I => \N__14115\
        );

    \I__2998\ : Span4Mux_h
    port map (
            O => \N__14163\,
            I => \N__14115\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__14156\,
            I => \N__14115\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__14153\,
            I => \N__14115\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__14146\,
            I => \N__14104\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14104\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__14138\,
            I => \N__14104\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__14129\,
            I => \N__14104\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__14126\,
            I => \N__14104\
        );

    \I__2990\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14099\
        );

    \I__2989\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14099\
        );

    \I__2988\ : Span4Mux_v
    port map (
            O => \N__14115\,
            I => \N__14096\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__14104\,
            I => \N__14093\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__14099\,
            I => \Lab_UT.Run\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__14096\,
            I => \Lab_UT.Run\
        );

    \I__2984\ : Odrv4
    port map (
            O => \N__14093\,
            I => \Lab_UT.Run\
        );

    \I__2983\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14082\
        );

    \I__2982\ : InMux
    port map (
            O => \N__14085\,
            I => \N__14079\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__14082\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__14079\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1\
        );

    \I__2979\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14069\
        );

    \I__2978\ : InMux
    port map (
            O => \N__14073\,
            I => \N__14064\
        );

    \I__2977\ : InMux
    port map (
            O => \N__14072\,
            I => \N__14064\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__14069\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__14064\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__14059\,
            I => \Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_\
        );

    \I__2973\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__14053\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa\
        );

    \I__2971\ : InMux
    port map (
            O => \N__14050\,
            I => \N__14047\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__2969\ : Odrv4
    port map (
            O => \N__14044\,
            I => \Lab_UT.didp.m34_nsZ0Z_1\
        );

    \I__2968\ : InMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2967\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14035\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__14035\,
            I => \N__14031\
        );

    \I__2965\ : InMux
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__2964\ : Span4Mux_h
    port map (
            O => \N__14031\,
            I => \N__14025\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__14028\,
            I => \Lab_UT.dictrl.next_state16Z0Z_4\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__14025\,
            I => \Lab_UT.dictrl.next_state16Z0Z_4\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__14020\,
            I => \Lab_UT.m34_ns_cascade_\
        );

    \I__2960\ : InMux
    port map (
            O => \N__14017\,
            I => \N__14014\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__14014\,
            I => \N__14011\
        );

    \I__2958\ : Span4Mux_s2_h
    port map (
            O => \N__14011\,
            I => \N__14008\
        );

    \I__2957\ : Span4Mux_h
    port map (
            O => \N__14008\,
            I => \N__14003\
        );

    \I__2956\ : InMux
    port map (
            O => \N__14007\,
            I => \N__14000\
        );

    \I__2955\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13997\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__14003\,
            I => \resetGen_escKey_4\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__14000\,
            I => \resetGen_escKey_4\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__13997\,
            I => \resetGen_escKey_4\
        );

    \I__2951\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13987\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__13987\,
            I => \N__13984\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__13984\,
            I => \N__13975\
        );

    \I__2948\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13970\
        );

    \I__2947\ : InMux
    port map (
            O => \N__13982\,
            I => \N__13970\
        );

    \I__2946\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13961\
        );

    \I__2945\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13961\
        );

    \I__2944\ : InMux
    port map (
            O => \N__13979\,
            I => \N__13961\
        );

    \I__2943\ : InMux
    port map (
            O => \N__13978\,
            I => \N__13961\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__13975\,
            I => bu_rx_data_1
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__13970\,
            I => bu_rx_data_1
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__13961\,
            I => bu_rx_data_1
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__13954\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13951\,
            I => \N__13948\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__13948\,
            I => \N__13943\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__13947\,
            I => \N__13940\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__13946\,
            I => \N__13934\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__13943\,
            I => \N__13931\
        );

    \I__2933\ : InMux
    port map (
            O => \N__13940\,
            I => \N__13920\
        );

    \I__2932\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13920\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13938\,
            I => \N__13920\
        );

    \I__2930\ : InMux
    port map (
            O => \N__13937\,
            I => \N__13920\
        );

    \I__2929\ : InMux
    port map (
            O => \N__13934\,
            I => \N__13920\
        );

    \I__2928\ : Span4Mux_h
    port map (
            O => \N__13931\,
            I => \N__13917\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__13920\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__13917\,
            I => \resetGen.reset_countZ0Z_4\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13909\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13909\,
            I => \Lab_UT.dictrl.next_state_out_3\
        );

    \I__2923\ : SRMux
    port map (
            O => \N__13906\,
            I => \N__13903\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__13903\,
            I => \N__13900\
        );

    \I__2921\ : Odrv12
    port map (
            O => \N__13900\,
            I => \Lab_UT.m34_ns\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__13897\,
            I => \Lab_UT.didp.N_164_cascade_\
        );

    \I__2919\ : SRMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__2917\ : Span4Mux_v
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__2916\ : Span4Mux_h
    port map (
            O => \N__13885\,
            I => \N__13881\
        );

    \I__2915\ : InMux
    port map (
            O => \N__13884\,
            I => \N__13878\
        );

    \I__2914\ : Odrv4
    port map (
            O => \N__13881\,
            I => \Lab_UT.m42\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13878\,
            I => \Lab_UT.m42\
        );

    \I__2912\ : InMux
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__13870\,
            I => \Lab_UT.bcd2segment2.segment_i_0Z0Z_1\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__13867\,
            I => \Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_\
        );

    \I__2909\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13861\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__2907\ : Odrv4
    port map (
            O => \N__13858\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__13855\,
            I => \Lab_UT.three_2_cascade_\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__13849\,
            I => \Lab_UT.didp.countrce1.un20_qPone\
        );

    \I__2903\ : InMux
    port map (
            O => \N__13846\,
            I => \N__13843\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__13843\,
            I => \uu2.mem0.g0_7_4_0\
        );

    \I__2901\ : CascadeMux
    port map (
            O => \N__13840\,
            I => \N__13835\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__13839\,
            I => \N__13832\
        );

    \I__2899\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13825\
        );

    \I__2898\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13817\
        );

    \I__2897\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13817\
        );

    \I__2896\ : InMux
    port map (
            O => \N__13831\,
            I => \N__13817\
        );

    \I__2895\ : InMux
    port map (
            O => \N__13830\,
            I => \N__13814\
        );

    \I__2894\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13811\
        );

    \I__2893\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13808\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__13825\,
            I => \N__13805\
        );

    \I__2891\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13797\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__13817\,
            I => \N__13792\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__13814\,
            I => \N__13792\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__13811\,
            I => \N__13789\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__13808\,
            I => \N__13786\
        );

    \I__2886\ : Span4Mux_h
    port map (
            O => \N__13805\,
            I => \N__13783\
        );

    \I__2885\ : InMux
    port map (
            O => \N__13804\,
            I => \N__13780\
        );

    \I__2884\ : InMux
    port map (
            O => \N__13803\,
            I => \N__13771\
        );

    \I__2883\ : InMux
    port map (
            O => \N__13802\,
            I => \N__13771\
        );

    \I__2882\ : InMux
    port map (
            O => \N__13801\,
            I => \N__13771\
        );

    \I__2881\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13771\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__13797\,
            I => \N__13764\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__13792\,
            I => \N__13764\
        );

    \I__2878\ : Span4Mux_h
    port map (
            O => \N__13789\,
            I => \N__13764\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__13786\,
            I => \uu2.N_46\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__13783\,
            I => \uu2.N_46\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__13780\,
            I => \uu2.N_46\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__13771\,
            I => \uu2.N_46\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__13764\,
            I => \uu2.N_46\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__13753\,
            I => \N__13748\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__13752\,
            I => \N__13743\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__13751\,
            I => \N__13740\
        );

    \I__2869\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13734\
        );

    \I__2868\ : InMux
    port map (
            O => \N__13747\,
            I => \N__13731\
        );

    \I__2867\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13728\
        );

    \I__2866\ : InMux
    port map (
            O => \N__13743\,
            I => \N__13723\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13740\,
            I => \N__13723\
        );

    \I__2864\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13720\
        );

    \I__2863\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13717\
        );

    \I__2862\ : InMux
    port map (
            O => \N__13737\,
            I => \N__13713\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__13734\,
            I => \N__13703\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__13731\,
            I => \N__13700\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__13728\,
            I => \N__13693\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__13723\,
            I => \N__13693\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__13720\,
            I => \N__13693\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__13717\,
            I => \N__13690\
        );

    \I__2855\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13687\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__13713\,
            I => \N__13684\
        );

    \I__2853\ : InMux
    port map (
            O => \N__13712\,
            I => \N__13671\
        );

    \I__2852\ : InMux
    port map (
            O => \N__13711\,
            I => \N__13671\
        );

    \I__2851\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13671\
        );

    \I__2850\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13671\
        );

    \I__2849\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13664\
        );

    \I__2848\ : InMux
    port map (
            O => \N__13707\,
            I => \N__13664\
        );

    \I__2847\ : InMux
    port map (
            O => \N__13706\,
            I => \N__13664\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__13703\,
            I => \N__13655\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__13700\,
            I => \N__13655\
        );

    \I__2844\ : Span4Mux_v
    port map (
            O => \N__13693\,
            I => \N__13655\
        );

    \I__2843\ : Span4Mux_v
    port map (
            O => \N__13690\,
            I => \N__13655\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N__13650\
        );

    \I__2841\ : Span4Mux_h
    port map (
            O => \N__13684\,
            I => \N__13650\
        );

    \I__2840\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13641\
        );

    \I__2839\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13641\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13641\
        );

    \I__2837\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13641\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__13671\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__13664\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2834\ : Odrv4
    port map (
            O => \N__13655\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__13650\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__13641\,
            I => \uu2.w_addr_displayingZ0Z_4\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__13630\,
            I => \N__13620\
        );

    \I__2830\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13616\
        );

    \I__2829\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13613\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__13627\,
            I => \N__13610\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__13626\,
            I => \N__13606\
        );

    \I__2826\ : InMux
    port map (
            O => \N__13625\,
            I => \N__13595\
        );

    \I__2825\ : InMux
    port map (
            O => \N__13624\,
            I => \N__13595\
        );

    \I__2824\ : InMux
    port map (
            O => \N__13623\,
            I => \N__13595\
        );

    \I__2823\ : InMux
    port map (
            O => \N__13620\,
            I => \N__13595\
        );

    \I__2822\ : InMux
    port map (
            O => \N__13619\,
            I => \N__13595\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__13616\,
            I => \N__13588\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__13613\,
            I => \N__13588\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13585\
        );

    \I__2818\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13580\
        );

    \I__2817\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13580\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__13595\,
            I => \N__13574\
        );

    \I__2815\ : InMux
    port map (
            O => \N__13594\,
            I => \N__13569\
        );

    \I__2814\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13569\
        );

    \I__2813\ : Span4Mux_v
    port map (
            O => \N__13588\,
            I => \N__13564\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__13585\,
            I => \N__13564\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13561\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13579\,
            I => \N__13554\
        );

    \I__2809\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13554\
        );

    \I__2808\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13554\
        );

    \I__2807\ : Span4Mux_v
    port map (
            O => \N__13574\,
            I => \N__13551\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__13569\,
            I => \N__13546\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__13564\,
            I => \N__13546\
        );

    \I__2804\ : Span4Mux_h
    port map (
            O => \N__13561\,
            I => \N__13541\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__13554\,
            I => \N__13541\
        );

    \I__2802\ : Odrv4
    port map (
            O => \N__13551\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__13546\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2800\ : Odrv4
    port map (
            O => \N__13541\,
            I => \uu2.w_addr_displayingZ0Z_3\
        );

    \I__2799\ : CEMux
    port map (
            O => \N__13534\,
            I => \N__13530\
        );

    \I__2798\ : CEMux
    port map (
            O => \N__13533\,
            I => \N__13527\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__13530\,
            I => \N__13524\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__13527\,
            I => \N__13520\
        );

    \I__2795\ : Span4Mux_v
    port map (
            O => \N__13524\,
            I => \N__13517\
        );

    \I__2794\ : CEMux
    port map (
            O => \N__13523\,
            I => \N__13514\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__13520\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__13517\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13514\,
            I => \uu2.un21_w_addr_displaying_i_0\
        );

    \I__2790\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13495\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__13506\,
            I => \N__13491\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__13505\,
            I => \N__13488\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__13504\,
            I => \N__13485\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__13503\,
            I => \N__13482\
        );

    \I__2785\ : InMux
    port map (
            O => \N__13502\,
            I => \N__13479\
        );

    \I__2784\ : InMux
    port map (
            O => \N__13501\,
            I => \N__13476\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13500\,
            I => \N__13471\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13471\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__13498\,
            I => \N__13468\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__13495\,
            I => \N__13465\
        );

    \I__2779\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13459\
        );

    \I__2778\ : InMux
    port map (
            O => \N__13491\,
            I => \N__13459\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13452\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13485\,
            I => \N__13452\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13482\,
            I => \N__13452\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__13479\,
            I => \N__13449\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__13476\,
            I => \N__13446\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__13471\,
            I => \N__13443\
        );

    \I__2771\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13440\
        );

    \I__2770\ : Span4Mux_v
    port map (
            O => \N__13465\,
            I => \N__13437\
        );

    \I__2769\ : InMux
    port map (
            O => \N__13464\,
            I => \N__13434\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__13459\,
            I => \N__13429\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__13452\,
            I => \N__13429\
        );

    \I__2766\ : Span4Mux_h
    port map (
            O => \N__13449\,
            I => \N__13422\
        );

    \I__2765\ : Span4Mux_h
    port map (
            O => \N__13446\,
            I => \N__13422\
        );

    \I__2764\ : Span4Mux_h
    port map (
            O => \N__13443\,
            I => \N__13422\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__13440\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__13437\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__13434\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__13429\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2759\ : Odrv4
    port map (
            O => \N__13422\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__2758\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13406\
        );

    \I__2757\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13403\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__13409\,
            I => \N__13399\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__13406\,
            I => \N__13391\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__13403\,
            I => \N__13388\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__13402\,
            I => \N__13385\
        );

    \I__2752\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13377\
        );

    \I__2751\ : InMux
    port map (
            O => \N__13398\,
            I => \N__13377\
        );

    \I__2750\ : InMux
    port map (
            O => \N__13397\,
            I => \N__13377\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__13396\,
            I => \N__13370\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__13395\,
            I => \N__13367\
        );

    \I__2747\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13364\
        );

    \I__2746\ : Span4Mux_h
    port map (
            O => \N__13391\,
            I => \N__13361\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__13388\,
            I => \N__13358\
        );

    \I__2744\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13353\
        );

    \I__2743\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13353\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__13377\,
            I => \N__13350\
        );

    \I__2741\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13343\
        );

    \I__2740\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13343\
        );

    \I__2739\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13343\
        );

    \I__2738\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13340\
        );

    \I__2737\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13335\
        );

    \I__2736\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13335\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__13364\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__13361\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2733\ : Odrv4
    port map (
            O => \N__13358\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__13353\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2731\ : Odrv4
    port map (
            O => \N__13350\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13343\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__13340\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__13335\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__2727\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13313\
        );

    \I__2726\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13310\
        );

    \I__2725\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13307\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__13313\,
            I => \N__13300\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__13310\,
            I => \N__13297\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__13307\,
            I => \N__13294\
        );

    \I__2721\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13291\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__13305\,
            I => \N__13284\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__13304\,
            I => \N__13281\
        );

    \I__2718\ : InMux
    port map (
            O => \N__13303\,
            I => \N__13277\
        );

    \I__2717\ : Span4Mux_h
    port map (
            O => \N__13300\,
            I => \N__13274\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__13297\,
            I => \N__13271\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__13294\,
            I => \N__13268\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__13291\,
            I => \N__13265\
        );

    \I__2713\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13260\
        );

    \I__2712\ : InMux
    port map (
            O => \N__13289\,
            I => \N__13260\
        );

    \I__2711\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13253\
        );

    \I__2710\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13253\
        );

    \I__2709\ : InMux
    port map (
            O => \N__13284\,
            I => \N__13253\
        );

    \I__2708\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13248\
        );

    \I__2707\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13248\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__13277\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__13274\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2704\ : Odrv4
    port map (
            O => \N__13271\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__13268\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__13265\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__13260\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__13253\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__13248\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__2698\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13226\
        );

    \I__2697\ : InMux
    port map (
            O => \N__13230\,
            I => \N__13220\
        );

    \I__2696\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13220\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13217\
        );

    \I__2694\ : InMux
    port map (
            O => \N__13225\,
            I => \N__13209\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13206\
        );

    \I__2692\ : Span4Mux_h
    port map (
            O => \N__13217\,
            I => \N__13197\
        );

    \I__2691\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13194\
        );

    \I__2690\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13191\
        );

    \I__2689\ : InMux
    port map (
            O => \N__13214\,
            I => \N__13186\
        );

    \I__2688\ : InMux
    port map (
            O => \N__13213\,
            I => \N__13186\
        );

    \I__2687\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13183\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__13209\,
            I => \N__13180\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__13206\,
            I => \N__13177\
        );

    \I__2684\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13168\
        );

    \I__2683\ : InMux
    port map (
            O => \N__13204\,
            I => \N__13168\
        );

    \I__2682\ : InMux
    port map (
            O => \N__13203\,
            I => \N__13168\
        );

    \I__2681\ : InMux
    port map (
            O => \N__13202\,
            I => \N__13168\
        );

    \I__2680\ : InMux
    port map (
            O => \N__13201\,
            I => \N__13163\
        );

    \I__2679\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13163\
        );

    \I__2678\ : Span4Mux_v
    port map (
            O => \N__13197\,
            I => \N__13154\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__13194\,
            I => \N__13154\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13154\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__13186\,
            I => \N__13154\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__13183\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__13180\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__13177\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__13168\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__13163\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__13154\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__2668\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13138\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__13138\,
            I => \N__13135\
        );

    \I__2666\ : Odrv12
    port map (
            O => \N__13135\,
            I => \uu2.mem0.g0_16_1\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__13132\,
            I => \Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13126\
        );

    \I__2663\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13123\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__13123\,
            I => \N__13120\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__13120\,
            I => \N__13117\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__13117\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__13114\,
            I => \Lab_UT.nine_cascade_\
        );

    \I__2658\ : CascadeMux
    port map (
            O => \N__13111\,
            I => \N__13106\
        );

    \I__2657\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13099\
        );

    \I__2656\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13099\
        );

    \I__2655\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13099\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__13099\,
            I => \N__13096\
        );

    \I__2653\ : Span4Mux_h
    port map (
            O => \N__13096\,
            I => \N__13093\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__13093\,
            I => \uu2.N_49\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__13090\,
            I => \uu2.mem0.g0_7_5_0_cascade_\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__13087\,
            I => \uu2.mem0.un31_w_data_displaying_1_0_0_cascade_\
        );

    \I__2649\ : InMux
    port map (
            O => \N__13084\,
            I => \N__13081\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__13081\,
            I => \N__13078\
        );

    \I__2647\ : Span4Mux_v
    port map (
            O => \N__13078\,
            I => \N__13075\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__13075\,
            I => \uu2.mem0.g1_0_1\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__13072\,
            I => \N__13066\
        );

    \I__2644\ : InMux
    port map (
            O => \N__13071\,
            I => \N__13059\
        );

    \I__2643\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13056\
        );

    \I__2642\ : InMux
    port map (
            O => \N__13069\,
            I => \N__13053\
        );

    \I__2641\ : InMux
    port map (
            O => \N__13066\,
            I => \N__13043\
        );

    \I__2640\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13043\
        );

    \I__2639\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13043\
        );

    \I__2638\ : InMux
    port map (
            O => \N__13063\,
            I => \N__13038\
        );

    \I__2637\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13038\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__13059\,
            I => \N__13033\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__13056\,
            I => \N__13033\
        );

    \I__2634\ : LocalMux
    port map (
            O => \N__13053\,
            I => \N__13024\
        );

    \I__2633\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13021\
        );

    \I__2632\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13018\
        );

    \I__2631\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13015\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__13043\,
            I => \N__13008\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__13038\,
            I => \N__13008\
        );

    \I__2628\ : Span4Mux_v
    port map (
            O => \N__13033\,
            I => \N__13008\
        );

    \I__2627\ : InMux
    port map (
            O => \N__13032\,
            I => \N__13003\
        );

    \I__2626\ : InMux
    port map (
            O => \N__13031\,
            I => \N__13003\
        );

    \I__2625\ : InMux
    port map (
            O => \N__13030\,
            I => \N__12994\
        );

    \I__2624\ : InMux
    port map (
            O => \N__13029\,
            I => \N__12994\
        );

    \I__2623\ : InMux
    port map (
            O => \N__13028\,
            I => \N__12994\
        );

    \I__2622\ : InMux
    port map (
            O => \N__13027\,
            I => \N__12994\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__13024\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__13021\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__13018\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__13015\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__13008\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__13003\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__12994\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__12979\,
            I => \N__12975\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12978\,
            I => \N__12966\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12975\,
            I => \N__12959\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12959\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12973\,
            I => \N__12959\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__12972\,
            I => \N__12956\
        );

    \I__2608\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12949\
        );

    \I__2607\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12949\
        );

    \I__2606\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12942\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__12966\,
            I => \N__12937\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12959\,
            I => \N__12937\
        );

    \I__2603\ : InMux
    port map (
            O => \N__12956\,
            I => \N__12934\
        );

    \I__2602\ : InMux
    port map (
            O => \N__12955\,
            I => \N__12931\
        );

    \I__2601\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12928\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__12949\,
            I => \N__12925\
        );

    \I__2599\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12918\
        );

    \I__2598\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12918\
        );

    \I__2597\ : InMux
    port map (
            O => \N__12946\,
            I => \N__12918\
        );

    \I__2596\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12915\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__12942\,
            I => \N__12910\
        );

    \I__2594\ : Span4Mux_h
    port map (
            O => \N__12937\,
            I => \N__12910\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__12934\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__12931\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__12928\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2590\ : Odrv12
    port map (
            O => \N__12925\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__12918\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__12915\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2587\ : Odrv4
    port map (
            O => \N__12910\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__2586\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12889\
        );

    \I__2585\ : InMux
    port map (
            O => \N__12894\,
            I => \N__12885\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12893\,
            I => \N__12869\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12892\,
            I => \N__12869\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__12889\,
            I => \N__12861\
        );

    \I__2581\ : InMux
    port map (
            O => \N__12888\,
            I => \N__12856\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__12885\,
            I => \N__12853\
        );

    \I__2579\ : InMux
    port map (
            O => \N__12884\,
            I => \N__12849\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12883\,
            I => \N__12846\
        );

    \I__2577\ : InMux
    port map (
            O => \N__12882\,
            I => \N__12841\
        );

    \I__2576\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12841\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12880\,
            I => \N__12826\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12879\,
            I => \N__12826\
        );

    \I__2573\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12826\
        );

    \I__2572\ : InMux
    port map (
            O => \N__12877\,
            I => \N__12826\
        );

    \I__2571\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12826\
        );

    \I__2570\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12826\
        );

    \I__2569\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12823\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__12869\,
            I => \N__12820\
        );

    \I__2567\ : InMux
    port map (
            O => \N__12868\,
            I => \N__12817\
        );

    \I__2566\ : InMux
    port map (
            O => \N__12867\,
            I => \N__12810\
        );

    \I__2565\ : InMux
    port map (
            O => \N__12866\,
            I => \N__12810\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12865\,
            I => \N__12810\
        );

    \I__2563\ : InMux
    port map (
            O => \N__12864\,
            I => \N__12807\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__12861\,
            I => \N__12804\
        );

    \I__2561\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12799\
        );

    \I__2560\ : InMux
    port map (
            O => \N__12859\,
            I => \N__12799\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12856\,
            I => \N__12794\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__12853\,
            I => \N__12794\
        );

    \I__2557\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12791\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__12849\,
            I => \N__12784\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__12846\,
            I => \N__12784\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__12841\,
            I => \N__12784\
        );

    \I__2553\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12779\
        );

    \I__2552\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12779\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__12826\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__12823\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2549\ : Odrv4
    port map (
            O => \N__12820\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__12817\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__12810\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__12807\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2545\ : Odrv4
    port map (
            O => \N__12804\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__12799\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__12794\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__12791\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__12784\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__12779\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12751\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__12751\,
            I => \uu2.mem0.g1_0_1_1\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12745\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__12745\,
            I => \uu2.mem0.g1_5_5\
        );

    \I__2535\ : CascadeMux
    port map (
            O => \N__12742\,
            I => \N__12735\
        );

    \I__2534\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12730\
        );

    \I__2533\ : InMux
    port map (
            O => \N__12740\,
            I => \N__12727\
        );

    \I__2532\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12720\
        );

    \I__2531\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12720\
        );

    \I__2530\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12720\
        );

    \I__2529\ : InMux
    port map (
            O => \N__12734\,
            I => \N__12713\
        );

    \I__2528\ : InMux
    port map (
            O => \N__12733\,
            I => \N__12710\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__12730\,
            I => \N__12707\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12704\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12701\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__12719\,
            I => \N__12697\
        );

    \I__2523\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12689\
        );

    \I__2522\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12689\
        );

    \I__2521\ : InMux
    port map (
            O => \N__12716\,
            I => \N__12689\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12686\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__12710\,
            I => \N__12677\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__12707\,
            I => \N__12677\
        );

    \I__2517\ : Span4Mux_v
    port map (
            O => \N__12704\,
            I => \N__12677\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__12701\,
            I => \N__12677\
        );

    \I__2515\ : InMux
    port map (
            O => \N__12700\,
            I => \N__12670\
        );

    \I__2514\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12670\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12670\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__12689\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__2511\ : Odrv4
    port map (
            O => \N__12686\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__12677\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__12670\,
            I => \uu2.w_addr_displaying_3_repZ0Z2\
        );

    \I__2508\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12654\
        );

    \I__2507\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12654\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__12659\,
            I => \N__12650\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__12654\,
            I => \N__12645\
        );

    \I__2504\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12642\
        );

    \I__2503\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12639\
        );

    \I__2502\ : InMux
    port map (
            O => \N__12649\,
            I => \N__12634\
        );

    \I__2501\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12634\
        );

    \I__2500\ : Span4Mux_v
    port map (
            O => \N__12645\,
            I => \N__12631\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__12642\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__12639\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__12634\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__12631\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__12622\,
            I => \N__12619\
        );

    \I__2494\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12616\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__12616\,
            I => \N__12613\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__12613\,
            I => \uu2.mem0.N_74_i\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12604\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__12604\,
            I => \Lab_UT.dispString.dOutP_0_iv_3_0\
        );

    \I__2488\ : CascadeMux
    port map (
            O => \N__12601\,
            I => \uu2.N_84_cascade_\
        );

    \I__2487\ : InMux
    port map (
            O => \N__12598\,
            I => \N__12589\
        );

    \I__2486\ : InMux
    port map (
            O => \N__12597\,
            I => \N__12589\
        );

    \I__2485\ : InMux
    port map (
            O => \N__12596\,
            I => \N__12589\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__12589\,
            I => \N__12583\
        );

    \I__2483\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12573\
        );

    \I__2482\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12573\
        );

    \I__2481\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12573\
        );

    \I__2480\ : Span4Mux_h
    port map (
            O => \N__12583\,
            I => \N__12570\
        );

    \I__2479\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12563\
        );

    \I__2478\ : InMux
    port map (
            O => \N__12581\,
            I => \N__12563\
        );

    \I__2477\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12563\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12560\
        );

    \I__2475\ : Odrv4
    port map (
            O => \N__12570\,
            I => \uu2.N_97\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__12563\,
            I => \uu2.N_97\
        );

    \I__2473\ : Odrv12
    port map (
            O => \N__12560\,
            I => \uu2.N_97\
        );

    \I__2472\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12549\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__12552\,
            I => \N__12545\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__12549\,
            I => \N__12541\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12533\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12533\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12533\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__12541\,
            I => \N__12530\
        );

    \I__2465\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12527\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__12533\,
            I => \N__12520\
        );

    \I__2463\ : Span4Mux_s3_h
    port map (
            O => \N__12530\,
            I => \N__12520\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__12527\,
            I => \N__12520\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__12520\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__12517\,
            I => \uu2.N_97_cascade_\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__12514\,
            I => \N__12511\
        );

    \I__2458\ : InMux
    port map (
            O => \N__12511\,
            I => \N__12506\
        );

    \I__2457\ : InMux
    port map (
            O => \N__12510\,
            I => \N__12503\
        );

    \I__2456\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12500\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__12506\,
            I => \N__12497\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12494\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__12500\,
            I => \uu2.N_159\
        );

    \I__2452\ : Odrv4
    port map (
            O => \N__12497\,
            I => \uu2.N_159\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__12494\,
            I => \uu2.N_159\
        );

    \I__2450\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12478\
        );

    \I__2449\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12478\
        );

    \I__2448\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12478\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__12478\,
            I => \N__12474\
        );

    \I__2446\ : InMux
    port map (
            O => \N__12477\,
            I => \N__12471\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__12474\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__12471\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__2443\ : InMux
    port map (
            O => \N__12466\,
            I => \N__12463\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__12463\,
            I => \N__12460\
        );

    \I__2441\ : Span12Mux_s5_v
    port map (
            O => \N__12460\,
            I => \N__12454\
        );

    \I__2440\ : InMux
    port map (
            O => \N__12459\,
            I => \N__12451\
        );

    \I__2439\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12446\
        );

    \I__2438\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12446\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__12454\,
            I => \L3_tx_data_0\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__12451\,
            I => \L3_tx_data_0\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__12446\,
            I => \L3_tx_data_0\
        );

    \I__2434\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12436\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12432\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__12435\,
            I => \N__12429\
        );

    \I__2431\ : Span4Mux_h
    port map (
            O => \N__12432\,
            I => \N__12426\
        );

    \I__2430\ : InMux
    port map (
            O => \N__12429\,
            I => \N__12423\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__12426\,
            I => \N__12420\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__2427\ : Odrv4
    port map (
            O => \N__12420\,
            I => \uu2.N_86\
        );

    \I__2426\ : Odrv12
    port map (
            O => \N__12417\,
            I => \uu2.N_86\
        );

    \I__2425\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12400\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12400\
        );

    \I__2423\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12400\
        );

    \I__2422\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12400\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__12400\,
            I => \N__12397\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__12397\,
            I => \N__12392\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12387\
        );

    \I__2418\ : InMux
    port map (
            O => \N__12395\,
            I => \N__12387\
        );

    \I__2417\ : Odrv4
    port map (
            O => \N__12392\,
            I => \L3_tx_data_rdy\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__12387\,
            I => \L3_tx_data_rdy\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__12382\,
            I => \uu2.N_86_cascade_\
        );

    \I__2414\ : InMux
    port map (
            O => \N__12379\,
            I => \N__12373\
        );

    \I__2413\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12373\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__12373\,
            I => \N__12370\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__12370\,
            I => \N__12367\
        );

    \I__2410\ : Span4Mux_h
    port map (
            O => \N__12367\,
            I => \N__12362\
        );

    \I__2409\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12359\
        );

    \I__2408\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12356\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__12362\,
            I => \uu2.N_84\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__12359\,
            I => \uu2.N_84\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__12356\,
            I => \uu2.N_84\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__12349\,
            I => \N__12345\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__12348\,
            I => \N__12340\
        );

    \I__2402\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12332\
        );

    \I__2401\ : InMux
    port map (
            O => \N__12344\,
            I => \N__12332\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12343\,
            I => \N__12329\
        );

    \I__2399\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12324\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12324\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12318\
        );

    \I__2396\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12315\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__12332\,
            I => \N__12308\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12329\,
            I => \N__12308\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__12324\,
            I => \N__12308\
        );

    \I__2392\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12305\
        );

    \I__2391\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12302\
        );

    \I__2390\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12299\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__12318\,
            I => \N__12296\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12293\
        );

    \I__2387\ : Span4Mux_v
    port map (
            O => \N__12308\,
            I => \N__12290\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__12305\,
            I => \N__12283\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__12302\,
            I => \N__12283\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12283\
        );

    \I__2383\ : Span4Mux_h
    port map (
            O => \N__12296\,
            I => \N__12277\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__12293\,
            I => \N__12270\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__12290\,
            I => \N__12270\
        );

    \I__2380\ : Span4Mux_h
    port map (
            O => \N__12283\,
            I => \N__12270\
        );

    \I__2379\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12267\
        );

    \I__2378\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12262\
        );

    \I__2377\ : InMux
    port map (
            O => \N__12280\,
            I => \N__12262\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__12277\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__12270\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__12267\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__12262\,
            I => \uu2.w_addr_i_0_tzZ0Z_0\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__12253\,
            I => \uu2.w_addr_i_0_tzZ0Z_0_cascade_\
        );

    \I__2371\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12247\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__12247\,
            I => \N__12243\
        );

    \I__2369\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12240\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__12243\,
            I => \N__12236\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__12240\,
            I => \N__12233\
        );

    \I__2366\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12230\
        );

    \I__2365\ : Odrv4
    port map (
            O => \N__12236\,
            I => \uu2.N_61\
        );

    \I__2364\ : Odrv12
    port map (
            O => \N__12233\,
            I => \uu2.N_61\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__12230\,
            I => \uu2.N_61\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \N__12216\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__12222\,
            I => \N__12212\
        );

    \I__2360\ : CascadeMux
    port map (
            O => \N__12221\,
            I => \N__12207\
        );

    \I__2359\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12201\
        );

    \I__2358\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12201\
        );

    \I__2357\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12198\
        );

    \I__2356\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12181\
        );

    \I__2355\ : InMux
    port map (
            O => \N__12212\,
            I => \N__12181\
        );

    \I__2354\ : InMux
    port map (
            O => \N__12211\,
            I => \N__12181\
        );

    \I__2353\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12181\
        );

    \I__2352\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12181\
        );

    \I__2351\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12181\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__12201\,
            I => \N__12176\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__12198\,
            I => \N__12176\
        );

    \I__2348\ : InMux
    port map (
            O => \N__12197\,
            I => \N__12167\
        );

    \I__2347\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12167\
        );

    \I__2346\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12167\
        );

    \I__2345\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12167\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__12181\,
            I => \N__12164\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__12176\,
            I => \N__12158\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__12167\,
            I => \N__12158\
        );

    \I__2341\ : Span4Mux_h
    port map (
            O => \N__12164\,
            I => \N__12155\
        );

    \I__2340\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12152\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__12158\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2338\ : Odrv4
    port map (
            O => \N__12155\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__12152\,
            I => \uu2.un21_w_addr_displaying_i\
        );

    \I__2336\ : InMux
    port map (
            O => \N__12145\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__2335\ : InMux
    port map (
            O => \N__12142\,
            I => \N__12139\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__12139\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__12136\,
            I => \N__12130\
        );

    \I__2332\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12125\
        );

    \I__2331\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12125\
        );

    \I__2330\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12120\
        );

    \I__2329\ : InMux
    port map (
            O => \N__12130\,
            I => \N__12120\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__12125\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__12120\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__2326\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__2325\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12109\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__12109\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__12106\,
            I => \N__12102\
        );

    \I__2322\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12097\
        );

    \I__2321\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12097\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__12097\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__2319\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12085\
        );

    \I__2318\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12085\
        );

    \I__2317\ : InMux
    port map (
            O => \N__12092\,
            I => \N__12085\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__12085\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__12082\,
            I => \N__12077\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__12081\,
            I => \N__12074\
        );

    \I__2313\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12070\
        );

    \I__2312\ : InMux
    port map (
            O => \N__12077\,
            I => \N__12063\
        );

    \I__2311\ : InMux
    port map (
            O => \N__12074\,
            I => \N__12063\
        );

    \I__2310\ : InMux
    port map (
            O => \N__12073\,
            I => \N__12063\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__12070\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__12063\,
            I => \buart.Z_rx.ser_clk_2\
        );

    \I__2307\ : InMux
    port map (
            O => \N__12058\,
            I => \N__12055\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__12055\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__12052\,
            I => \N__12049\
        );

    \I__2304\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12042\
        );

    \I__2303\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12033\
        );

    \I__2302\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12033\
        );

    \I__2301\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12033\
        );

    \I__2300\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12033\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__12042\,
            I => \buart.Z_rx.ser_clk_3\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__12033\,
            I => \buart.Z_rx.ser_clk_3\
        );

    \I__2297\ : InMux
    port map (
            O => \N__12028\,
            I => \N__12019\
        );

    \I__2296\ : InMux
    port map (
            O => \N__12027\,
            I => \N__12019\
        );

    \I__2295\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12019\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__12013\
        );

    \I__2293\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12006\
        );

    \I__2292\ : InMux
    port map (
            O => \N__12017\,
            I => \N__12006\
        );

    \I__2291\ : InMux
    port map (
            O => \N__12016\,
            I => \N__12006\
        );

    \I__2290\ : Span4Mux_v
    port map (
            O => \N__12013\,
            I => \N__11991\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__12006\,
            I => \N__11991\
        );

    \I__2288\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11976\
        );

    \I__2287\ : InMux
    port map (
            O => \N__12004\,
            I => \N__11976\
        );

    \I__2286\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11976\
        );

    \I__2285\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11976\
        );

    \I__2284\ : InMux
    port map (
            O => \N__12001\,
            I => \N__11976\
        );

    \I__2283\ : InMux
    port map (
            O => \N__12000\,
            I => \N__11976\
        );

    \I__2282\ : InMux
    port map (
            O => \N__11999\,
            I => \N__11976\
        );

    \I__2281\ : InMux
    port map (
            O => \N__11998\,
            I => \N__11971\
        );

    \I__2280\ : InMux
    port map (
            O => \N__11997\,
            I => \N__11971\
        );

    \I__2279\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11968\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__11991\,
            I => \buart.Z_rx.startbit\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__11976\,
            I => \buart.Z_rx.startbit\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__11971\,
            I => \buart.Z_rx.startbit\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__11968\,
            I => \buart.Z_rx.startbit\
        );

    \I__2274\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11953\
        );

    \I__2273\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11953\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__11953\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__2271\ : InMux
    port map (
            O => \N__11950\,
            I => \N__11947\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__11947\,
            I => \N__11944\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__11944\,
            I => \N__11941\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__11941\,
            I => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_2\
        );

    \I__2267\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11933\
        );

    \I__2266\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11927\
        );

    \I__2265\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11927\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__11933\,
            I => \N__11924\
        );

    \I__2263\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11921\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__11927\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__11924\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__11921\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__2259\ : CascadeMux
    port map (
            O => \N__11914\,
            I => \N__11907\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11904\
        );

    \I__2257\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11899\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11899\
        );

    \I__2255\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11896\
        );

    \I__2254\ : InMux
    port map (
            O => \N__11907\,
            I => \N__11893\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__11904\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__11899\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__11896\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__11893\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__2249\ : InMux
    port map (
            O => \N__11884\,
            I => \N__11881\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__11881\,
            I => \N__11875\
        );

    \I__2247\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11867\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11867\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11867\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__11875\,
            I => \N__11864\
        );

    \I__2243\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11861\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__11867\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__11864\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__11861\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__2239\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11851\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__11851\,
            I => \uu2.w_addr_user_3_i_a2_2_6\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__11848\,
            I => \N__11845\
        );

    \I__2236\ : InMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__11842\,
            I => \N__11839\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__11839\,
            I => \N__11836\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__11836\,
            I => \uu2.mem0.N_72_i\
        );

    \I__2232\ : CascadeMux
    port map (
            O => \N__11833\,
            I => \N__11830\
        );

    \I__2231\ : InMux
    port map (
            O => \N__11830\,
            I => \N__11827\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11827\,
            I => \N__11822\
        );

    \I__2229\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11819\
        );

    \I__2228\ : InMux
    port map (
            O => \N__11825\,
            I => \N__11816\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__11822\,
            I => \buart.Z_rx.idle\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__11819\,
            I => \buart.Z_rx.idle\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__11816\,
            I => \buart.Z_rx.idle\
        );

    \I__2224\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11806\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__11806\,
            I => \N__11802\
        );

    \I__2222\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__2221\ : Span4Mux_v
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11799\,
            I => \N__11792\
        );

    \I__2219\ : Span4Mux_v
    port map (
            O => \N__11796\,
            I => \N__11789\
        );

    \I__2218\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11786\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__11792\,
            I => bu_rx_data_rdy
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__11789\,
            I => bu_rx_data_rdy
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__11786\,
            I => bu_rx_data_rdy
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__2213\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11763\
        );

    \I__2212\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11763\
        );

    \I__2211\ : InMux
    port map (
            O => \N__11774\,
            I => \N__11763\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11763\
        );

    \I__2209\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11760\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__11763\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11760\,
            I => \buart.Z_rx.bitcountlde_0\
        );

    \I__2206\ : InMux
    port map (
            O => \N__11755\,
            I => \N__11752\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__11752\,
            I => \buart.Z_rx.un1_sample_0\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__11749\,
            I => \buart.Z_rx.ser_clk_2_cascade_\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__11746\,
            I => \N__11740\
        );

    \I__2202\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11735\
        );

    \I__2201\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11730\
        );

    \I__2200\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11730\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11727\
        );

    \I__2198\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11722\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11722\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__11735\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__11730\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__11727\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__11722\,
            I => \buart.Z_rx.bitcountZ0Z_0\
        );

    \I__2192\ : CEMux
    port map (
            O => \N__11713\,
            I => \N__11709\
        );

    \I__2191\ : CEMux
    port map (
            O => \N__11712\,
            I => \N__11706\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__11709\,
            I => \N__11700\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__11706\,
            I => \N__11700\
        );

    \I__2188\ : CEMux
    port map (
            O => \N__11705\,
            I => \N__11697\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__11700\,
            I => \N__11694\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__11697\,
            I => \N__11691\
        );

    \I__2185\ : Sp12to4
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__2184\ : Sp12to4
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__2183\ : Span12Mux_s7_h
    port map (
            O => \N__11688\,
            I => \N__11680\
        );

    \I__2182\ : Span12Mux_s7_v
    port map (
            O => \N__11685\,
            I => \N__11680\
        );

    \I__2181\ : Odrv12
    port map (
            O => \N__11680\,
            I => \buart.Z_rx.sample\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11673\
        );

    \I__2179\ : InMux
    port map (
            O => \N__11676\,
            I => \N__11670\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__11673\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__11670\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__2176\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11662\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__11662\,
            I => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\
        );

    \I__2174\ : InMux
    port map (
            O => \N__11659\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__2173\ : InMux
    port map (
            O => \N__11656\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11653\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \N__11647\
        );

    \I__2170\ : InMux
    port map (
            O => \N__11647\,
            I => \N__11644\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__11644\,
            I => \N__11641\
        );

    \I__2168\ : Odrv12
    port map (
            O => \N__11641\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11632\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__2164\ : Span4Mux_h
    port map (
            O => \N__11629\,
            I => \N__11626\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__11626\,
            I => \N__11622\
        );

    \I__2162\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11619\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__11622\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__11619\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__2159\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11611\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__11611\,
            I => \Lab_UT.dictrl.next_state_out_0\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__11608\,
            I => \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__11605\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\
        );

    \I__2155\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11599\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11596\
        );

    \I__2153\ : Span12Mux_s8_v
    port map (
            O => \N__11596\,
            I => \N__11593\
        );

    \I__2152\ : Odrv12
    port map (
            O => \N__11593\,
            I => \Lab_UT.dictrl.dicRun_2_reti\
        );

    \I__2151\ : InMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__11587\,
            I => \N__11583\
        );

    \I__2149\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__11583\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_1\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__11580\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_1\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__11575\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_cascade_\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \Lab_UT.m37_ns_cascade_\
        );

    \I__2144\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__11566\,
            I => \Lab_UT.dictrl.next_state_out_2\
        );

    \I__2142\ : SRMux
    port map (
            O => \N__11563\,
            I => \N__11560\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__11560\,
            I => \N__11556\
        );

    \I__2140\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11553\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__11556\,
            I => \N__11550\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__11553\,
            I => \N__11547\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__11550\,
            I => \Lab_UT.m45\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__11547\,
            I => \Lab_UT.m45\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__11542\,
            I => \Lab_UT.m40_cascade_\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__11539\,
            I => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__11536\,
            I => \resetGen_escKey_4_cascade_\
        );

    \I__2132\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11525\
        );

    \I__2131\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11525\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__11531\,
            I => \N__11521\
        );

    \I__2129\ : InMux
    port map (
            O => \N__11530\,
            I => \N__11518\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__11525\,
            I => \N__11515\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11510\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11521\,
            I => \N__11510\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11518\,
            I => \N__11505\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__11515\,
            I => \N__11505\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__11510\,
            I => bu_rx_data_5
        );

    \I__2122\ : Odrv4
    port map (
            O => \N__11505\,
            I => bu_rx_data_5
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__11500\,
            I => \N__11494\
        );

    \I__2120\ : InMux
    port map (
            O => \N__11499\,
            I => \N__11488\
        );

    \I__2119\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11485\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11474\
        );

    \I__2117\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11474\
        );

    \I__2116\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11474\
        );

    \I__2115\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11474\
        );

    \I__2114\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11474\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__11488\,
            I => bu_rx_data_2
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__11485\,
            I => bu_rx_data_2
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__11474\,
            I => bu_rx_data_2
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_\
        );

    \I__2109\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11456\
        );

    \I__2108\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11445\
        );

    \I__2107\ : InMux
    port map (
            O => \N__11462\,
            I => \N__11445\
        );

    \I__2106\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11445\
        );

    \I__2105\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11445\
        );

    \I__2104\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11445\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__11456\,
            I => bu_rx_data_4
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__11445\,
            I => bu_rx_data_4
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__11440\,
            I => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\
        );

    \I__2100\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__11434\,
            I => \resetGen_escKey_2_0\
        );

    \I__2098\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11423\
        );

    \I__2097\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11423\
        );

    \I__2096\ : CascadeMux
    port map (
            O => \N__11429\,
            I => \N__11420\
        );

    \I__2095\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11416\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11423\,
            I => \N__11413\
        );

    \I__2093\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11408\
        );

    \I__2092\ : InMux
    port map (
            O => \N__11419\,
            I => \N__11408\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__11416\,
            I => \N__11401\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__11413\,
            I => \N__11401\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__11408\,
            I => \N__11401\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__11401\,
            I => bu_rx_data_6
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__11398\,
            I => \N__11391\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__11397\,
            I => \N__11388\
        );

    \I__2085\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11383\
        );

    \I__2084\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11374\
        );

    \I__2083\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11374\
        );

    \I__2082\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11374\
        );

    \I__2081\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11374\
        );

    \I__2080\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11369\
        );

    \I__2079\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11369\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__11383\,
            I => bu_rx_data_3
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__11374\,
            I => bu_rx_data_3
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__11369\,
            I => bu_rx_data_3
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__11362\,
            I => \N__11358\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11352\
        );

    \I__2073\ : InMux
    port map (
            O => \N__11358\,
            I => \N__11352\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__11357\,
            I => \N__11348\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__11352\,
            I => \N__11344\
        );

    \I__2070\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11339\
        );

    \I__2069\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11339\
        );

    \I__2068\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11336\
        );

    \I__2067\ : Span4Mux_h
    port map (
            O => \N__11344\,
            I => \N__11333\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11330\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__11336\,
            I => bu_rx_data_7
        );

    \I__2064\ : Odrv4
    port map (
            O => \N__11333\,
            I => bu_rx_data_7
        );

    \I__2063\ : Odrv12
    port map (
            O => \N__11330\,
            I => bu_rx_data_7
        );

    \I__2062\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__11320\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxa_2\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__11317\,
            I => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11311\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11308\
        );

    \I__2057\ : Span4Mux_v
    port map (
            O => \N__11308\,
            I => \N__11305\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__11305\,
            I => \Lab_UT.didp.countrce2.N_183\
        );

    \I__2055\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11299\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__11299\,
            I => \Lab_UT.didp.countrce2.N_180\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__11296\,
            I => \Lab_UT.didp.countrce4.N_80_i_cascade_\
        );

    \I__2052\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11290\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__11290\,
            I => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_3\
        );

    \I__2050\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__11284\,
            I => \Lab_UT.bcd2segment4.segment_i_0Z0Z_6\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__11278\,
            I => \Lab_UT.dictrl.next_alarmstate4_1Z0Z_0\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__11275\,
            I => \Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_\
        );

    \I__2045\ : InMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__11269\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__2043\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11259\
        );

    \I__2042\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11253\
        );

    \I__2041\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11250\
        );

    \I__2040\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11247\
        );

    \I__2039\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11244\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__11259\,
            I => \N__11241\
        );

    \I__2037\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11234\
        );

    \I__2036\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11234\
        );

    \I__2035\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11234\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__11253\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__11250\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__11247\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__11244\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2030\ : Odrv4
    port map (
            O => \N__11241\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__11234\,
            I => \uu2.w_addr_displaying_1_repZ0Z1\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__11221\,
            I => \uu2.N_7_cascade_\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__11218\,
            I => \N__11215\
        );

    \I__2026\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11212\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11209\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__11209\,
            I => \uu2.N_10\
        );

    \I__2023\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11202\
        );

    \I__2022\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11195\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__11202\,
            I => \N__11192\
        );

    \I__2020\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11187\
        );

    \I__2019\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11187\
        );

    \I__2018\ : InMux
    port map (
            O => \N__11199\,
            I => \N__11182\
        );

    \I__2017\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11182\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__11195\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__11192\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__11187\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__11182\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__2012\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11170\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__11170\,
            I => \uu2.N_8\
        );

    \I__2010\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11164\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__11164\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__2008\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11158\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__11158\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__2006\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11152\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__11152\,
            I => \Lab_UT.didp.countrce2.N_178\
        );

    \I__2004\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__11146\,
            I => \N__11143\
        );

    \I__2002\ : Odrv12
    port map (
            O => \N__11143\,
            I => \Lab_UT.didp.countrce2.N_175\
        );

    \I__2001\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11137\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__11137\,
            I => \N__11134\
        );

    \I__1999\ : Span4Mux_h
    port map (
            O => \N__11134\,
            I => \N__11131\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__11131\,
            I => \Lab_UT.didp.countrce2.N_170\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_\
        );

    \I__1996\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11122\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__11122\,
            I => \N__11119\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__11119\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_45\
        );

    \I__1993\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11106\
        );

    \I__1992\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11103\
        );

    \I__1991\ : InMux
    port map (
            O => \N__11114\,
            I => \N__11100\
        );

    \I__1990\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11095\
        );

    \I__1989\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11095\
        );

    \I__1988\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11090\
        );

    \I__1987\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11090\
        );

    \I__1986\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11087\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__11106\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__11103\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__11100\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__11095\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__11090\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__11087\,
            I => \uu2.w_addr_displaying_2_repZ0Z1\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__1978\ : InMux
    port map (
            O => \N__11071\,
            I => \N__11068\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__11068\,
            I => \N__11060\
        );

    \I__1976\ : InMux
    port map (
            O => \N__11067\,
            I => \N__11054\
        );

    \I__1975\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11051\
        );

    \I__1974\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11048\
        );

    \I__1973\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11045\
        );

    \I__1972\ : InMux
    port map (
            O => \N__11063\,
            I => \N__11042\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__11060\,
            I => \N__11039\
        );

    \I__1970\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11032\
        );

    \I__1969\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11032\
        );

    \I__1968\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11032\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__11054\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__11051\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__11048\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__11045\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__11042\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1962\ : Odrv4
    port map (
            O => \N__11039\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__11032\,
            I => \uu2.w_addr_displaying_3_repZ0Z1\
        );

    \I__1960\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11014\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__11014\,
            I => \uu2.bitmap_pmux_sn_N_31_0\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__11011\,
            I => \uu2.bitmap_pmux_sn_N_31_0_cascade_\
        );

    \I__1957\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10999\
        );

    \I__1956\ : InMux
    port map (
            O => \N__11007\,
            I => \N__10999\
        );

    \I__1955\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10999\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__10999\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__1953\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10993\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__10993\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_48\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__10990\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_\
        );

    \I__1950\ : InMux
    port map (
            O => \N__10987\,
            I => \N__10984\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10984\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_47\
        );

    \I__1948\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__10978\,
            I => \N__10975\
        );

    \I__1946\ : Odrv4
    port map (
            O => \N__10975\,
            I => \uu2.mem0.bitmap_pmux_u_ns_1\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__10972\,
            I => \uu2.mem0.g0_5_3_cascade_\
        );

    \I__1944\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10966\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__10966\,
            I => \uu2.mem0.g0_5_6\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__10963\,
            I => \Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__10960\,
            I => \uu2.un31_w_data_displaying_0_a2_1_cascade_\
        );

    \I__1940\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10950\
        );

    \I__1939\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10950\
        );

    \I__1938\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10947\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__10950\,
            I => \N__10944\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__10947\,
            I => \N__10941\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__10944\,
            I => \N__10936\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__10941\,
            I => \N__10936\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__10936\,
            I => \uu2.un31_w_data_displaying\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__10930\,
            I => \uu2.un15_w_data_displaying_6\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__10927\,
            I => \uu2.un15_w_data_displaying_6_cascade_\
        );

    \I__1929\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10920\
        );

    \I__1928\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10917\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__10920\,
            I => \N__10912\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10912\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__10912\,
            I => \uu2.un49_w_data_displaying_1\
        );

    \I__1924\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10905\
        );

    \I__1923\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10902\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__10905\,
            I => \N__10899\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__10902\,
            I => \N__10896\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__10899\,
            I => \N__10893\
        );

    \I__1919\ : Span4Mux_h
    port map (
            O => \N__10896\,
            I => \N__10890\
        );

    \I__1918\ : Odrv4
    port map (
            O => \N__10893\,
            I => \uu2.un49_w_data_displaying\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__10890\,
            I => \uu2.un49_w_data_displaying\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__10885\,
            I => \N__10881\
        );

    \I__1915\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10877\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10872\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10872\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__10877\,
            I => \N__10869\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__10872\,
            I => \N__10864\
        );

    \I__1910\ : Span4Mux_h
    port map (
            O => \N__10869\,
            I => \N__10864\
        );

    \I__1909\ : Odrv4
    port map (
            O => \N__10864\,
            I => \uu2.un15_w_data_displaying_i_i_o2_0\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__10861\,
            I => \uu2.un15_w_data_displaying_i_i_o2_0_cascade_\
        );

    \I__1907\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10855\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__10855\,
            I => \uu2.mem0.un49_w_data_displaying_0\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__10852\,
            I => \N__10849\
        );

    \I__1904\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10843\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__10843\,
            I => \uu2.mem0.g0_5_5\
        );

    \I__1901\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10837\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__10837\,
            I => \uu2.mem0.un31_w_data_displaying_0\
        );

    \I__1899\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10831\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__10831\,
            I => \N__10828\
        );

    \I__1897\ : Span4Mux_h
    port map (
            O => \N__10828\,
            I => \N__10825\
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__10825\,
            I => \uu2.mem0.g1_1_1\
        );

    \I__1895\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10818\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__10818\,
            I => \N__10810\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10807\
        );

    \I__1891\ : CascadeMux
    port map (
            O => \N__10814\,
            I => \N__10800\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10796\
        );

    \I__1889\ : Span4Mux_h
    port map (
            O => \N__10810\,
            I => \N__10791\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__10807\,
            I => \N__10791\
        );

    \I__1887\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10788\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10783\
        );

    \I__1885\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10783\
        );

    \I__1884\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10776\
        );

    \I__1883\ : InMux
    port map (
            O => \N__10800\,
            I => \N__10776\
        );

    \I__1882\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10776\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10796\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__10791\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__10788\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__10783\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__10776\,
            I => \uu2.w_addr_displaying_7_repZ0Z1\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10765\,
            I => \N__10753\
        );

    \I__1875\ : InMux
    port map (
            O => \N__10764\,
            I => \N__10753\
        );

    \I__1874\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10748\
        );

    \I__1873\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10748\
        );

    \I__1872\ : InMux
    port map (
            O => \N__10761\,
            I => \N__10745\
        );

    \I__1871\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10742\
        );

    \I__1870\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10737\
        );

    \I__1869\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10737\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__10753\,
            I => \N__10734\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__10748\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__10745\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__10742\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__10737\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__10734\,
            I => \uu2.w_addr_displaying_8_repZ0Z1\
        );

    \I__1862\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10720\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__10720\,
            I => \N__10711\
        );

    \I__1860\ : InMux
    port map (
            O => \N__10719\,
            I => \N__10704\
        );

    \I__1859\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10704\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10704\
        );

    \I__1857\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10701\
        );

    \I__1856\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10696\
        );

    \I__1855\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10696\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__10711\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__10704\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10701\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__10696\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__10687\,
            I => \N__10679\
        );

    \I__1849\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10676\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__10685\,
            I => \N__10673\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__10684\,
            I => \N__10670\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__10683\,
            I => \N__10667\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__10682\,
            I => \N__10664\
        );

    \I__1844\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10661\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__10676\,
            I => \N__10658\
        );

    \I__1842\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10655\
        );

    \I__1841\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10648\
        );

    \I__1840\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10648\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10648\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__10661\,
            I => \N__10645\
        );

    \I__1837\ : Span4Mux_h
    port map (
            O => \N__10658\,
            I => \N__10642\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__10655\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__10648\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__10645\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__10642\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__1832\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10630\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__1830\ : Span4Mux_h
    port map (
            O => \N__10627\,
            I => \N__10624\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__10624\,
            I => \uu2.mem0.N_111\
        );

    \I__1828\ : CEMux
    port map (
            O => \N__10621\,
            I => \N__10618\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__10618\,
            I => \N__10614\
        );

    \I__1826\ : CEMux
    port map (
            O => \N__10617\,
            I => \N__10611\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__10614\,
            I => \N__10608\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__10611\,
            I => \N__10605\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__10608\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__1822\ : Odrv12
    port map (
            O => \N__10605\,
            I => \uu2.un28_w_addr_user_i_0_0\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__10600\,
            I => \N__10597\
        );

    \I__1820\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10594\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__10594\,
            I => \N__10591\
        );

    \I__1818\ : Span4Mux_h
    port map (
            O => \N__10591\,
            I => \N__10588\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__10588\,
            I => \uu2.mem0.N_73_i\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__10585\,
            I => \buart.Z_rx.bitcount_lm_2_cascade_\
        );

    \I__1815\ : InMux
    port map (
            O => \N__10582\,
            I => \N__10572\
        );

    \I__1814\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10572\
        );

    \I__1813\ : InMux
    port map (
            O => \N__10580\,
            I => \N__10569\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10566\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10561\
        );

    \I__1810\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10561\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__10572\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__10569\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__10566\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__10561\,
            I => \buart.Z_rx.bitcountZ0Z_2\
        );

    \I__1805\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10549\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__10549\,
            I => \buart.Z_rx.bitcount_lm_4\
        );

    \I__1803\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10539\
        );

    \I__1802\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10536\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10533\
        );

    \I__1800\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10528\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10542\,
            I => \N__10528\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__10539\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10536\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__10533\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__10528\,
            I => \buart.Z_rx.bitcountZ0Z_4\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__10519\,
            I => \N__10516\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10513\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__10513\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__1791\ : CascadeMux
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__1790\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10497\
        );

    \I__1789\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10497\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10497\
        );

    \I__1787\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10494\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__10497\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__10494\,
            I => \buart.Z_rx.N_27_0_i\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__10489\,
            I => \buart.Z_rx.bitcount_lm_3_cascade_\
        );

    \I__1783\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10476\
        );

    \I__1782\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10476\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10473\
        );

    \I__1780\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10470\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10465\
        );

    \I__1778\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10465\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__10476\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10473\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__10470\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__10465\,
            I => \buart.Z_rx.bitcountZ0Z_3\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10453\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__10453\,
            I => \uu2.N_153\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__10450\,
            I => \uu2.N_90_cascade_\
        );

    \I__1770\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10444\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__10444\,
            I => \uu2.N_105\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__10441\,
            I => \N__10436\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__10440\,
            I => \N__10432\
        );

    \I__1766\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10429\
        );

    \I__1765\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10426\
        );

    \I__1764\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10421\
        );

    \I__1763\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10421\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__10429\,
            I => \uu2.N_90\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__10426\,
            I => \uu2.N_90\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10421\,
            I => \uu2.N_90\
        );

    \I__1759\ : SRMux
    port map (
            O => \N__10414\,
            I => \N__10409\
        );

    \I__1758\ : IoInMux
    port map (
            O => \N__10413\,
            I => \N__10406\
        );

    \I__1757\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10403\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__10409\,
            I => \N__10400\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__10406\,
            I => \N__10397\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__10403\,
            I => \N__10394\
        );

    \I__1753\ : Span4Mux_v
    port map (
            O => \N__10400\,
            I => \N__10391\
        );

    \I__1752\ : Span4Mux_s2_v
    port map (
            O => \N__10397\,
            I => \N__10388\
        );

    \I__1751\ : Span4Mux_s2_v
    port map (
            O => \N__10394\,
            I => \N__10383\
        );

    \I__1750\ : Span4Mux_s2_v
    port map (
            O => \N__10391\,
            I => \N__10383\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__10388\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__10383\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__10378\,
            I => \buart.Z_rx.N_27_0_i_cascade_\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__10375\,
            I => \buart.Z_rx.bitcount_lm_0_cascade_\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__10372\,
            I => \N__10369\
        );

    \I__1744\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10366\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__10366\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__10363\,
            I => \buart.Z_rx.bitcount_lm_1_cascade_\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__10360\,
            I => \N__10352\
        );

    \I__1740\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10347\
        );

    \I__1739\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10347\
        );

    \I__1738\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10344\
        );

    \I__1737\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10339\
        );

    \I__1736\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10339\
        );

    \I__1735\ : InMux
    port map (
            O => \N__10352\,
            I => \N__10336\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__10347\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__10344\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__10339\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__10336\,
            I => \buart.Z_rx.bitcountZ0Z_1\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__10327\,
            I => \N__10324\
        );

    \I__1729\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10321\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__10321\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__10318\,
            I => \Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_\
        );

    \I__1726\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10312\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10312\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__1724\ : InMux
    port map (
            O => \N__10309\,
            I => \N__10306\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__10306\,
            I => \Lab_UT.bcd2segment3.segment_i_0Z0Z_1\
        );

    \I__1722\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10300\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__10300\,
            I => \Lab_UT.bcd2segment3.segment_i_0Z0Z_2\
        );

    \I__1720\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__1718\ : Span4Mux_h
    port map (
            O => \N__10291\,
            I => \N__10288\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__10288\,
            I => \resetGen.escKeyZ0Z_3\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__10285\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__10282\,
            I => \uu2.N_4_cascade_\
        );

    \I__1714\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__10276\,
            I => \N__10273\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__10273\,
            I => \uu2.g0_17_1\
        );

    \I__1711\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10267\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__10267\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__1709\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10261\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__10261\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__1707\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10255\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__10255\,
            I => \uu2.N_5\
        );

    \I__1705\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10249\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__10249\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__10246\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_\
        );

    \I__1702\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10236\
        );

    \I__1701\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10233\
        );

    \I__1700\ : InMux
    port map (
            O => \N__10241\,
            I => \N__10226\
        );

    \I__1699\ : InMux
    port map (
            O => \N__10240\,
            I => \N__10226\
        );

    \I__1698\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10226\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__10236\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__10233\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__10226\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__1694\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10216\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__10216\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__1692\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10210\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__10210\,
            I => \uu2.bitmap_RNISSSNZ0Z_162\
        );

    \I__1690\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__10204\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__10201\,
            I => \uu2.N_46_cascade_\
        );

    \I__1687\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10193\
        );

    \I__1686\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10190\
        );

    \I__1685\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10187\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__10193\,
            I => \N__10184\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__10190\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__10187\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__10184\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__1680\ : InMux
    port map (
            O => \N__10177\,
            I => \N__10171\
        );

    \I__1679\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10171\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__10168\
        );

    \I__1677\ : Span4Mux_h
    port map (
            O => \N__10168\,
            I => \N__10165\
        );

    \I__1676\ : Odrv4
    port map (
            O => \N__10165\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__10162\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__10159\,
            I => \N__10156\
        );

    \I__1673\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10153\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__10153\,
            I => \N__10150\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__10150\,
            I => \N__10147\
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__10147\,
            I => \uu2.un426_ci\
        );

    \I__1669\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__1668\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10133\
        );

    \I__1667\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10133\
        );

    \I__1666\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10130\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__10138\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__10133\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__10130\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__1662\ : InMux
    port map (
            O => \N__10123\,
            I => \N__10120\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10117\
        );

    \I__1660\ : Span4Mux_h
    port map (
            O => \N__10117\,
            I => \N__10114\
        );

    \I__1659\ : Odrv4
    port map (
            O => \N__10114\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_2\
        );

    \I__1658\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10108\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__10108\,
            I => \N__10105\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__10105\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \uu2.mem0.g0_7_3_cascade_\
        );

    \I__1654\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10096\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__10096\,
            I => \uu2.bitmap_pmux_27_ns_1_0\
        );

    \I__1652\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10090\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__10090\,
            I => \uu2.mem0.g0_6_4\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__10087\,
            I => \uu2.mem0.g0_6_5_cascade_\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__10084\,
            I => \uu2.N_150_cascade_\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__10081\,
            I => \N__10078\
        );

    \I__1647\ : InMux
    port map (
            O => \N__10078\,
            I => \N__10073\
        );

    \I__1646\ : InMux
    port map (
            O => \N__10077\,
            I => \N__10070\
        );

    \I__1645\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10067\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__10073\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__10070\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__10067\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__1640\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10054\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__1638\ : Odrv4
    port map (
            O => \N__10051\,
            I => \uu2.mem0.N_78_i_0\
        );

    \I__1637\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10044\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__10047\,
            I => \N__10041\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__10044\,
            I => \N__10038\
        );

    \I__1634\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10035\
        );

    \I__1633\ : Span4Mux_v
    port map (
            O => \N__10038\,
            I => \N__10032\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__10035\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__10032\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__10027\,
            I => \N__10024\
        );

    \I__1629\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10019\
        );

    \I__1628\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10014\
        );

    \I__1627\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10014\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__10019\,
            I => \uu2.N_93\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__10014\,
            I => \uu2.N_93\
        );

    \I__1624\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10003\
        );

    \I__1623\ : InMux
    port map (
            O => \N__10008\,
            I => \N__10000\
        );

    \I__1622\ : InMux
    port map (
            O => \N__10007\,
            I => \N__9997\
        );

    \I__1621\ : InMux
    port map (
            O => \N__10006\,
            I => \N__9994\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__10003\,
            I => \N__9991\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__10000\,
            I => \N__9988\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__9997\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__9994\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__9991\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__9988\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__1614\ : InMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__9976\,
            I => \N__9973\
        );

    \I__1612\ : Span12Mux_s7_v
    port map (
            O => \N__9973\,
            I => \N__9969\
        );

    \I__1611\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9966\
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__9969\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__9966\,
            I => \buart.Z_rx.hhZ0Z_1\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9957\
        );

    \I__1607\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9954\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9951\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__9954\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1604\ : Odrv4
    port map (
            O => \N__9951\,
            I => \buart.Z_rx.hhZ0Z_0\
        );

    \I__1603\ : InMux
    port map (
            O => \N__9946\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__1602\ : InMux
    port map (
            O => \N__9943\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__1601\ : InMux
    port map (
            O => \N__9940\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9937\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9934\,
            I => \N__9931\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__9931\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__9928\,
            I => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\
        );

    \I__1596\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__9922\,
            I => \N__9919\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__9919\,
            I => \uu2.bitmap_pmux_sn_N_15\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__9916\,
            I => \uu2.N_395_cascade_\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__9910\,
            I => \uu2.N_56\
        );

    \I__1590\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9904\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__9904\,
            I => \N__9900\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9897\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9891\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__9894\,
            I => \uu2.N_401\
        );

    \I__1584\ : Odrv12
    port map (
            O => \N__9891\,
            I => \uu2.N_401\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__9886\,
            I => \buart.Z_rx.idle_1_cascade_\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \buart.Z_rx.valid_1_cascade_\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__9880\,
            I => \N__9875\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__9879\,
            I => \N__9872\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \N__9869\
        );

    \I__1578\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9864\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9864\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9869\,
            I => \N__9861\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__9864\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__9861\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9850\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9850\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__9850\,
            I => \uu2.N_383\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9847\,
            I => \N__9844\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__9844\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__9841\,
            I => \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__9838\,
            I => \Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9832\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__9832\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9826\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__9826\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__1562\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9820\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__9820\,
            I => \uu2.bitmap_pmux_15_i_m2_ns_1\
        );

    \I__1560\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9814\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__9814\,
            I => \uu2.mem0.g1_3_0\
        );

    \I__1558\ : InMux
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__1557\ : InMux
    port map (
            O => \N__9810\,
            I => \N__9805\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9802\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__9802\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__1554\ : InMux
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__1553\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9793\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9790\
        );

    \I__1551\ : Odrv4
    port map (
            O => \N__9790\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__9787\,
            I => \uu2.N_247_cascade_\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__1548\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9775\
        );

    \I__1547\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9775\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__9775\,
            I => \uu2.N_2171_0\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__9769\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_44\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__9763\,
            I => \Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_\
        );

    \I__1541\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9757\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__9757\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__1538\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9748\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__9748\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__9745\,
            I => \uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__9742\,
            I => \N__9738\
        );

    \I__1534\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9735\
        );

    \I__1533\ : InMux
    port map (
            O => \N__9738\,
            I => \N__9732\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__9735\,
            I => \uu2.g2_0_0\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__9732\,
            I => \uu2.g2_0_0\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__9727\,
            I => \uu2.mem0.g1_6_cascade_\
        );

    \I__1529\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9721\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__9721\,
            I => \uu2.mem0.N_1201_0_0_0\
        );

    \I__1527\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9715\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__9715\,
            I => \uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9706\
        );

    \I__1524\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9706\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__9706\,
            I => \uu2.bitmap_pmux_sn_N_20_0\
        );

    \I__1522\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9700\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__9700\,
            I => \N__9697\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__9697\,
            I => \uu2.bitmap_pmux_19_i_m2_ns_1\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9691\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__9691\,
            I => \uu2.N_55_0\
        );

    \I__1517\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__9685\,
            I => \uu2.mem0.bitmap_pmux_sn_N_20_1_0_1\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9679\,
            I => \uu2.mem0.N_2166_1_0_1\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__9676\,
            I => \uu2.mem0.N_247_0_cascade_\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \uu2.mem0.N_2171_1_0_1_cascade_\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9667\
        );

    \I__1510\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1509\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9661\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__9661\,
            I => \N__9657\
        );

    \I__1507\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9654\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__9657\,
            I => \uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__9654\,
            I => \uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7\
        );

    \I__1504\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9646\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__9646\,
            I => \uu2.mem0.N_397_1_0_1\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__9643\,
            I => \uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_\
        );

    \I__1501\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9637\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__9637\,
            I => \uu2.mem0.g1_2_0\
        );

    \I__1499\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9631\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__9631\,
            I => \uu2.N_40_0\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__9628\,
            I => \N__9625\
        );

    \I__1496\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__9622\,
            I => \uu2.N_48_i_0\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9616\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__9616\,
            I => \uu2.N_404\
        );

    \I__1492\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__9610\,
            I => \uu2.mem0.g1_1_1_0\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__9607\,
            I => \uu2.N_404_cascade_\
        );

    \I__1489\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9601\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__9601\,
            I => \uu2.mem0.bitmap_pmux_1_0_0\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__9598\,
            I => \uu2.mem0.bitmap_pmux_sn_N_42_cascade_\
        );

    \I__1486\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9592\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__9592\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_46\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__9589\,
            I => \uu2.bitmap_pmux_20_ns_1_cascade_\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__9586\,
            I => \N__9583\
        );

    \I__1482\ : InMux
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__9580\,
            I => \Lab_UT.bcd2segment4.segment_0Z0Z_2\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9574\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__9574\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__9571\,
            I => \Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9565\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__9565\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__1475\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9559\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__9559\,
            I => \Lab_UT.bcd2segment4.N_217\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__9556\,
            I => \N__9553\
        );

    \I__1472\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__9550\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__1470\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9544\
        );

    \I__1469\ : LocalMux
    port map (
            O => \N__9544\,
            I => \Lab_UT.bcd2segment4.segment_i_1Z0Z_5\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9538\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__9538\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__9535\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__9532\,
            I => \N__9529\
        );

    \I__1464\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__9523\,
            I => \N__9516\
        );

    \I__1461\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9511\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9511\
        );

    \I__1459\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9506\
        );

    \I__1458\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9506\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__9516\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__9511\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__9506\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__9499\,
            I => \N__9496\
        );

    \I__1453\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9493\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__9493\,
            I => \N__9490\
        );

    \I__1451\ : Span4Mux_s3_h
    port map (
            O => \N__9490\,
            I => \N__9484\
        );

    \I__1450\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9481\
        );

    \I__1449\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9478\
        );

    \I__1448\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9475\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__9484\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__9481\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__9478\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__9475\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1443\ : CEMux
    port map (
            O => \N__9466\,
            I => \N__9463\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__9463\,
            I => \N__9460\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__9460\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__9457\,
            I => \N__9454\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9451\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__9451\,
            I => \N__9448\
        );

    \I__1437\ : Span4Mux_s3_h
    port map (
            O => \N__9448\,
            I => \N__9445\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__9445\,
            I => \uu2.mem0.N_70_i\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__9442\,
            I => \N__9439\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9436\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__9436\,
            I => \N__9431\
        );

    \I__1432\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9425\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9425\
        );

    \I__1430\ : Span4Mux_h
    port map (
            O => \N__9431\,
            I => \N__9422\
        );

    \I__1429\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9419\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__9425\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1427\ : Odrv4
    port map (
            O => \N__9422\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__9419\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__9412\,
            I => \N__9409\
        );

    \I__1424\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9401\
        );

    \I__1422\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9398\
        );

    \I__1421\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9395\
        );

    \I__1420\ : Span4Mux_v
    port map (
            O => \N__9401\,
            I => \N__9392\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__9398\,
            I => \N__9387\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__9395\,
            I => \N__9387\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__9392\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__9387\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1415\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__9379\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__1413\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9372\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__9375\,
            I => \N__9367\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9372\,
            I => \N__9364\
        );

    \I__1410\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9361\
        );

    \I__1409\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9358\
        );

    \I__1408\ : InMux
    port map (
            O => \N__9367\,
            I => \N__9355\
        );

    \I__1407\ : Span4Mux_h
    port map (
            O => \N__9364\,
            I => \N__9352\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__9361\,
            I => \N__9347\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__9358\,
            I => \N__9347\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__9355\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__9352\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__9347\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1401\ : InMux
    port map (
            O => \N__9340\,
            I => \N__9336\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__9339\,
            I => \N__9332\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9329\
        );

    \I__1398\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9324\
        );

    \I__1397\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9321\
        );

    \I__1396\ : Span4Mux_h
    port map (
            O => \N__9329\,
            I => \N__9318\
        );

    \I__1395\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9313\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9313\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9324\,
            I => \N__9310\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__9321\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__9318\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__9313\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1389\ : Odrv12
    port map (
            O => \N__9310\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__1387\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9295\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__9295\,
            I => \N__9290\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__9294\,
            I => \N__9287\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__9293\,
            I => \N__9284\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__9290\,
            I => \N__9281\
        );

    \I__1382\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9278\
        );

    \I__1381\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9275\
        );

    \I__1380\ : Odrv4
    port map (
            O => \N__9281\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__9278\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__9275\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1377\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9264\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__9267\,
            I => \N__9260\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__9264\,
            I => \N__9257\
        );

    \I__1374\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9251\
        );

    \I__1373\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9248\
        );

    \I__1372\ : Span4Mux_h
    port map (
            O => \N__9257\,
            I => \N__9245\
        );

    \I__1371\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9238\
        );

    \I__1370\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9238\
        );

    \I__1369\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9238\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9235\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__9248\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__9245\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__9238\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1364\ : Odrv12
    port map (
            O => \N__9235\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1362\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9216\
        );

    \I__1361\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9211\
        );

    \I__1360\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9211\
        );

    \I__1359\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9206\
        );

    \I__1358\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9206\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__9216\,
            I => \uu2.un404_ci\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__9211\,
            I => \uu2.un404_ci\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__9206\,
            I => \uu2.un404_ci\
        );

    \I__1354\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9196\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__9196\,
            I => \N__9190\
        );

    \I__1352\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9187\
        );

    \I__1351\ : InMux
    port map (
            O => \N__9194\,
            I => \N__9182\
        );

    \I__1350\ : InMux
    port map (
            O => \N__9193\,
            I => \N__9182\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__9190\,
            I => \N__9179\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__9187\,
            I => \o_One_Sec_Pulse\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__9182\,
            I => \o_One_Sec_Pulse\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__9179\,
            I => \o_One_Sec_Pulse\
        );

    \I__1345\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__9169\,
            I => \N__9165\
        );

    \I__1343\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9162\
        );

    \I__1342\ : Span4Mux_s3_h
    port map (
            O => \N__9165\,
            I => \N__9159\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__9162\,
            I => \N__9154\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__9159\,
            I => \N__9151\
        );

    \I__1339\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9146\
        );

    \I__1338\ : InMux
    port map (
            O => \N__9157\,
            I => \N__9146\
        );

    \I__1337\ : Span4Mux_v
    port map (
            O => \N__9154\,
            I => \N__9143\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__9151\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__9146\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__9143\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__1333\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9133\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__9133\,
            I => \N__9129\
        );

    \I__1331\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9126\
        );

    \I__1330\ : Span4Mux_s3_h
    port map (
            O => \N__9129\,
            I => \N__9123\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__9126\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__9123\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__1327\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__1324\ : Odrv4
    port map (
            O => \N__9109\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__1322\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9092\
        );

    \I__1321\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9092\
        );

    \I__1320\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9092\
        );

    \I__1319\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9089\
        );

    \I__1318\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9086\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9082\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9079\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__9086\,
            I => \N__9076\
        );

    \I__1314\ : InMux
    port map (
            O => \N__9085\,
            I => \N__9073\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__9082\,
            I => \N__9070\
        );

    \I__1312\ : Span4Mux_s3_h
    port map (
            O => \N__9079\,
            I => \N__9067\
        );

    \I__1311\ : Span4Mux_s3_h
    port map (
            O => \N__9076\,
            I => \N__9064\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__9073\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1309\ : Odrv4
    port map (
            O => \N__9070\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__9067\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__9064\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__1306\ : InMux
    port map (
            O => \N__9055\,
            I => \N__9052\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__1304\ : IoSpan4Mux
    port map (
            O => \N__9049\,
            I => \N__9046\
        );

    \I__1303\ : IoSpan4Mux
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__1302\ : IoSpan4Mux
    port map (
            O => \N__9043\,
            I => \N__9040\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__9040\,
            I => \uart_RXD\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__1299\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__1297\ : Span4Mux_h
    port map (
            O => \N__9028\,
            I => \N__9024\
        );

    \I__1296\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9021\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__9024\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__9021\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__1292\ : InMux
    port map (
            O => \N__9013\,
            I => \N__9010\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__9010\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1290\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__9004\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__1288\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8998\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__8998\,
            I => \uu2.bitmap_RNI8LB51Z0Z_186\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__8995\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__8992\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__8989\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__8983\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__1280\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8974\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__8974\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__1278\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8968\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__8968\,
            I => \uu2.mem0.bitmap_pmux_sn_i7_mux_0\
        );

    \I__1276\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8962\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__8962\,
            I => \N__8959\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__8959\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__8956\,
            I => \Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_\
        );

    \I__1272\ : CascadeMux
    port map (
            O => \N__8953\,
            I => \uu2.bitmap_RNIMQ601Z0Z_58_cascade_\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__8950\,
            I => \Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__8944\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__1268\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8938\
        );

    \I__1267\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8935\,
            I => \uu2.mem0.N_71_i\
        );

    \I__1265\ : InMux
    port map (
            O => \N__8932\,
            I => \N__8929\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8929\,
            I => \uu2.mem0.w_data_1\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__8926\,
            I => \N__8923\
        );

    \I__1262\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8920\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8917\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__8917\,
            I => \uu2.mem0.N_76_i_0\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__8914\,
            I => \uu2.mem0.N_2166_0_cascade_\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__8911\,
            I => \uu2.mem0.bitmap_pmux_0_cascade_\
        );

    \I__1257\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__8905\,
            I => \N__8902\
        );

    \I__1255\ : Span4Mux_s3_h
    port map (
            O => \N__8902\,
            I => \N__8899\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__8899\,
            I => \uu2.mem0.w_data_3\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8893\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__8893\,
            I => \uu2.mem0.ram512X8_inst_RNOZ0Z_42\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__8884\,
            I => \N__8881\
        );

    \I__1248\ : Odrv4
    port map (
            O => \N__8881\,
            I => \uu2.mem0.N_75_i\
        );

    \I__1247\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8875\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__8875\,
            I => \uu2.N_361\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__8872\,
            I => \uu2.N_361_cascade_\
        );

    \I__1244\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__8866\,
            I => \uu2.mem0.w_data_4\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8860\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__8860\,
            I => \N__8857\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__8857\,
            I => \uu2.mem0.N_69_i\
        );

    \I__1239\ : InMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__8851\,
            I => \uu2.mem0.w_data_0_a3_0_4\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__8848\,
            I => \uu2.N_61_cascade_\
        );

    \I__1236\ : CascadeMux
    port map (
            O => \N__8845\,
            I => \uu2.mem0.un51_w_data_displaying_cascade_\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8839\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__8839\,
            I => \uu2.mem0.w_data_5\
        );

    \I__1233\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__8833\,
            I => \uu2.mem0.w_data_6\
        );

    \I__1231\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8826\
        );

    \I__1230\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8823\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__8826\,
            I => \N__8820\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__8823\,
            I => \N__8817\
        );

    \I__1227\ : Span4Mux_h
    port map (
            O => \N__8820\,
            I => \N__8814\
        );

    \I__1226\ : Odrv12
    port map (
            O => \N__8817\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1225\ : Odrv4
    port map (
            O => \N__8814\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__8806\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8797\
        );

    \I__1221\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8797\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__8797\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__8794\,
            I => \N__8791\
        );

    \I__1218\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8783\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8783\
        );

    \I__1216\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8780\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8777\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8771\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__8780\,
            I => \N__8771\
        );

    \I__1212\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8766\
        );

    \I__1211\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8766\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__8771\,
            I => \N__8763\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__8766\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1208\ : Odrv4
    port map (
            O => \N__8763\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__8758\,
            I => \uu2.trig_rd_is_det_cascade_\
        );

    \I__1206\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8750\
        );

    \I__1205\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8745\
        );

    \I__1204\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8745\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8742\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8737\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__8742\,
            I => \N__8737\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__8737\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__1198\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8728\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__8728\,
            I => \uu2.mem0.N_77_i\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__8725\,
            I => \uu2.mem0.w_data_i_a3_1_0_cascade_\
        );

    \I__1195\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__8719\,
            I => \uu2.mem0.N_79_i_0\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__1192\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8709\
        );

    \I__1191\ : IoInMux
    port map (
            O => \N__8712\,
            I => \N__8706\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__8709\,
            I => \N__8703\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8706\,
            I => \N__8700\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__8703\,
            I => \N__8697\
        );

    \I__1187\ : Span12Mux_s9_v
    port map (
            O => \N__8700\,
            I => \N__8692\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__8697\,
            I => \N__8692\
        );

    \I__1185\ : Odrv12
    port map (
            O => \N__8692\,
            I => clk
        );

    \I__1184\ : SRMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__1182\ : Span4Mux_s3_h
    port map (
            O => \N__8683\,
            I => \N__8680\
        );

    \I__1181\ : Span4Mux_h
    port map (
            O => \N__8680\,
            I => \N__8676\
        );

    \I__1180\ : CEMux
    port map (
            O => \N__8679\,
            I => \N__8673\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__8676\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__8673\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__8668\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__8665\,
            I => \uu0.un220_ci_cascade_\
        );

    \I__1175\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8658\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8655\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8652\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__8655\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__8652\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1169\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8638\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__8638\,
            I => \uu0.un99_ci_0\
        );

    \I__1166\ : InMux
    port map (
            O => \N__8635\,
            I => \N__8626\
        );

    \I__1165\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8626\
        );

    \I__1164\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8626\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__8626\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__8623\,
            I => \N__8619\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__8622\,
            I => \N__8616\
        );

    \I__1160\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8613\
        );

    \I__1159\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8610\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__8613\,
            I => \N__8607\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8604\
        );

    \I__1156\ : Odrv12
    port map (
            O => \N__8607\,
            I => \uu0.un88_ci_3\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__8604\,
            I => \uu0.un88_ci_3\
        );

    \I__1154\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8585\
        );

    \I__1153\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8578\
        );

    \I__1152\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8578\
        );

    \I__1151\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8578\
        );

    \I__1150\ : InMux
    port map (
            O => \N__8595\,
            I => \N__8569\
        );

    \I__1149\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8569\
        );

    \I__1148\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8569\
        );

    \I__1147\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8569\
        );

    \I__1146\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8566\
        );

    \I__1145\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8559\
        );

    \I__1144\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8559\
        );

    \I__1143\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8559\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8556\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8551\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8551\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__8566\,
            I => \uu0.un4_l_count_0\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8559\,
            I => \uu0.un4_l_count_0\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__8556\,
            I => \uu0.un4_l_count_0\
        );

    \I__1136\ : Odrv4
    port map (
            O => \N__8551\,
            I => \uu0.un4_l_count_0\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8536\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8541\,
            I => \N__8533\
        );

    \I__1133\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8528\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8539\,
            I => \N__8528\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8523\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8523\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__8528\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__8523\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1127\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8511\
        );

    \I__1126\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8508\
        );

    \I__1125\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8501\
        );

    \I__1124\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8501\
        );

    \I__1123\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8501\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__8511\,
            I => \N__8494\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__8508\,
            I => \N__8494\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__8501\,
            I => \N__8494\
        );

    \I__1119\ : Odrv4
    port map (
            O => \N__8494\,
            I => \uu0.un66_ci\
        );

    \I__1118\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8488\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__8488\,
            I => \N__8482\
        );

    \I__1116\ : InMux
    port map (
            O => \N__8487\,
            I => \N__8479\
        );

    \I__1115\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8476\
        );

    \I__1114\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8473\
        );

    \I__1113\ : Span4Mux_h
    port map (
            O => \N__8482\,
            I => \N__8470\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__8479\,
            I => \N__8467\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__8476\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8473\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__8470\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__8467\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1107\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8453\
        );

    \I__1106\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8450\
        );

    \I__1105\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8447\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8442\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__8450\,
            I => \N__8442\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__8447\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__8442\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1100\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8432\
        );

    \I__1099\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8427\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8427\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__8432\,
            I => \uu0.un198_ci_2\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__8427\,
            I => \uu0.un198_ci_2\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__8422\,
            I => \N__8417\
        );

    \I__1094\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8413\
        );

    \I__1093\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8408\
        );

    \I__1092\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8408\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__8416\,
            I => \N__8401\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8396\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8396\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__8407\,
            I => \N__8393\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__8406\,
            I => \N__8390\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__8405\,
            I => \N__8387\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__8404\,
            I => \N__8384\
        );

    \I__1084\ : InMux
    port map (
            O => \N__8401\,
            I => \N__8379\
        );

    \I__1083\ : Span4Mux_s2_h
    port map (
            O => \N__8396\,
            I => \N__8376\
        );

    \I__1082\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8373\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8370\
        );

    \I__1080\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8361\
        );

    \I__1079\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8361\
        );

    \I__1078\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8361\
        );

    \I__1077\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8361\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8358\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__8376\,
            I => \uu0.un110_ci\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__8373\,
            I => \uu0.un110_ci\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__8370\,
            I => \uu0.un110_ci\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__8361\,
            I => \uu0.un110_ci\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__8358\,
            I => \uu0.un110_ci\
        );

    \I__1070\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8344\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__8344\,
            I => \N__8338\
        );

    \I__1068\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8333\
        );

    \I__1067\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8333\
        );

    \I__1066\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8330\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__8338\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__8333\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__8330\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__8323\,
            I => \N__8319\
        );

    \I__1061\ : InMux
    port map (
            O => \N__8322\,
            I => \N__8313\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8313\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8310\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__8313\,
            I => \N__8307\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8310\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1056\ : Odrv4
    port map (
            O => \N__8307\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1055\ : CEMux
    port map (
            O => \N__8302\,
            I => \N__8284\
        );

    \I__1054\ : CEMux
    port map (
            O => \N__8301\,
            I => \N__8284\
        );

    \I__1053\ : CEMux
    port map (
            O => \N__8300\,
            I => \N__8284\
        );

    \I__1052\ : CEMux
    port map (
            O => \N__8299\,
            I => \N__8284\
        );

    \I__1051\ : CEMux
    port map (
            O => \N__8298\,
            I => \N__8284\
        );

    \I__1050\ : CEMux
    port map (
            O => \N__8297\,
            I => \N__8284\
        );

    \I__1049\ : GlobalMux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1048\ : gio2CtrlBuf
    port map (
            O => \N__8281\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__8278\,
            I => \resetGen.escKeyZ0_cascade_\
        );

    \I__1046\ : CascadeMux
    port map (
            O => \N__8275\,
            I => \resetGen.un252_ci_cascade_\
        );

    \I__1045\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__8269\,
            I => \N__8265\
        );

    \I__1043\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8262\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__8265\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__8262\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1040\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8247\
        );

    \I__1039\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8247\
        );

    \I__1038\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8247\
        );

    \I__1037\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8244\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__8247\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__8244\,
            I => \resetGen.reset_countZ0Z_0\
        );

    \I__1034\ : InMux
    port map (
            O => \N__8239\,
            I => \N__8232\
        );

    \I__1033\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8232\
        );

    \I__1032\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8229\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__8232\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__8229\,
            I => \resetGen.reset_countZ0Z_1\
        );

    \I__1029\ : CascadeMux
    port map (
            O => \N__8224\,
            I => \N__8221\
        );

    \I__1028\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8214\
        );

    \I__1027\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8214\
        );

    \I__1026\ : InMux
    port map (
            O => \N__8219\,
            I => \N__8211\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__8214\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__8211\,
            I => \resetGen.reset_countZ0Z_2\
        );

    \I__1023\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__1022\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8200\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__8200\,
            I => \N__8197\
        );

    \I__1020\ : Odrv12
    port map (
            O => \N__8197\,
            I => \resetGen.un241_ci\
        );

    \I__1019\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8191\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__8191\,
            I => \resetGen.reset_count_2_0_4\
        );

    \I__1017\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8176\
        );

    \I__1016\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8176\
        );

    \I__1015\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8176\
        );

    \I__1014\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8176\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__8176\,
            I => \resetGen.escKeyZ0\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__8172\,
            I => \N__8164\
        );

    \I__1010\ : InMux
    port map (
            O => \N__8171\,
            I => \N__8154\
        );

    \I__1009\ : InMux
    port map (
            O => \N__8170\,
            I => \N__8154\
        );

    \I__1008\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8154\
        );

    \I__1007\ : InMux
    port map (
            O => \N__8164\,
            I => \N__8154\
        );

    \I__1006\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8151\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__8154\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__8151\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1003\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8139\
        );

    \I__1002\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8139\
        );

    \I__1001\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8136\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__8139\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__8136\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__998\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__8128\,
            I => \N__8125\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__8125\,
            I => \uu0.un4_l_count_12\
        );

    \I__995\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8118\
        );

    \I__994\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8115\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__8118\,
            I => \N__8107\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8107\
        );

    \I__991\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8100\
        );

    \I__990\ : InMux
    port map (
            O => \N__8113\,
            I => \N__8100\
        );

    \I__989\ : InMux
    port map (
            O => \N__8112\,
            I => \N__8100\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__8107\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__8100\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__986\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8090\
        );

    \I__985\ : InMux
    port map (
            O => \N__8094\,
            I => \N__8087\
        );

    \I__984\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8084\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8081\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__8087\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__8084\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__8081\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__979\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8067\
        );

    \I__978\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8067\
        );

    \I__977\ : InMux
    port map (
            O => \N__8072\,
            I => \N__8064\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8061\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__8064\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__974\ : Odrv4
    port map (
            O => \N__8061\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__973\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__8050\,
            I => vbuf_tx_data_6
        );

    \I__970\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8044\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__8044\,
            I => \N__8041\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__8041\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__967\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8032\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__8032\,
            I => vbuf_tx_data_7
        );

    \I__964\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8026\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__8026\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__962\ : CEMux
    port map (
            O => \N__8023\,
            I => \N__8019\
        );

    \I__961\ : CEMux
    port map (
            O => \N__8022\,
            I => \N__8016\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__8019\,
            I => \N__8013\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__8016\,
            I => \N__8010\
        );

    \I__958\ : Span4Mux_v
    port map (
            O => \N__8013\,
            I => \N__8006\
        );

    \I__957\ : Span4Mux_v
    port map (
            O => \N__8010\,
            I => \N__8003\
        );

    \I__956\ : CEMux
    port map (
            O => \N__8009\,
            I => \N__8000\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__8006\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__8003\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__8000\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__7993\,
            I => \uu0.un88_ci_3_cascade_\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__7990\,
            I => \N__7978\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7975\
        );

    \I__949\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7958\
        );

    \I__948\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7958\
        );

    \I__947\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7958\
        );

    \I__946\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7958\
        );

    \I__945\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7958\
        );

    \I__944\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7958\
        );

    \I__943\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7953\
        );

    \I__942\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7953\
        );

    \I__941\ : InMux
    port map (
            O => \N__7978\,
            I => \N__7942\
        );

    \I__940\ : InMux
    port map (
            O => \N__7975\,
            I => \N__7942\
        );

    \I__939\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7942\
        );

    \I__938\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7942\
        );

    \I__937\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7942\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__7971\,
            I => \N__7939\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7930\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7930\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7942\,
            I => \N__7930\
        );

    \I__932\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7927\
        );

    \I__931\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7922\
        );

    \I__930\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7922\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__7930\,
            I => \N__7919\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__7927\,
            I => vbuf_tx_data_rdy
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7922\,
            I => vbuf_tx_data_rdy
        );

    \I__926\ : Odrv4
    port map (
            O => \N__7919\,
            I => vbuf_tx_data_rdy
        );

    \I__925\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7909\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__7906\,
            I => \uu2.r_data_wire_2\
        );

    \I__922\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__7900\,
            I => vbuf_tx_data_2
        );

    \I__920\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__7891\,
            I => \uu2.r_data_wire_3\
        );

    \I__917\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7885\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__7885\,
            I => vbuf_tx_data_3
        );

    \I__915\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7879\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7879\,
            I => \uu2.r_data_wire_4\
        );

    \I__913\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__7873\,
            I => vbuf_tx_data_4
        );

    \I__911\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7867\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__7867\,
            I => \uu2.r_data_wire_5\
        );

    \I__909\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7861\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__7861\,
            I => vbuf_tx_data_5
        );

    \I__907\ : InMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__7855\,
            I => \uu2.r_data_wire_6\
        );

    \I__905\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__7849\,
            I => \uu2.r_data_wire_7\
        );

    \I__903\ : CEMux
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__901\ : Span4Mux_v
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__7837\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__899\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7831\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__7831\,
            I => \uu0.sec_clkDZ0\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__7828\,
            I => \uu2.un1_l_count_2_2_cascade_\
        );

    \I__896\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7822\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__7822\,
            I => \uu2.un284_ci\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__893\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7809\
        );

    \I__892\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7809\
        );

    \I__891\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7806\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__7809\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__7806\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__7801\,
            I => \N__7798\
        );

    \I__887\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7793\
        );

    \I__886\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7790\
        );

    \I__885\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7787\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__7793\,
            I => \N__7784\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__7790\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__7787\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__7784\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__880\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7772\
        );

    \I__879\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7767\
        );

    \I__878\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7767\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__7772\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7767\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__875\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7753\
        );

    \I__874\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7753\
        );

    \I__873\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7748\
        );

    \I__872\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7748\
        );

    \I__871\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7745\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__7753\,
            I => \N__7742\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__7748\,
            I => \N__7739\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__7745\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__867\ : Odrv4
    port map (
            O => \N__7742\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__7739\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__7732\,
            I => \N__7727\
        );

    \I__864\ : CascadeMux
    port map (
            O => \N__7731\,
            I => \N__7724\
        );

    \I__863\ : InMux
    port map (
            O => \N__7730\,
            I => \N__7717\
        );

    \I__862\ : InMux
    port map (
            O => \N__7727\,
            I => \N__7717\
        );

    \I__861\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7717\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__7717\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__859\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7700\
        );

    \I__858\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7700\
        );

    \I__857\ : InMux
    port map (
            O => \N__7712\,
            I => \N__7700\
        );

    \I__856\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7700\
        );

    \I__855\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7695\
        );

    \I__854\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7695\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__7700\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7695\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__851\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7680\
        );

    \I__850\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7680\
        );

    \I__849\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7680\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__7687\,
            I => \N__7676\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__7680\,
            I => \N__7673\
        );

    \I__846\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7668\
        );

    \I__845\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7668\
        );

    \I__844\ : Odrv4
    port map (
            O => \N__7673\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__7668\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__842\ : InMux
    port map (
            O => \N__7663\,
            I => \N__7654\
        );

    \I__841\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7654\
        );

    \I__840\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7647\
        );

    \I__839\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7647\
        );

    \I__838\ : InMux
    port map (
            O => \N__7659\,
            I => \N__7647\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__7654\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__7647\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__7642\,
            I => \uu2.un1_l_count_1_2_0_cascade_\
        );

    \I__834\ : InMux
    port map (
            O => \N__7639\,
            I => \N__7633\
        );

    \I__833\ : InMux
    port map (
            O => \N__7638\,
            I => \N__7633\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__7633\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__7630\,
            I => \N__7624\
        );

    \I__830\ : InMux
    port map (
            O => \N__7629\,
            I => \N__7619\
        );

    \I__829\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7619\
        );

    \I__828\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7616\
        );

    \I__827\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7613\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__7619\,
            I => \N__7610\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__7616\,
            I => \uu2.un306_ci\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__7613\,
            I => \uu2.un306_ci\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__7610\,
            I => \uu2.un306_ci\
        );

    \I__822\ : InMux
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__7597\,
            I => \uu2.r_data_wire_0\
        );

    \I__819\ : InMux
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__7591\,
            I => vbuf_tx_data_0
        );

    \I__817\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7582\
        );

    \I__815\ : Odrv4
    port map (
            O => \N__7582\,
            I => \uu2.r_data_wire_1\
        );

    \I__814\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7576\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7576\,
            I => vbuf_tx_data_1
        );

    \I__812\ : InMux
    port map (
            O => \N__7573\,
            I => \N__7564\
        );

    \I__811\ : InMux
    port map (
            O => \N__7572\,
            I => \N__7564\
        );

    \I__810\ : InMux
    port map (
            O => \N__7571\,
            I => \N__7557\
        );

    \I__809\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7557\
        );

    \I__808\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7557\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__7564\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__7557\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__805\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__7549\,
            I => \buart.Z_tx.un1_bitcount_c3\
        );

    \I__803\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7542\
        );

    \I__802\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7539\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__7542\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__7539\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__799\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7521\
        );

    \I__798\ : InMux
    port map (
            O => \N__7533\,
            I => \N__7521\
        );

    \I__797\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7521\
        );

    \I__796\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7521\
        );

    \I__795\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7518\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__7521\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__7518\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__792\ : InMux
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7510\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__7507\,
            I => \N__7503\
        );

    \I__789\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7495\
        );

    \I__788\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7495\
        );

    \I__787\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7495\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__7495\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__784\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7486\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__7486\,
            I => \uu2.un350_ci\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__7483\,
            I => \N__7479\
        );

    \I__781\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7474\
        );

    \I__780\ : InMux
    port map (
            O => \N__7479\,
            I => \N__7474\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__7474\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__778\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7465\
        );

    \I__777\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7465\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__7465\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__775\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7456\
        );

    \I__774\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7456\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__7456\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__7453\,
            I => \N__7449\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__7452\,
            I => \N__7446\
        );

    \I__770\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7441\
        );

    \I__769\ : InMux
    port map (
            O => \N__7446\,
            I => \N__7441\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__7441\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__766\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7429\
        );

    \I__765\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7429\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__7429\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__763\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7423\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__7423\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__7420\,
            I => \N__7416\
        );

    \I__760\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7412\
        );

    \I__759\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7407\
        );

    \I__758\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7407\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__7412\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7407\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__755\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7394\
        );

    \I__754\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7394\
        );

    \I__753\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7389\
        );

    \I__752\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7389\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__7394\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__7389\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__7384\,
            I => \buart.Z_tx.uart_busy_0_0_cascade_\
        );

    \I__748\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7371\
        );

    \I__747\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7371\
        );

    \I__746\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7371\
        );

    \I__745\ : InMux
    port map (
            O => \N__7378\,
            I => \N__7368\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__7371\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__7368\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__7363\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__741\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7354\
        );

    \I__740\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7347\
        );

    \I__739\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7347\
        );

    \I__738\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7347\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__7354\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__7347\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__735\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7334\
        );

    \I__734\ : InMux
    port map (
            O => \N__7341\,
            I => \N__7334\
        );

    \I__733\ : InMux
    port map (
            O => \N__7340\,
            I => \N__7329\
        );

    \I__732\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7329\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__7334\,
            I => \uu0.un154_ci_9\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__7329\,
            I => \uu0.un154_ci_9\
        );

    \I__729\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7319\
        );

    \I__728\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7314\
        );

    \I__727\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7314\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__7319\,
            I => \N__7311\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__7314\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__7311\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__7306\,
            I => \uu0.un4_l_count_0_8_cascade_\
        );

    \I__722\ : CascadeMux
    port map (
            O => \N__7303\,
            I => \N__7297\
        );

    \I__721\ : InMux
    port map (
            O => \N__7302\,
            I => \N__7292\
        );

    \I__720\ : InMux
    port map (
            O => \N__7301\,
            I => \N__7292\
        );

    \I__719\ : InMux
    port map (
            O => \N__7300\,
            I => \N__7287\
        );

    \I__718\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7287\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7292\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__7287\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__715\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7269\
        );

    \I__714\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7269\
        );

    \I__713\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7269\
        );

    \I__712\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7269\
        );

    \I__711\ : InMux
    port map (
            O => \N__7278\,
            I => \N__7266\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__7269\,
            I => \N__7263\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__7266\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__708\ : Odrv12
    port map (
            O => \N__7263\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__707\ : InMux
    port map (
            O => \N__7258\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__706\ : InMux
    port map (
            O => \N__7255\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__705\ : InMux
    port map (
            O => \N__7252\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__704\ : InMux
    port map (
            O => \N__7249\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__703\ : InMux
    port map (
            O => \N__7246\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__702\ : InMux
    port map (
            O => \N__7243\,
            I => \N__7231\
        );

    \I__701\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7231\
        );

    \I__700\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7231\
        );

    \I__699\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7231\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__7231\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__697\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7225\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__7225\,
            I => \uu0.un143_ci_0\
        );

    \I__695\ : InMux
    port map (
            O => \N__7222\,
            I => \N__7204\
        );

    \I__694\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7204\
        );

    \I__693\ : InMux
    port map (
            O => \N__7220\,
            I => \N__7204\
        );

    \I__692\ : InMux
    port map (
            O => \N__7219\,
            I => \N__7204\
        );

    \I__691\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7204\
        );

    \I__690\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7204\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__7204\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__7201\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__7198\,
            I => \N__7195\
        );

    \I__686\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7192\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__7192\,
            I => \uu0.un165_ci_0\
        );

    \I__684\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7185\
        );

    \I__683\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7182\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__7185\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__7182\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__680\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7168\
        );

    \I__679\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7168\
        );

    \I__678\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7168\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__7168\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__676\ : InMux
    port map (
            O => \N__7165\,
            I => \N__7160\
        );

    \I__675\ : InMux
    port map (
            O => \N__7164\,
            I => \N__7155\
        );

    \I__674\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7155\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__7160\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__7155\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__7150\,
            I => \uu0.un55_ci_cascade_\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \N__7140\
        );

    \I__669\ : InMux
    port map (
            O => \N__7146\,
            I => \N__7126\
        );

    \I__668\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7126\
        );

    \I__667\ : InMux
    port map (
            O => \N__7144\,
            I => \N__7126\
        );

    \I__666\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7126\
        );

    \I__665\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7126\
        );

    \I__664\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7126\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__7126\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__662\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7110\
        );

    \I__661\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7110\
        );

    \I__660\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7110\
        );

    \I__659\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7110\
        );

    \I__658\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7107\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__7110\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__7107\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__7102\,
            I => \N__7098\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__7101\,
            I => \N__7095\
        );

    \I__653\ : InMux
    port map (
            O => \N__7098\,
            I => \N__7086\
        );

    \I__652\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7086\
        );

    \I__651\ : InMux
    port map (
            O => \N__7094\,
            I => \N__7086\
        );

    \I__650\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7083\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__7086\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__7083\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__7078\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__646\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__7069\,
            I => \uu0.un4_l_count_18\
        );

    \I__643\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7061\
        );

    \I__642\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7058\
        );

    \I__641\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7055\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__7061\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__7058\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__7055\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__7048\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \N__7040\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__7044\,
            I => \N__7037\
        );

    \I__634\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7030\
        );

    \I__633\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7030\
        );

    \I__632\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7030\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__7030\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__7027\,
            I => \uu0.un4_l_count_11_cascade_\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__7024\,
            I => \uu0.un4_l_count_16_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__7021\,
            I => \N__7017\
        );

    \I__627\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7014\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__7017\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__7014\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__623\ : InMux
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__7003\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__621\ : IoInMux
    port map (
            O => \N__7000\,
            I => \N__6997\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__6997\,
            I => \uu0.un11_l_count_i\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__618\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6981\
        );

    \I__617\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6981\
        );

    \I__616\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6981\
        );

    \I__615\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6978\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__6981\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__6978\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__612\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6970\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__6970\,
            I => \uu0.un4_l_count_13\
        );

    \I__610\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6964\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__608\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__6958\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__606\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6952\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6952\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__6949\,
            I => \uu2.un284_ci_cascade_\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__6946\,
            I => \uu2.un306_ci_cascade_\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__601\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6937\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6934\
        );

    \I__599\ : Odrv4
    port map (
            O => \N__6934\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__598\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__6928\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__596\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__6922\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__594\ : InMux
    port map (
            O => \N__6919\,
            I => \N__6916\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__6916\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__592\ : IoInMux
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__590\ : IoSpan4Mux
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__589\ : Odrv4
    port map (
            O => \N__6904\,
            I => o_serial_data_c
        );

    \I__588\ : IoInMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__6898\,
            I => \N__6895\
        );

    \I__586\ : Span12Mux_s5_h
    port map (
            O => \N__6895\,
            I => \N__6892\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__6889\,
            I => clk_in_c
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__18050\
        );

    \INVuu2.w_addr_displaying_nesr_5C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_5C_net\,
            I => \N__18056\
        );

    \INVuu2.bitmap_215C\ : INV
    port map (
            O => \INVuu2.bitmap_215C_net\,
            I => \N__18044\
        );

    \INVuu2.w_addr_displaying_nesr_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_8C_net\,
            I => \N__18055\
        );

    \INVuu2.w_addr_user_nesr_3C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_3C_net\,
            I => \N__18067\
        );

    \INVuu2.bitmap_168C\ : INV
    port map (
            O => \INVuu2.bitmap_168C_net\,
            I => \N__18024\
        );

    \INVuu2.bitmap_200C\ : INV
    port map (
            O => \INVuu2.bitmap_200C_net\,
            I => \N__18029\
        );

    \INVuu2.w_addr_displaying_fast_nesr_8C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            I => \N__18033\
        );

    \INVuu2.w_addr_displaying_2_rep1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_2_rep1C_net\,
            I => \N__18040\
        );

    \INVuu2.w_addr_displaying_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4C_net\,
            I => \N__18052\
        );

    \INVuu2.w_addr_user_nesr_6C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_6C_net\,
            I => \N__18058\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__18031\
        );

    \INVuu2.bitmap_290C\ : INV
    port map (
            O => \INVuu2.bitmap_290C_net\,
            I => \N__18036\
        );

    \INVuu2.bitmap_197C\ : INV
    port map (
            O => \INVuu2.bitmap_197C_net\,
            I => \N__18061\
        );

    \INVuu2.bitmap_308C\ : INV
    port map (
            O => \INVuu2.bitmap_308C_net\,
            I => \N__18035\
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__18043\
        );

    \INVuu2.bitmap_186C\ : INV
    port map (
            O => \INVuu2.bitmap_186C_net\,
            I => \N__18049\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__18072\
        );

    \IN_MUX_bfv_2_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_3_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8712\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7000\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__17647\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \buart.Z_tx.shifter_0_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__7982\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18094\,
            ce => \N__8009\,
            sr => \N__17820\
        );

    \buart.Z_tx.uart_tx_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7981\,
            in2 => \_gnd_net_\,
            in3 => \N__6919\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18094\,
            ce => \N__8009\,
            sr => \N__17820\
        );

    \uu2.l_count_7_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__8074\,
            in1 => \N__7762\,
            in2 => \N__7630\,
            in3 => \N__7816\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18088\,
            ce => 'H',
            sr => \N__17817\
        );

    \uu2.l_count_1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7714\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18088\,
            ce => 'H',
            sr => \N__17817\
        );

    \uu2.l_count_0_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__7713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18088\,
            ce => 'H',
            sr => \N__17817\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7660\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7712\,
            lcout => \uu2.un284_ci\,
            ltout => \uu2.un284_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_2_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6949\,
            in3 => \N__7679\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18088\,
            ce => 'H',
            sr => \N__17817\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7659\,
            in1 => \N__7711\,
            in2 => \N__7687\,
            in3 => \N__7777\,
            lcout => \uu2.un306_ci\,
            ltout => \uu2.un306_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8073\,
            in1 => \N__7761\,
            in2 => \N__6946\,
            in3 => \N__7815\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_8_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6943\,
            in3 => \N__7796\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18088\,
            ce => 'H',
            sr => \N__17817\
        );

    \buart.Z_tx.shifter_1_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7983\,
            in1 => \N__6931\,
            in2 => \_gnd_net_\,
            in3 => \N__7594\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \buart.Z_tx.shifter_2_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__6925\,
            in1 => \N__7986\,
            in2 => \_gnd_net_\,
            in3 => \N__7579\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \buart.Z_tx.shifter_3_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7984\,
            in1 => \N__6967\,
            in2 => \_gnd_net_\,
            in3 => \N__7903\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \buart.Z_tx.shifter_4_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7888\,
            in1 => \N__6961\,
            in2 => \_gnd_net_\,
            in3 => \N__7988\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \buart.Z_tx.shifter_5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__6955\,
            in2 => \_gnd_net_\,
            in3 => \N__7876\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \buart.Z_tx.shifter_6_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__8047\,
            in1 => \N__7987\,
            in2 => \_gnd_net_\,
            in3 => \N__7864\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18078\,
            ce => \N__8022\,
            sr => \N__17814\
        );

    \uu2.l_count_5_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__8094\,
            in1 => \N__8122\,
            in2 => \_gnd_net_\,
            in3 => \N__7629\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \uu2.l_count_6_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7628\,
            in1 => \N__8072\,
            in2 => \_gnd_net_\,
            in3 => \N__7758\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \Lab_UT.dispString.cnt_1_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__15290\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15206\,
            lcout => \Lab_UT.cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \Lab_UT.dispString.cnt_0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15289\,
            lcout => \Lab_UT.cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \uu0.sec_clk_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9195\,
            in2 => \_gnd_net_\,
            in3 => \N__8591\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \uu0.delay_line_1_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7021\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18071\,
            ce => 'H',
            sr => \N__17805\
        );

    \uu0.delay_line_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7280\,
            in1 => \N__9101\,
            in2 => \N__7045\,
            in3 => \N__6991\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18065\,
            ce => 'H',
            sr => \N__17815\
        );

    \uu0.l_precount_3_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__6993\,
            in1 => \N__7043\,
            in2 => \N__9106\,
            in3 => \N__7282\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18065\,
            ce => 'H',
            sr => \N__17815\
        );

    \uu0.l_precount_2_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__7281\,
            in1 => \N__9102\,
            in2 => \_gnd_net_\,
            in3 => \N__6992\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18065\,
            ce => 'H',
            sr => \N__17815\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7279\,
            in1 => \N__8457\,
            in2 => \N__7044\,
            in3 => \N__7119\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI96A32_18_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7324\,
            in1 => \N__8662\,
            in2 => \N__7027\,
            in3 => \N__8541\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_11_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6973\,
            in1 => \N__8131\,
            in2 => \N__7024\,
            in3 => \N__7075\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_RNILLLG7_1_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111010"
        )
    port map (
            in0 => \N__7020\,
            in1 => \_gnd_net_\,
            in2 => \N__7009\,
            in3 => \N__7006\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2CNU_11_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8341\,
            in1 => \N__7064\,
            in2 => \N__6994\,
            in3 => \N__7139\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8145\,
            in1 => \N__7094\,
            in2 => \N__7147\,
            in3 => \N__7120\,
            lcout => \uu0.un66_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__7123\,
            in1 => \_gnd_net_\,
            in2 => \N__7102\,
            in3 => \N__7146\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18059\,
            ce => \N__8297\,
            sr => \N__17816\
        );

    \uu0.l_count_0_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7144\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18059\,
            ce => \N__8297\,
            sr => \N__17816\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7121\,
            in1 => \_gnd_net_\,
            in2 => \N__7101\,
            in3 => \N__7143\,
            lcout => OPEN,
            ltout => \uu0.un55_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_3_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__8146\,
            in1 => \_gnd_net_\,
            in2 => \N__7150\,
            in3 => \N__8590\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18059\,
            ce => \N__8297\,
            sr => \N__17816\
        );

    \uu0.l_count_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7122\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7145\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18059\,
            ce => \N__8297\,
            sr => \N__17816\
        );

    \uu0.l_count_11_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__7228\,
            in1 => \N__7066\,
            in2 => \N__8407\,
            in3 => \N__8589\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18059\,
            ce => \N__8297\,
            sr => \N__17816\
        );

    \uu0.l_count_RNI04591_10_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7240\,
            in1 => \N__7217\,
            in2 => \N__7303\,
            in3 => \N__7093\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI2GS72_4_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9099\,
            in1 => \N__8487\,
            in2 => \N__7078\,
            in3 => \N__7163\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7241\,
            in1 => \N__7065\,
            in2 => \N__8172\,
            in3 => \N__7218\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_14_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8382\,
            in1 => \N__7300\,
            in2 => \N__7048\,
            in3 => \N__7164\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18053\,
            ce => \N__8298\,
            sr => \N__17819\
        );

    \uu0.l_count_8_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8383\,
            in2 => \_gnd_net_\,
            in3 => \N__7221\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18053\,
            ce => \N__8298\,
            sr => \N__17819\
        );

    \uu0.l_count_10_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__7220\,
            in1 => \N__8170\,
            in2 => \N__8405\,
            in3 => \N__7243\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18053\,
            ce => \N__8298\,
            sr => \N__17819\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7242\,
            in1 => \_gnd_net_\,
            in2 => \N__8173\,
            in3 => \N__7219\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_9_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__7222\,
            in1 => \_gnd_net_\,
            in2 => \N__8404\,
            in3 => \N__8171\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18053\,
            ce => \N__8298\,
            sr => \N__17819\
        );

    \uu0.l_count_13_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__8597\,
            in1 => \N__7189\,
            in2 => \N__7198\,
            in3 => \N__8420\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18047\,
            ce => \N__8299\,
            sr => \N__17822\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7302\,
            in1 => \N__7340\,
            in2 => \_gnd_net_\,
            in3 => \N__7165\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8421\,
            in1 => \N__8599\,
            in2 => \N__7201\,
            in3 => \N__7323\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18047\,
            ce => \N__8299\,
            sr => \N__17822\
        );

    \uu0.l_count_12_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7342\,
            in1 => \N__8596\,
            in2 => \N__8422\,
            in3 => \N__7177\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18047\,
            ce => \N__8299\,
            sr => \N__17822\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7341\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIFAQ9_13_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7188\,
            in2 => \_gnd_net_\,
            in3 => \N__7175\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => \uu0.un4_l_count_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7339\,
            in1 => \N__7322\,
            in2 => \N__7306\,
            in3 => \N__7301\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_4_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8517\,
            in1 => \N__8598\,
            in2 => \_gnd_net_\,
            in3 => \N__8485\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18047\,
            ce => \N__8299\,
            sr => \N__17822\
        );

    \uu0.l_precount_1_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9100\,
            in2 => \_gnd_net_\,
            in3 => \N__7278\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18041\,
            ce => 'H',
            sr => \N__17824\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7400\,
            in2 => \N__7420\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_3_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7482\,
            in2 => \_gnd_net_\,
            in3 => \N__7258\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__18097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__7380\,
            in1 => \_gnd_net_\,
            in2 => \N__7438\,
            in3 => \N__7255\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__18097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7462\,
            in2 => \_gnd_net_\,
            in3 => \N__7252\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__18097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7381\,
            in1 => \N__7471\,
            in2 => \_gnd_net_\,
            in3 => \N__7249\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__18097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7379\,
            in2 => \N__7453\,
            in3 => \N__7246\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7415\,
            in1 => \N__7399\,
            in2 => \N__7483\,
            in3 => \N__7426\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7470\,
            in1 => \N__7461\,
            in2 => \N__7452\,
            in3 => \N__7434\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7419\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7401\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18095\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000111110000"
        )
    port map (
            in0 => \N__7570\,
            in1 => \N__7358\,
            in2 => \N__7507\,
            in3 => \N__7530\,
            lcout => \buart.Z_tx.bitcount_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7569\,
            in2 => \_gnd_net_\,
            in3 => \N__7545\,
            lcout => OPEN,
            ltout => \buart.Z_tx.uart_busy_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__7502\,
            in1 => \N__7357\,
            in2 => \N__7384\,
            in3 => \N__7378\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__7359\,
            in1 => \N__7571\,
            in2 => \N__7363\,
            in3 => \N__7506\,
            lcout => \buart.Z_tx.un1_bitcount_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111110010"
        )
    port map (
            in0 => \N__7533\,
            in1 => \N__7573\,
            in2 => \N__7989\,
            in3 => \N__7360\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \buart.Z_tx.bitcount_0_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__7572\,
            in1 => \N__7974\,
            in2 => \_gnd_net_\,
            in3 => \N__7532\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \buart.Z_tx.bitcount_3_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100111110110"
        )
    port map (
            in0 => \N__7534\,
            in1 => \N__7546\,
            in2 => \N__7990\,
            in3 => \N__7552\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7972\,
            in2 => \_gnd_net_\,
            in3 => \N__7531\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7513\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \uu2.r_addr_2_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9328\,
            in1 => \N__9371\,
            in2 => \N__8794\,
            in3 => \N__9256\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \uu2.r_addr_1_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__9255\,
            in1 => \N__8790\,
            in2 => \_gnd_net_\,
            in3 => \N__9327\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \uu2.r_addr_0_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8789\,
            in2 => \_gnd_net_\,
            in3 => \N__9254\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18089\,
            ce => 'H',
            sr => \N__17806\
        );

    \uu2.l_count_9_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__8754\,
            in1 => \N__7730\,
            in2 => \N__7492\,
            in3 => \N__7797\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18079\,
            ce => 'H',
            sr => \N__17821\
        );

    \uu2.l_count_RNIBCGK1_9_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7760\,
            in1 => \N__8113\,
            in2 => \N__7732\,
            in3 => \N__7710\,
            lcout => OPEN,
            ltout => \uu2.un1_l_count_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7689\,
            in1 => \N__7663\,
            in2 => \N__7828\,
            in3 => \N__7638\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_3_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__7776\,
            in1 => \N__7825\,
            in2 => \N__7819\,
            in3 => \N__7690\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18079\,
            ce => 'H',
            sr => \N__17821\
        );

    \uu2.l_count_RNIFGGK1_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7814\,
            in1 => \N__8095\,
            in2 => \N__7801\,
            in3 => \N__7775\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7759\,
            in1 => \N__8112\,
            in2 => \N__7731\,
            in3 => \N__7709\,
            lcout => OPEN,
            ltout => \uu2.un1_l_count_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_0_1_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7688\,
            in1 => \N__7662\,
            in2 => \N__7642\,
            in3 => \N__7639\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7627\,
            in1 => \N__8114\,
            in2 => \_gnd_net_\,
            in3 => \N__8753\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18079\,
            ce => 'H',
            sr => \N__17821\
        );

    \uu2.r_data_reg_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7588\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7912\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7897\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7882\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7858\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7852\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__7846\,
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__9118\,
            in1 => \N__9136\,
            in2 => \_gnd_net_\,
            in3 => \N__17852\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9194\,
            lcout => \uu0.sec_clkDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18066\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7834\,
            in2 => \_gnd_net_\,
            in3 => \N__9193\,
            lcout => \oneSecStrb_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8121\,
            in2 => \_gnd_net_\,
            in3 => \N__8093\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_7_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7937\,
            in1 => \N__8029\,
            in2 => \_gnd_net_\,
            in3 => \N__8056\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18060\,
            ce => \N__8023\,
            sr => \N__17818\
        );

    \buart.Z_tx.shifter_8_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7938\,
            in2 => \_gnd_net_\,
            in3 => \N__8038\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18060\,
            ce => \N__8023\,
            sr => \N__17818\
        );

    \resetGen.reset_count_RNO_0_4_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8219\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8268\,
            lcout => \resetGen.reset_count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8237\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8254\,
            lcout => \resetGen.un241_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8491\,
            in2 => \_gnd_net_\,
            in3 => \N__8458\,
            lcout => \uu0.un88_ci_3\,
            ltout => \uu0.un88_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7993\,
            in3 => \N__8542\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__9172\,
            in1 => \N__8829\,
            in2 => \N__7971\,
            in3 => \N__17855\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10297\,
            in1 => \N__11809\,
            in2 => \_gnd_net_\,
            in3 => \N__14017\,
            lcout => \resetGen.escKeyZ0\,
            ltout => \resetGen.escKeyZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__8256\,
            in1 => \_gnd_net_\,
            in2 => \N__8278\,
            in3 => \N__13937\,
            lcout => \resetGen.reset_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8238\,
            in1 => \N__8255\,
            in2 => \_gnd_net_\,
            in3 => \N__8220\,
            lcout => OPEN,
            ltout => \resetGen.un252_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010100"
        )
    port map (
            in0 => \N__8187\,
            in1 => \N__8272\,
            in2 => \N__8275\,
            in3 => \N__13939\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010100110"
        )
    port map (
            in0 => \N__8239\,
            in1 => \N__8257\,
            in2 => \N__13947\,
            in3 => \N__8185\,
            lcout => \resetGen.reset_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__8186\,
            in1 => \N__13938\,
            in2 => \N__8224\,
            in3 => \N__8205\,
            lcout => \resetGen.reset_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__8206\,
            in1 => \N__8194\,
            in2 => \N__13946\,
            in3 => \N__8188\,
            lcout => \resetGen.reset_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8163\,
            in1 => \N__8633\,
            in2 => \N__8323\,
            in3 => \N__8144\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__8436\,
            in1 => \N__8593\,
            in2 => \N__8406\,
            in3 => \N__8343\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18048\,
            ce => \N__8300\,
            sr => \N__17823\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8514\,
            in1 => \N__8539\,
            in2 => \N__8622\,
            in3 => \N__8634\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8435\,
            in1 => \N__8322\,
            in2 => \N__8668\,
            in3 => \N__8342\,
            lcout => OPEN,
            ltout => \uu0.un220_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_18_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__8592\,
            in1 => \_gnd_net_\,
            in2 => \N__8665\,
            in3 => \N__8661\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18048\,
            ce => \N__8300\,
            sr => \N__17823\
        );

    \uu0.l_count_7_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8635\,
            in1 => \N__8516\,
            in2 => \N__8647\,
            in3 => \N__8595\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18048\,
            ce => \N__8300\,
            sr => \N__17823\
        );

    \uu0.l_count_6_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__8540\,
            in1 => \N__8515\,
            in2 => \N__8623\,
            in3 => \N__8594\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18048\,
            ce => \N__8300\,
            sr => \N__17823\
        );

    \uu0.l_count_5_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__8518\,
            in1 => \N__8486\,
            in2 => \_gnd_net_\,
            in3 => \N__8456\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18042\,
            ce => \N__8301\,
            sr => \N__17825\
        );

    \uu0.l_count_17_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__8437\,
            in1 => \N__8318\,
            in2 => \N__8416\,
            in3 => \N__8347\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18034\,
            ce => \N__8302\,
            sr => \N__17826\
        );

    \CONSTANT_ONE_LUT4_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_5_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9219\,
            in1 => \N__9522\,
            in2 => \N__8788\,
            in3 => \N__9488\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18082\,
            ce => 'H',
            sr => \N__17807\
        );

    \uu2.r_addr_4_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__9521\,
            in1 => \N__8776\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18082\,
            ce => 'H',
            sr => \N__17807\
        );

    \uu2.trig_rd_det_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9157\,
            in2 => \_gnd_net_\,
            in3 => \N__8830\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18082\,
            ce => 'H',
            sr => \N__17807\
        );

    \uu2.trig_rd_det_1_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8803\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18082\,
            ce => 'H',
            sr => \N__17807\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8809\,
            in2 => \_gnd_net_\,
            in3 => \N__8802\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => \uu2.trig_rd_is_det_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8758\,
            in3 => \N__17854\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9158\,
            in2 => \_gnd_net_\,
            in3 => \N__8755\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18082\,
            ce => 'H',
            sr => \N__17807\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10686\,
            in1 => \N__12322\,
            in2 => \_gnd_net_\,
            in3 => \N__13071\,
            lcout => \uu2.mem0.N_77_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_21_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14706\,
            in1 => \N__14995\,
            in2 => \_gnd_net_\,
            in3 => \N__12378\,
            lcout => OPEN,
            ltout => \uu2.mem0.w_data_i_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100010001"
        )
    port map (
            in0 => \N__12412\,
            in1 => \N__8878\,
            in2 => \N__8725\,
            in3 => \N__12466\,
            lcout => \uu2.mem0.N_79_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__12439\,
            in1 => \N__12409\,
            in2 => \N__8716\,
            in3 => \N__12379\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12323\,
            in1 => \N__11938\,
            in2 => \_gnd_net_\,
            in3 => \N__13628\,
            lcout => \uu2.mem0.N_75_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIUGNM6_2_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10908\,
            in2 => \_gnd_net_\,
            in3 => \N__10955\,
            lcout => \uu2.N_361\,
            ltout => \uu2.N_361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100001101"
        )
    port map (
            in0 => \N__12411\,
            in1 => \N__8854\,
            in2 => \N__8872\,
            in3 => \N__14659\,
            lcout => \uu2.mem0.w_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__14707\,
            in1 => \N__10633\,
            in2 => \_gnd_net_\,
            in3 => \N__12410\,
            lcout => \uu2.mem0.N_69_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14685\,
            in1 => \N__14733\,
            in2 => \N__12435\,
            in3 => \N__14790\,
            lcout => \uu2.mem0.w_data_0_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIFOBB3_8_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13317\,
            in1 => \N__10884\,
            in2 => \N__13627\,
            in3 => \N__13829\,
            lcout => \uu2.N_61\,
            ltout => \uu2.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10909\,
            in2 => \N__8848\,
            in3 => \N__10956\,
            lcout => OPEN,
            ltout => \uu2.mem0.un51_w_data_displaying_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__14734\,
            in1 => \_gnd_net_\,
            in2 => \N__8845\,
            in3 => \N__12344\,
            lcout => \uu2.mem0.w_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__14686\,
            in1 => \N__12239\,
            in2 => \N__12349\,
            in3 => \N__10957\,
            lcout => \uu2.mem0.w_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10009\,
            in1 => \N__12339\,
            in2 => \_gnd_net_\,
            in3 => \N__13507\,
            lcout => \uu2.mem0.N_71_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__13084\,
            in1 => \N__14991\,
            in2 => \N__12348\,
            in3 => \N__9604\,
            lcout => \uu2.mem0.w_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12343\,
            in1 => \N__11884\,
            in2 => \_gnd_net_\,
            in3 => \N__12978\,
            lcout => \uu2.mem0.N_76_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIDKOL_1_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13070\,
            in2 => \_gnd_net_\,
            in3 => \N__12895\,
            lcout => \uu2.N_48_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_i_m4_4_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15512\,
            in1 => \N__17474\,
            in2 => \_gnd_net_\,
            in3 => \N__14943\,
            lcout => \Lab_UT.bcd2segment4.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_26_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__8965\,
            in1 => \N__9907\,
            in2 => \_gnd_net_\,
            in3 => \N__8896\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_2166_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_17_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__10981\,
            in1 => \N__8971\,
            in2 => \N__8914\,
            in3 => \N__9619\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__12338\,
            in1 => \N__10834\,
            in2 => \N__8911\,
            in3 => \N__14794\,
            lcout => \uu2.mem0.w_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_42_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001010000000"
        )
    port map (
            in0 => \N__9711\,
            in1 => \N__10176\,
            in2 => \N__9670\,
            in3 => \N__9780\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_27_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9772\,
            in1 => \N__11125\,
            in2 => \_gnd_net_\,
            in3 => \N__9595\,
            lcout => \uu2.mem0.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_25_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__13316\,
            in1 => \N__13502\,
            in2 => \N__9742\,
            in3 => \N__9640\,
            lcout => \uu2.mem0.g1_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_43_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011111111"
        )
    port map (
            in0 => \N__10177\,
            in1 => \N__9666\,
            in2 => \N__9784\,
            in3 => \N__9712\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_6_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011000011"
        )
    port map (
            in0 => \N__16500\,
            in1 => \N__16417\,
            in2 => \N__16647\,
            in3 => \N__16574\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_186_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8956\,
            in3 => \N__14241\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__17776\
        );

    \uu2.bitmap_RNIMQ601_58_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10765\,
            in2 => \N__9880\,
            in3 => \N__8947\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNIMQ601Z0Z_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_nesr_RNIV0V92_7_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11206\,
            in2 => \N__8953\,
            in3 => \N__9001\,
            lcout => \uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_0_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011101101101"
        )
    port map (
            in0 => \N__16501\,
            in1 => \N__16418\,
            in2 => \N__16648\,
            in3 => \N__16575\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_58_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8950\,
            in3 => \N__14242\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_186C_net\,
            ce => 'H',
            sr => \N__17776\
        );

    \uu2.bitmap_RNI8LB51_186_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10764\,
            in2 => \N__9879\,
            in3 => \N__9007\,
            lcout => \uu2.bitmap_RNI8LB51Z0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_0_2_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__16573\,
            in1 => \N__16636\,
            in2 => \N__16420\,
            in3 => \N__16499\,
            lcout => \Lab_UT.bcd2segment1.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segmentUQ_3_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010010010"
        )
    port map (
            in0 => \N__16643\,
            in1 => \N__16566\,
            in2 => \N__16502\,
            in3 => \N__16408\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_314_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8995\,
            in3 => \N__14230\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__17778\
        );

    \Lab_UT.bcd2segment1.segmentUQ_4_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__16567\,
            in2 => \N__16503\,
            in3 => \N__16409\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_218_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8992\,
            in3 => \N__14229\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__17778\
        );

    \Lab_UT.bcd2segment1.segmentUQ_5_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011010100"
        )
    port map (
            in0 => \N__16645\,
            in1 => \N__16568\,
            in2 => \N__16504\,
            in3 => \N__16410\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_90_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8989\,
            in3 => \N__14231\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__17778\
        );

    \uu2.bitmap_RNIARM01_90_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__8986\,
            in1 => \N__12894\,
            in2 => \N__8980\,
            in3 => \N__10822\,
            lcout => \uu2.bitmap_pmux_19_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_308_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14238\,
            in1 => \N__11314\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__17779\
        );

    \uu2.bitmap_52_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14237\,
            in2 => \_gnd_net_\,
            in3 => \N__11140\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__17779\
        );

    \uu2.bitmap_111_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9199\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__17779\
        );

    \uu2.vram_rd_clk_det_0_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9168\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__17779\
        );

    \uu2.vram_rd_clk_det_1_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9132\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_308C_net\,
            ce => 'H',
            sr => \N__17779\
        );

    \uu0.l_precount_0_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9085\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18030\,
            ce => 'H',
            sr => \N__17827\
        );

    \buart.Z_rx.hh_1_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => \buart.Z_rx.hhZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18090\,
            ce => 'H',
            sr => \N__17831\
        );

    \buart.Z_rx.hh_0_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9055\,
            lcout => \buart.Z_rx.hhZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18083\,
            ce => 'H',
            sr => \N__17829\
        );

    \uu2.r_addr_esr_8_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9382\,
            in1 => \N__9221\,
            in2 => \N__9016\,
            in3 => \N__9027\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18073\,
            ce => \N__9466\,
            sr => \N__17808\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9519\,
            in2 => \_gnd_net_\,
            in3 => \N__9487\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_7_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__9405\,
            in1 => \N__9434\,
            in2 => \N__9535\,
            in3 => \N__9222\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18073\,
            ce => \N__9466\,
            sr => \N__17808\
        );

    \uu2.r_addr_esr_6_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9520\,
            in1 => \N__9489\,
            in2 => \N__9226\,
            in3 => \N__9435\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18073\,
            ce => \N__9466\,
            sr => \N__17808\
        );

    \uu2.r_addr_esr_3_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__9376\,
            in1 => \N__9340\,
            in2 => \N__9294\,
            in3 => \N__9268\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18073\,
            ce => \N__9466\,
            sr => \N__17808\
        );

    \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un426_ci_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13830\,
            in1 => \N__13231\,
            in2 => \N__13753\,
            in3 => \N__13629\,
            lcout => \uu2.un426_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12337\,
            in1 => \N__10077\,
            in2 => \_gnd_net_\,
            in3 => \N__13318\,
            lcout => \uu2.mem0.N_70_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9404\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9370\,
            in1 => \N__9335\,
            in2 => \N__9293\,
            in3 => \N__9263\,
            lcout => \uu2.un404_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_i_1_5_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110101100"
        )
    port map (
            in0 => \N__17492\,
            in1 => \N__14944\,
            in2 => \N__15490\,
            in3 => \N__17252\,
            lcout => \Lab_UT.bcd2segment4.segment_i_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_0_2_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__17488\,
            in1 => \N__14937\,
            in2 => \N__15511\,
            in3 => \N__17248\,
            lcout => \Lab_UT.bcd2segment4.segment_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIG4PV_66_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__9541\,
            in1 => \N__12881\,
            in2 => \N__9556\,
            in3 => \N__10821\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_20_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIKJFQ1_69_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__12882\,
            in1 => \N__9577\,
            in2 => \N__9589\,
            in3 => \N__9568\,
            lcout => \uu2.N_40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_197_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14227\,
            in1 => \_gnd_net_\,
            in2 => \N__9586\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__17781\
        );

    \Lab_UT.bcd2segment4.segment_0_1_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__14941\,
            in1 => \N__17249\,
            in2 => \N__17494\,
            in3 => \N__14226\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_69_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000010110000"
        )
    port map (
            in0 => \N__17251\,
            in1 => \N__15494\,
            in2 => \N__9571\,
            in3 => \N__14344\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__17781\
        );

    \uu2.bitmap_194_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14239\,
            in1 => \N__17250\,
            in2 => \_gnd_net_\,
            in3 => \N__9562\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__17781\
        );

    \uu2.bitmap_66_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14228\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9547\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__17781\
        );

    \uu2.mem0.ram512X8_inst_RNO_38_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__13710\,
            in1 => \N__12974\,
            in2 => \_gnd_net_\,
            in3 => \N__13028\,
            lcout => \uu2.mem0.N_1201_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_53_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__12840\,
            in1 => \N__12696\,
            in2 => \_gnd_net_\,
            in3 => \N__11114\,
            lcout => \uu2.mem0.g0_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep2_RNI1HJ81_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__13709\,
            in1 => \N__12973\,
            in2 => \N__12719\,
            in3 => \N__13030\,
            lcout => \uu2.g2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_37_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011100000"
        )
    port map (
            in0 => \N__13027\,
            in1 => \N__13711\,
            in2 => \N__12979\,
            in3 => \N__12700\,
            lcout => \uu2.mem0.bitmap_pmux_sn_N_20_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_59_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12839\,
            in2 => \_gnd_net_\,
            in3 => \N__11065\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_41_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010010010010"
        )
    port map (
            in0 => \N__13029\,
            in1 => \N__13712\,
            in2 => \N__9643\,
            in3 => \N__12954\,
            lcout => \uu2.mem0.g1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI5R5D8_69_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__9694\,
            in1 => \N__9634\,
            in2 => \N__9628\,
            in3 => \N__10099\,
            lcout => \uu2.N_404\,
            ltout => \uu2.N_404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_16_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__9718\,
            in1 => \N__9613\,
            in2 => \N__9607\,
            in3 => \N__9682\,
            lcout => \uu2.mem0.bitmap_pmux_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_61_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__13213\,
            in1 => \N__10804\,
            in2 => \N__13395\,
            in3 => \N__10762\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_46_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__12738\,
            in1 => \N__12866\,
            in2 => \N__9598\,
            in3 => \N__11113\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_58_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001000"
        )
    port map (
            in0 => \N__13214\,
            in1 => \N__10805\,
            in2 => \N__13396\,
            in3 => \N__10763\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__12739\,
            in1 => \N__12955\,
            in2 => \N__9745\,
            in3 => \N__12865\,
            lcout => OPEN,
            ltout => \uu2.mem0.g1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__9741\,
            in1 => \N__13141\,
            in2 => \N__9727\,
            in3 => \N__9724\,
            lcout => \uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNIT4P31_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110010001000"
        )
    port map (
            in0 => \N__13737\,
            in1 => \N__11112\,
            in2 => \N__12742\,
            in3 => \N__11264\,
            lcout => \uu2.bitmap_pmux_sn_N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIVOBS1_93_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__12867\,
            in1 => \N__10111\,
            in2 => \N__13129\,
            in3 => \N__9703\,
            lcout => \uu2.N_55_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_23_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9688\,
            in1 => \N__9903\,
            in2 => \_gnd_net_\,
            in3 => \N__9649\,
            lcout => \uu2.mem0.N_2166_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNIKIVT_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000110"
        )
    port map (
            in0 => \N__11256\,
            in1 => \N__11110\,
            in2 => \N__10814\,
            in3 => \N__11058\,
            lcout => \uu2.bitmap_pmux_sn_N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_62_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__9811\,
            in2 => \_gnd_net_\,
            in3 => \N__9798\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_247_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_56_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__10799\,
            in1 => \N__11057\,
            in2 => \N__9676\,
            in3 => \N__9855\,
            lcout => OPEN,
            ltout => \uu2.mem0.N_2171_1_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_36_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__12741\,
            in1 => \N__9817\,
            in2 => \N__9673\,
            in3 => \N__9660\,
            lcout => \uu2.mem0.N_397_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__11257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10760\,
            lcout => \uu2.mem0.g1_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI232M_52_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10142\,
            in1 => \N__9810\,
            in2 => \_gnd_net_\,
            in3 => \N__9799\,
            lcout => OPEN,
            ltout => \uu2.N_247_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_7_rep1_nesr_RNI023T1_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__10803\,
            in1 => \N__11059\,
            in2 => \N__9787\,
            in3 => \N__9856\,
            lcout => \uu2.N_2171_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_44_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001000100"
        )
    port map (
            in0 => \N__11111\,
            in1 => \N__13738\,
            in2 => \_gnd_net_\,
            in3 => \N__11258\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.N_198_i_1_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000111"
        )
    port map (
            in0 => \N__17486\,
            in1 => \N__14935\,
            in2 => \N__15526\,
            in3 => \N__17253\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_290_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9766\,
            in3 => \N__14235\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__17780\
        );

    \Lab_UT.bcd2segment4.segment_i_0_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100100010000"
        )
    port map (
            in0 => \N__17487\,
            in1 => \N__14936\,
            in2 => \N__15527\,
            in3 => \N__17254\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_34_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9763\,
            in3 => \N__14236\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__17780\
        );

    \uu2.bitmap_RNI8LAO_34_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100011101"
        )
    port map (
            in0 => \N__9760\,
            in1 => \N__10141\,
            in2 => \N__9754\,
            in3 => \N__10239\,
            lcout => \uu2.bitmap_pmux_15_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_3_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__10241\,
            in1 => \_gnd_net_\,
            in2 => \N__12223\,
            in3 => \N__13804\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__17780\
        );

    \uu2.bitmap_RNILMVP_180_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10240\,
            in2 => \N__9878\,
            in3 => \N__9847\,
            lcout => \uu2.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_180_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14234\,
            in2 => \_gnd_net_\,
            in3 => \N__11149\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_290C_net\,
            ce => 'H',
            sr => \N__17780\
        );

    \Lab_UT.bcd2segment3.segmentUQ_3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100110"
        )
    port map (
            in0 => \N__15730\,
            in1 => \N__15981\,
            in2 => \N__16080\,
            in3 => \N__15819\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9841\,
            in3 => \N__14232\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__17784\
        );

    \Lab_UT.bcd2segment3.segment_0_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111101111001"
        )
    port map (
            in0 => \N__15731\,
            in1 => \N__15982\,
            in2 => \N__16081\,
            in3 => \N__15820\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_40_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9838\,
            in3 => \N__14233\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__17784\
        );

    \uu2.bitmap_RNI2S3H1_40_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101111"
        )
    port map (
            in0 => \N__9835\,
            in1 => \N__9829\,
            in2 => \N__11074\,
            in3 => \N__9823\,
            lcout => \uu2.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__10048\,
            in1 => \N__10243\,
            in2 => \_gnd_net_\,
            in3 => \N__10198\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_sn_N_54_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNITQGB1_111_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9934\,
            in2 => \N__9928\,
            in3 => \N__10213\,
            lcout => OPEN,
            ltout => \uu2.N_395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNIJ9KQ3_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9925\,
            in2 => \N__9916\,
            in3 => \N__9913\,
            lcout => \uu2.N_401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18025\,
            ce => \N__11713\,
            sr => \N__17828\
        );

    \buart.Z_rx.shifter_6_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11347\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18025\,
            ce => \N__11713\,
            sr => \N__17828\
        );

    \buart.Z_rx.shifter_7_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9979\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18025\,
            ce => \N__11713\,
            sr => \N__17828\
        );

    \buart.Z_rx.bitcount_RNI9OJJ_1_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10577\,
            in2 => \_gnd_net_\,
            in3 => \N__10356\,
            lcout => OPEN,
            ltout => \buart.Z_rx.idle_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_4_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10482\,
            in1 => \N__10543\,
            in2 => \N__9886\,
            in3 => \N__11739\,
            lcout => \buart.Z_rx.idle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIAPJJ_1_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10481\,
            in2 => \_gnd_net_\,
            in3 => \N__10355\,
            lcout => OPEN,
            ltout => \buart.Z_rx.valid_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNI9F1H1_0_4_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__10542\,
            in2 => \N__9883\,
            in3 => \N__11738\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_RNI065O1_0_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9972\,
            in1 => \N__9961\,
            in2 => \_gnd_net_\,
            in3 => \N__11825\,
            lcout => \buart.Z_rx.startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11746\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10357\,
            in2 => \_gnd_net_\,
            in3 => \N__9946\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10579\,
            in2 => \_gnd_net_\,
            in3 => \N__9943\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10484\,
            in2 => \_gnd_net_\,
            in3 => \N__9940\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010100111010"
        )
    port map (
            in0 => \N__10545\,
            in1 => \N__11996\,
            in2 => \N__10510\,
            in3 => \N__9937\,
            lcout => \buart.Z_rx.bitcount_lm_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI8NF3_8_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10076\,
            in2 => \_gnd_net_\,
            in3 => \N__10008\,
            lcout => \uu2.N_153\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__12648\,
            in1 => \N__12544\,
            in2 => \N__10440\,
            in3 => \N__11911\,
            lcout => \uu2.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNO_0_6_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__11912\,
            in1 => \N__10435\,
            in2 => \N__12552\,
            in3 => \N__12649\,
            lcout => OPEN,
            ltout => \uu2.N_150_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_6_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10022\,
            in1 => \N__12509\,
            in2 => \N__10084\,
            in3 => \N__12597\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_6C_net\,
            ce => \N__10621\,
            sr => \N__17790\
        );

    \uu2.w_addr_user_nesr_8_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101010000"
        )
    port map (
            in0 => \N__12598\,
            in1 => \N__10023\,
            in2 => \N__10081\,
            in3 => \N__10007\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_6C_net\,
            ce => \N__10621\,
            sr => \N__17790\
        );

    \uu2.w_addr_user_nesr_0_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__10715\,
            in1 => \N__12548\,
            in2 => \N__12514\,
            in3 => \N__12596\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_6C_net\,
            ce => \N__10621\,
            sr => \N__17790\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10714\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__12883\,
            lcout => \uu2.mem0.N_78_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__12196\,
            in1 => \N__13594\,
            in2 => \N__13840\,
            in3 => \N__13716\,
            lcout => \uu2.w_addr_displayingZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_displaying_3_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__13593\,
            in1 => \N__13831\,
            in2 => \_gnd_net_\,
            in3 => \N__12194\,
            lcout => \uu2.w_addr_displayingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_displaying_3_rep2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__12195\,
            in1 => \_gnd_net_\,
            in2 => \N__13839\,
            in3 => \N__12733\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_displaying_fast_2_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13069\,
            in1 => \N__12884\,
            in2 => \N__10047\,
            in3 => \N__12197\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_user_1_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010011110000"
        )
    port map (
            in0 => \N__12586\,
            in1 => \N__10723\,
            in2 => \N__10685\,
            in3 => \N__12485\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_user_7_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100000010"
        )
    port map (
            in0 => \N__12487\,
            in1 => \N__12588\,
            in2 => \N__10027\,
            in3 => \N__10006\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.w_addr_user_4_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000111110000"
        )
    port map (
            in0 => \N__12587\,
            in1 => \N__10439\,
            in2 => \N__12659\,
            in3 => \N__12486\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.bitmap_221_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10123\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14240\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__17786\
        );

    \uu2.mem0.ram512X8_inst_RNO_48_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13682\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11115\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_55_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12716\,
            in1 => \N__12945\,
            in2 => \N__13506\,
            in3 => \N__13384\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_35_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13683\,
            in1 => \N__10923\,
            in2 => \N__10102\,
            in3 => \N__13230\,
            lcout => \uu2.mem0.un49_w_data_displaying_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_rep1_RNI5QH04_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110001010000"
        )
    port map (
            in0 => \N__12718\,
            in1 => \N__11066\,
            in2 => \N__11218\,
            in3 => \N__10279\,
            lcout => \uu2.bitmap_pmux_27_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_54_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13681\,
            in1 => \N__13494\,
            in2 => \N__13402\,
            in3 => \N__13229\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_6_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_34_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10093\,
            in1 => \N__13306\,
            in2 => \N__10087\,
            in3 => \N__13052\,
            lcout => \uu2.mem0.un31_w_data_displaying_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNIFG6E_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13680\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11262\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_47_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12717\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12868\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12220\,
            in1 => \N__12879\,
            in2 => \N__13072\,
            in3 => \N__11116\,
            lcout => \uu2.w_addr_displaying_2_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12876\,
            in1 => \_gnd_net_\,
            in2 => \N__12221\,
            in3 => \N__13064\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_6_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011111111001000"
        )
    port map (
            in0 => \N__12250\,
            in1 => \N__12215\,
            in2 => \N__10159\,
            in3 => \N__13394\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12878\,
            in1 => \N__13065\,
            in2 => \N__12972\,
            in3 => \N__12219\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_0_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12206\,
            in2 => \_gnd_net_\,
            in3 => \N__12875\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_fast_1_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__12880\,
            in1 => \_gnd_net_\,
            in2 => \N__12222\,
            in3 => \N__10197\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_1_rep1_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__11265\,
            in1 => \N__12877\,
            in2 => \_gnd_net_\,
            in3 => \N__12210\,
            lcout => \uu2.w_addr_displaying_1_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_3_rep1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__12211\,
            in1 => \N__13824\,
            in2 => \_gnd_net_\,
            in3 => \N__11067\,
            lcout => \uu2.w_addr_displaying_3_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_2_rep1C_net\,
            ce => 'H',
            sr => \N__17777\
        );

    \uu2.w_addr_displaying_fast_nesr_8_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000100"
        )
    port map (
            in0 => \N__13802\,
            in1 => \N__13624\,
            in2 => \N__10885\,
            in3 => \N__10144\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            ce => \N__13533\,
            sr => \N__17782\
        );

    \uu2.w_addr_displaying_RNI50L01_2_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__12969\,
            in1 => \N__13050\,
            in2 => \_gnd_net_\,
            in3 => \N__12864\,
            lcout => \uu2.N_46\,
            ltout => \uu2.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_nesr_7_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100110"
        )
    port map (
            in0 => \N__11205\,
            in1 => \N__13623\,
            in2 => \N__10201\,
            in3 => \N__13109\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            ce => \N__13533\,
            sr => \N__17782\
        );

    \uu2.w_addr_displaying_8_rep1_nesr_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__10759\,
            in1 => \N__10880\,
            in2 => \N__13630\,
            in3 => \N__13801\,
            lcout => \uu2.w_addr_displaying_8_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            ce => \N__13533\,
            sr => \N__17782\
        );

    \uu2.w_addr_displaying_nesr_7_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110100"
        )
    port map (
            in0 => \N__13803\,
            in1 => \N__13625\,
            in2 => \N__13498\,
            in3 => \N__13110\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            ce => \N__13533\,
            sr => \N__17782\
        );

    \uu2.w_addr_displaying_7_rep1_nesr_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000010"
        )
    port map (
            in0 => \N__13619\,
            in1 => \N__13800\,
            in2 => \N__13111\,
            in3 => \N__10813\,
            lcout => \uu2.w_addr_displaying_7_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_fast_nesr_8C_net\,
            ce => \N__13533\,
            sr => \N__17782\
        );

    \uu2.w_addr_displaying_fast_RNIETIP_1_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__11064\,
            in1 => \N__10196\,
            in2 => \_gnd_net_\,
            in3 => \N__10758\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segmentUQ_4_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__15821\,
            in2 => \N__15738\,
            in3 => \N__16078\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_200_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10162\,
            in3 => \N__14223\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_200C_net\,
            ce => 'H',
            sr => \N__17785\
        );

    \Lab_UT.bcd2segment3.segmentUQ_5_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011010100"
        )
    port map (
            in0 => \N__15984\,
            in1 => \N__15822\,
            in2 => \N__15739\,
            in3 => \N__16079\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_72_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10285\,
            in3 => \N__14225\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_200C_net\,
            ce => 'H',
            sr => \N__17785\
        );

    \uu2.bitmap_RNI011L_75_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10315\,
            in1 => \N__11201\,
            in2 => \_gnd_net_\,
            in3 => \N__10252\,
            lcout => OPEN,
            ltout => \uu2.N_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNI588O1_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000011001"
        )
    port map (
            in0 => \N__12888\,
            in1 => \N__11266\,
            in2 => \N__10282\,
            in3 => \N__10258\,
            lcout => \uu2.g0_17_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIQQ0L_72_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10270\,
            in1 => \N__10264\,
            in2 => \_gnd_net_\,
            in3 => \N__11200\,
            lcout => \uu2.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_203_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10303\,
            in2 => \_gnd_net_\,
            in3 => \N__14224\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_200C_net\,
            ce => 'H',
            sr => \N__17785\
        );

    \Lab_UT.bcd2segment3.segmentUQ_6_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100111100001"
        )
    port map (
            in0 => \N__15980\,
            in1 => \N__15818\,
            in2 => \N__16071\,
            in3 => \N__15729\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_168_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__14217\,
            in1 => \_gnd_net_\,
            in2 => \N__10246\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__17789\
        );

    \uu2.bitmap_RNISSSN_162_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10207\,
            in1 => \N__10242\,
            in2 => \_gnd_net_\,
            in3 => \N__10219\,
            lcout => \uu2.bitmap_RNISSSNZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14216\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11287\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__17789\
        );

    \Lab_UT.bcd2segment3.segment_i_1_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011111111"
        )
    port map (
            in0 => \N__15979\,
            in1 => \N__15898\,
            in2 => \N__16070\,
            in3 => \N__14215\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10318\,
            in3 => \N__10309\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_168C_net\,
            ce => 'H',
            sr => \N__17789\
        );

    \Lab_UT.bcd2segment3.segment_i_0_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101000"
        )
    port map (
            in0 => \N__15977\,
            in1 => \N__15814\,
            in2 => \N__16069\,
            in3 => \N__15728\,
            lcout => \Lab_UT.bcd2segment3.segment_i_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.segment_i_0_2_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000010000"
        )
    port map (
            in0 => \N__15727\,
            in1 => \N__16049\,
            in2 => \N__15823\,
            in3 => \N__15978\,
            lcout => \Lab_UT.bcd2segment3.segment_i_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_1_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11461\,
            in1 => \N__11493\,
            in2 => \N__11398\,
            in3 => \N__13980\,
            lcout => \Lab_UT.dictrl.next_alarmstate4_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_3_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__13981\,
            in1 => \N__11394\,
            in2 => \N__11500\,
            in3 => \N__11462\,
            lcout => \resetGen.escKeyZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state16_4_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11460\,
            in1 => \N__11492\,
            in2 => \N__11397\,
            in3 => \N__13979\,
            lcout => \Lab_UT.dictrl.next_state16Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11497\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18021\,
            ce => \N__11712\,
            sr => \N__17830\
        );

    \Lab_UT.dictrl.next_state_1_sqmuxa_2_0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11459\,
            in1 => \N__11491\,
            in2 => \N__11531\,
            in3 => \N__13978\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxa_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_2_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11395\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18021\,
            ce => \N__11712\,
            sr => \N__17830\
        );

    \buart.Z_rx.shifter_4_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11524\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18021\,
            ce => \N__11712\,
            sr => \N__17830\
        );

    \buart.Z_rx.shifter_3_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11463\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18021\,
            ce => \N__11712\,
            sr => \N__17830\
        );

    \buart.Z_rx.bitcount_RNIMK771_4_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10580\,
            in1 => \N__10483\,
            in2 => \N__10360\,
            in3 => \N__10544\,
            lcout => \buart.Z_rx.un1_sample_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIIU223_4_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11826\,
            in2 => \_gnd_net_\,
            in3 => \N__11795\,
            lcout => \buart.Z_rx.N_27_0_i\,
            ltout => \buart.Z_rx.N_27_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNO_0_0_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__11997\,
            in1 => \N__10412\,
            in2 => \N__10378\,
            in3 => \N__11743\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_0_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__11744\,
            in1 => \N__11772\,
            in2 => \N__10375\,
            in3 => \N__11998\,
            lcout => \buart.Z_rx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18091\,
            ce => 'H',
            sr => \N__17834\
        );

    \buart.Z_rx.bitcount_RNO_0_1_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__11999\,
            in1 => \N__10358\,
            in2 => \N__10372\,
            in3 => \N__10507\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_1_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__10359\,
            in1 => \N__11773\,
            in2 => \N__10363\,
            in3 => \N__12002\,
            lcout => \buart.Z_rx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18084\,
            ce => 'H',
            sr => \N__17833\
        );

    \buart.Z_rx.bitcount_RNO_0_2_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__12000\,
            in1 => \N__10581\,
            in2 => \N__10327\,
            in3 => \N__10508\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_2_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__10582\,
            in1 => \N__11774\,
            in2 => \N__10585\,
            in3 => \N__12003\,
            lcout => \buart.Z_rx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18084\,
            ce => 'H',
            sr => \N__17833\
        );

    \buart.Z_rx.bitcount_4_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__12005\,
            in1 => \N__10546\,
            in2 => \N__11779\,
            in3 => \N__10552\,
            lcout => \buart.Z_rx.bitcountZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18084\,
            ce => 'H',
            sr => \N__17833\
        );

    \buart.Z_rx.bitcount_RNO_0_3_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111100"
        )
    port map (
            in0 => \N__12001\,
            in1 => \N__10485\,
            in2 => \N__10519\,
            in3 => \N__10509\,
            lcout => OPEN,
            ltout => \buart.Z_rx.bitcount_lm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_3_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__10486\,
            in1 => \N__11775\,
            in2 => \N__10489\,
            in3 => \N__12004\,
            lcout => \buart.Z_rx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18084\,
            ce => 'H',
            sr => \N__17833\
        );

    \uu2.w_addr_user_RNIPJCC_1_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10716\,
            in1 => \N__11854\,
            in2 => \N__10687\,
            in3 => \N__10456\,
            lcout => \uu2.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIFBD5_3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__10717\,
            in1 => \N__11936\,
            in2 => \N__10682\,
            in3 => \N__11878\,
            lcout => \uu2.N_90\,
            ltout => \uu2.N_90_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_3_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__12581\,
            in1 => \_gnd_net_\,
            in2 => \N__10450\,
            in3 => \N__10447\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__10617\,
            sr => \N__17792\
        );

    \uu2.w_addr_user_nesr_RNO_0_3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__10718\,
            in1 => \N__11937\,
            in2 => \N__10683\,
            in3 => \N__11879\,
            lcout => \uu2.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_5_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101000100"
        )
    port map (
            in0 => \N__12582\,
            in1 => \N__11913\,
            in2 => \N__10441\,
            in3 => \N__12653\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__10617\,
            sr => \N__17792\
        );

    \uu2.w_addr_user_nesr_2_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__10719\,
            in1 => \N__11880\,
            in2 => \N__10684\,
            in3 => \N__12580\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_3C_net\,
            ce => \N__10617\,
            sr => \N__17792\
        );

    \Lab_UT.dictrl.state_ret_4_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101110101011"
        )
    port map (
            in0 => \N__17644\,
            in1 => \N__11635\,
            in2 => \N__11650\,
            in3 => \N__11602\,
            lcout => \Lab_UT.dictrl.state_retZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111010101"
        )
    port map (
            in0 => \N__15171\,
            in1 => \N__15243\,
            in2 => \N__16255\,
            in3 => \N__15381\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_18_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__14987\,
            in1 => \N__12459\,
            in2 => \_gnd_net_\,
            in3 => \N__12366\,
            lcout => \uu2.mem0.N_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI34K17_8_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17642\,
            in2 => \_gnd_net_\,
            in3 => \N__12163\,
            lcout => \uu2.un21_w_addr_displaying_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNIB4K34_6_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12477\,
            lcout => \uu2.un28_w_addr_user_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11910\,
            in1 => \N__12282\,
            in2 => \_gnd_net_\,
            in3 => \N__13225\,
            lcout => \uu2.mem0.N_73_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15316\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18062\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_32_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13376\,
            in1 => \N__12946\,
            in2 => \N__13504\,
            in3 => \N__13707\,
            lcout => \uu2.mem0.g0_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI25P31_0_8_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13032\,
            in1 => \N__13280\,
            in2 => \_gnd_net_\,
            in3 => \N__12859\,
            lcout => \uu2.un49_w_data_displaying_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNI25P31_8_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__12860\,
            in1 => \_gnd_net_\,
            in2 => \N__13304\,
            in3 => \N__13031\,
            lcout => OPEN,
            ltout => \uu2.un31_w_data_displaying_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIFOBB3_2_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12947\,
            in1 => \N__13577\,
            in2 => \N__10960\,
            in3 => \N__10933\,
            lcout => \uu2.un31_w_data_displaying\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNISQPH1_7_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13374\,
            in1 => \N__13200\,
            in2 => \N__13503\,
            in3 => \N__13706\,
            lcout => \uu2.un15_w_data_displaying_6\,
            ltout => \uu2.un15_w_data_displaying_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIFOBB3_0_2_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12948\,
            in1 => \N__13578\,
            in2 => \N__10927\,
            in3 => \N__10924\,
            lcout => \uu2.un49_w_data_displaying\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNISQPH1_0_7_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__13375\,
            in1 => \N__13201\,
            in2 => \N__13505\,
            in3 => \N__13708\,
            lcout => \uu2.un15_w_data_displaying_i_i_o2_0\,
            ltout => \uu2.un15_w_data_displaying_i_i_o2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_8_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100110"
        )
    port map (
            in0 => \N__13303\,
            in1 => \N__13579\,
            in2 => \N__10861\,
            in3 => \N__13828\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_8C_net\,
            ce => \N__13523\,
            sr => \N__17787\
        );

    \uu2.mem0.ram512X8_inst_RNO_20_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__10858\,
            in1 => \N__10969\,
            in2 => \N__10852\,
            in3 => \N__10840\,
            lcout => \uu2.mem0.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_60_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__13373\,
            in1 => \N__10806\,
            in2 => \_gnd_net_\,
            in3 => \N__10761\,
            lcout => OPEN,
            ltout => \uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_45_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__13216\,
            in1 => \N__11006\,
            in2 => \N__11128\,
            in3 => \N__11017\,
            lcout => \uu2.mem0.ram512X8_inst_RNOZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_rep1_RNIDKIL_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11109\,
            in2 => \_gnd_net_\,
            in3 => \N__11063\,
            lcout => \uu2.bitmap_pmux_sn_N_31_0\,
            ltout => \uu2.bitmap_pmux_sn_N_31_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_49_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100000"
        )
    port map (
            in0 => \N__13464\,
            in1 => \N__13290\,
            in2 => \N__11011\,
            in3 => \N__11007\,
            lcout => OPEN,
            ltout => \uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_28_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000100000"
        )
    port map (
            in0 => \N__11008\,
            in1 => \N__10996\,
            in2 => \N__10990\,
            in3 => \N__10987\,
            lcout => \uu2.mem0.bitmap_pmux_u_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_52_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12734\,
            in2 => \_gnd_net_\,
            in3 => \N__13215\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_33_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13289\,
            in1 => \N__13051\,
            in2 => \N__10972\,
            in3 => \N__12874\,
            lcout => \uu2.mem0.g0_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_i_0_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010000000"
        )
    port map (
            in0 => \N__17548\,
            in1 => \N__16243\,
            in2 => \N__16319\,
            in3 => \N__16155\,
            lcout => \Lab_UT.bcd2segment2.segment_i_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_i_0_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000100"
        )
    port map (
            in0 => \N__16156\,
            in1 => \N__16308\,
            in2 => \N__16251\,
            in3 => \N__17549\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10963\,
            in3 => \N__14209\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__17788\
        );

    \uu2.bitmap_RNI693L_87_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13864\,
            in1 => \N__11199\,
            in2 => \_gnd_net_\,
            in3 => \N__11272\,
            lcout => OPEN,
            ltout => \uu2.N_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_rep1_RNIHOCO1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111001111111"
        )
    port map (
            in0 => \N__12852\,
            in1 => \N__11263\,
            in2 => \N__11221\,
            in3 => \N__11173\,
            lcout => \uu2.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI033L_84_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11161\,
            in1 => \N__11167\,
            in2 => \_gnd_net_\,
            in3 => \N__11198\,
            lcout => \uu2.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_84_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14210\,
            in2 => \_gnd_net_\,
            in3 => \N__11155\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__17788\
        );

    \uu2.bitmap_212_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__14211\,
            in1 => \N__11302\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__17788\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_1_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101001101"
        )
    port map (
            in0 => \N__16223\,
            in1 => \N__16145\,
            in2 => \N__16311\,
            in3 => \N__17546\,
            lcout => \Lab_UT.didp.countrce2.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_0_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011001010110"
        )
    port map (
            in0 => \N__17544\,
            in1 => \N__16291\,
            in2 => \N__16163\,
            in3 => \N__16222\,
            lcout => \Lab_UT.didp.countrce2.N_175\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010100000000110"
        )
    port map (
            in0 => \N__16221\,
            in1 => \N__16138\,
            in2 => \N__16310\,
            in3 => \N__17543\,
            lcout => \Lab_UT.didp.countrce2.N_170\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.un1_num_7_1_0_a2_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17452\,
            lcout => \Lab_UT.N_68_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_2_1_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101111001"
        )
    port map (
            in0 => \N__16220\,
            in1 => \N__16137\,
            in2 => \N__16309\,
            in3 => \N__17542\,
            lcout => \Lab_UT.didp.countrce2.N_183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_1_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000111"
        )
    port map (
            in0 => \N__17545\,
            in1 => \N__16292\,
            in2 => \N__16164\,
            in3 => \N__16224\,
            lcout => \Lab_UT.didp.countrce2.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001010"
        )
    port map (
            in0 => \N__17453\,
            in1 => \N__11293\,
            in2 => \N__17341\,
            in3 => \N__17285\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__16348\,
            in1 => \N__16296\,
            in2 => \N__15859\,
            in3 => \N__16225\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101010101"
        )
    port map (
            in0 => \N__17473\,
            in1 => \N__14916\,
            in2 => \N__15529\,
            in3 => \N__17221\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.N_80_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__17363\,
            in1 => \_gnd_net_\,
            in2 => \N__11296\,
            in3 => \N__11396\,
            lcout => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.segment_i_0_6_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100110101001"
        )
    port map (
            in0 => \N__17472\,
            in1 => \N__14915\,
            in2 => \N__15528\,
            in3 => \N__17220\,
            lcout => \Lab_UT.bcd2segment4.segment_i_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11361\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate4_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11431\,
            in1 => \N__11281\,
            in2 => \N__11275\,
            in3 => \N__17386\,
            lcout => \Lab_UT.next_alarmstate4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__17362\,
            in1 => \N__14350\,
            in2 => \_gnd_net_\,
            in3 => \N__11499\,
            lcout => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state16_5_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11430\,
            in1 => \N__11532\,
            in2 => \N__11362\,
            in3 => \N__17385\,
            lcout => \resetGen_escKey_4\,
            ltout => \resetGen_escKey_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14604\,
            in2 => \N__11536\,
            in3 => \N__14034\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_sqmuxa_2_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11530\,
            in1 => \N__11498\,
            in2 => \N__11429\,
            in3 => \N__13982\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11387\,
            in1 => \N__11437\,
            in2 => \N__11467\,
            in3 => \N__11464\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNI0C5J6_2_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__14125\,
            in1 => \N__11590\,
            in2 => \N__11440\,
            in3 => \N__13884\,
            lcout => \Lab_UT.dictrl.next_state_set\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.escKey_2_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__17388\,
            in1 => \N__11351\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \resetGen_escKey_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_sqmuxa_3_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__11419\,
            in1 => \N__11386\,
            in2 => \N__11357\,
            in3 => \N__17387\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_RNICD593_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11323\,
            in2 => \N__11317\,
            in3 => \N__14124\,
            lcout => \Lab_UT.dictrl.next_state_1_sqmuxa\,
            ltout => \Lab_UT.dictrl.next_state_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNI1GK36_2_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__11586\,
            in1 => \_gnd_net_\,
            in2 => \N__11575\,
            in3 => \N__11559\,
            lcout => \Lab_UT.dictrl.next_state_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13983\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18026\,
            ce => \N__11705\,
            sr => \N__17832\
        );

    \Lab_UT.dictrl.next_state_RNIN0UD1_2_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14260\,
            in2 => \_gnd_net_\,
            in3 => \N__11569\,
            lcout => \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m37_ns_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000011"
        )
    port map (
            in0 => \N__17073\,
            in1 => \N__14641\,
            in2 => \N__14603\,
            in3 => \N__17008\,
            lcout => \Lab_UT.m37_ns\,
            ltout => \Lab_UT.m37_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_2_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__14492\,
            in1 => \N__14282\,
            in2 => \N__11572\,
            in3 => \N__14308\,
            lcout => \Lab_UT.dictrl.next_state_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18022\,
            ce => \N__14389\,
            sr => \N__11563\
        );

    \Lab_UT.didp.m45_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011000000"
        )
    port map (
            in0 => \N__17072\,
            in1 => \N__17009\,
            in2 => \N__14602\,
            in3 => \N__16786\,
            lcout => \Lab_UT.m45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m40_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001100000"
        )
    port map (
            in0 => \N__16785\,
            in1 => \N__14587\,
            in2 => \N__17018\,
            in3 => \N__17074\,
            lcout => \Lab_UT.m40\,
            ltout => \Lab_UT.m40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI970U_3_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13912\,
            in2 => \N__11542\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3\,
            ltout => \Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNISML65_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__16863\,
            in1 => \N__15622\,
            in2 => \N__11539\,
            in3 => \N__15569\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m34_ns_1_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__17071\,
            in1 => \N__17004\,
            in2 => \_gnd_net_\,
            in3 => \N__16784\,
            lcout => \Lab_UT.didp.m34_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNI919D9_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__16961\,
            in1 => \N__16941\,
            in2 => \N__16911\,
            in3 => \N__16805\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_0\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNI4EJF21_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__11625\,
            in1 => \N__14085\,
            in2 => \N__11638\,
            in3 => \N__14073\,
            lcout => \Lab_UT.dictrl.un1_state_21_reti_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__16962\,
            in1 => \N__16942\,
            in2 => \N__14497\,
            in3 => \N__16806\,
            lcout => \Lab_UT.dictrl.next_state_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18020\,
            ce => \N__14383\,
            sr => \N__13894\
        );

    \Lab_UT.dictrl.state_ret_4_RNI4Q509_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__14261\,
            in1 => \N__14281\,
            in2 => \N__16887\,
            in3 => \N__14311\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11614\,
            in2 => \_gnd_net_\,
            in3 => \N__16940\,
            lcout => \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIO0LS1_1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14395\,
            in2 => \_gnd_net_\,
            in3 => \N__14445\,
            lcout => \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1\,
            ltout => \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNIRRERA_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__14416\,
            in1 => \N__16867\,
            in2 => \N__11608\,
            in3 => \N__14446\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_1\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNINI42G_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11605\,
            in3 => \N__14072\,
            lcout => \Lab_UT.dictrl.dicRun_2_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__12017\,
            in1 => \N__11665\,
            in2 => \N__12081\,
            in3 => \N__12048\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__12018\,
            in1 => \N__12047\,
            in2 => \N__12082\,
            in3 => \N__12142\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12135\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12016\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNILM873_4_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__12073\,
            in1 => \N__12046\,
            in2 => \N__11833\,
            in3 => \N__11805\,
            lcout => \buart.Z_rx.bitcountlde_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNIU4N1_2_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11677\,
            in2 => \_gnd_net_\,
            in3 => \N__12134\,
            lcout => \buart.Z_rx.ser_clk_2\,
            ltout => \buart.Z_rx.ser_clk_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__11755\,
            in2 => \N__11749\,
            in3 => \N__11745\,
            lcout => \buart.Z_rx.sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12092\,
            in2 => \N__12136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11676\,
            in2 => \_gnd_net_\,
            in3 => \N__11659\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12026\,
            in1 => \N__12114\,
            in2 => \_gnd_net_\,
            in3 => \N__11656\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__18092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11959\,
            in2 => \_gnd_net_\,
            in3 => \N__11653\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12105\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12145\,
            lcout => \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__12094\,
            in1 => \N__12133\,
            in2 => \_gnd_net_\,
            in3 => \N__12028\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11958\,
            in1 => \N__12115\,
            in2 => \N__12106\,
            in3 => \N__12093\,
            lcout => \buart.Z_rx.ser_clk_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__12080\,
            in1 => \N__12058\,
            in2 => \N__12052\,
            in3 => \N__12027\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18092\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__17293\,
            in1 => \N__11950\,
            in2 => \N__17336\,
            in3 => \N__15486\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18074\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m24_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__15382\,
            in1 => \N__15174\,
            in2 => \_gnd_net_\,
            in3 => \N__15271\,
            lcout => \Lab_UT.m24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNINJD5_3_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12660\,
            in1 => \N__11932\,
            in2 => \N__11914\,
            in3 => \N__11874\,
            lcout => \uu2.w_addr_user_3_i_a2_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12540\,
            in1 => \N__12281\,
            in2 => \_gnd_net_\,
            in3 => \N__13410\,
            lcout => \uu2.mem0.N_72_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13747\,
            in1 => \N__12280\,
            in2 => \_gnd_net_\,
            in3 => \N__12661\,
            lcout => \uu2.mem0.N_74_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__15029\,
            in1 => \N__15037\,
            in2 => \N__12610\,
            in3 => \N__16481\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18068\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_o2_0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__14721\,
            in1 => \N__14655\,
            in2 => \N__14676\,
            in3 => \N__14777\,
            lcout => \uu2.N_84\,
            ltout => \uu2.N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un28_w_addr_user_i_0_a3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000100"
        )
    port map (
            in0 => \N__14700\,
            in1 => \N__14977\,
            in2 => \N__12601\,
            in3 => \N__12458\,
            lcout => \uu2.N_97\,
            ltout => \uu2.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI7BP14_6_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__12396\,
            in1 => \N__12553\,
            in2 => \N__12517\,
            in3 => \N__12510\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_data_0_o2_0_4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__14699\,
            in1 => \N__14976\,
            in2 => \_gnd_net_\,
            in3 => \N__12457\,
            lcout => \uu2.N_86\,
            ltout => \uu2.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_i_0_tz_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101011111"
        )
    port map (
            in0 => \N__12395\,
            in1 => \_gnd_net_\,
            in2 => \N__12382\,
            in3 => \N__12365\,
            lcout => \uu2.w_addr_i_0_tzZ0Z_0\,
            ltout => \uu2.w_addr_i_0_tzZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_RNIVAPV6_8_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12253\,
            in3 => \N__12246\,
            lcout => \uu2.un21_w_addr_displaying_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIRJ7L_3_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15377\,
            in1 => \N__15170\,
            in2 => \_gnd_net_\,
            in3 => \N__15241\,
            lcout => \Lab_UT.dispString.un22_dOutP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__17638\,
            in1 => \_gnd_net_\,
            in2 => \N__15655\,
            in3 => \N__14323\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18063\,
            ce => 'H',
            sr => \N__17126\
        );

    \Lab_UT.didp.reset_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15651\,
            in2 => \_gnd_net_\,
            in3 => \N__17637\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18063\,
            ce => 'H',
            sr => \N__17126\
        );

    \uu2.w_addr_displaying_RNI8BP31_6_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__13746\,
            in1 => \N__13411\,
            in2 => \_gnd_net_\,
            in3 => \N__13212\,
            lcout => \uu2.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_51_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13501\,
            in1 => \N__13062\,
            in2 => \N__13751\,
            in3 => \N__13287\,
            lcout => OPEN,
            ltout => \uu2.mem0.g0_7_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_31_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__13846\,
            in1 => \N__12971\,
            in2 => \N__13090\,
            in3 => \N__12893\,
            lcout => OPEN,
            ltout => \uu2.mem0.un31_w_data_displaying_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_19_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__12748\,
            in1 => \N__12754\,
            in2 => \N__13087\,
            in3 => \N__13288\,
            lcout => \uu2.mem0.g1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_29_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13063\,
            in1 => \N__12970\,
            in2 => \N__13626\,
            in3 => \N__12892\,
            lcout => \uu2.mem0.g1_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_30_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13204\,
            in1 => \N__13500\,
            in2 => \N__13409\,
            in3 => \N__13739\,
            lcout => \uu2.mem0.g1_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_50_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12740\,
            in1 => \N__13398\,
            in2 => \_gnd_net_\,
            in3 => \N__13203\,
            lcout => \uu2.mem0.g0_7_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_5_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__13205\,
            in1 => \N__13838\,
            in2 => \N__13752\,
            in3 => \N__13609\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_5C_net\,
            ce => \N__13534\,
            sr => \N__17783\
        );

    \uu2.mem0.ram512X8_inst_RNO_39_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__13499\,
            in1 => \N__13397\,
            in2 => \N__13305\,
            in3 => \N__13202\,
            lcout => \uu2.mem0.g0_16_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.segment_1_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110111010111"
        )
    port map (
            in0 => \N__16611\,
            in1 => \N__16460\,
            in2 => \N__16406\,
            in3 => \N__16548\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__14208\,
            in1 => \_gnd_net_\,
            in2 => \N__13132\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__17791\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__16461\,
            in1 => \_gnd_net_\,
            in2 => \N__16569\,
            in3 => \N__16613\,
            lcout => \Lab_UT.didp.countrce1.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.un1_num_11_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16612\,
            in1 => \N__16459\,
            in2 => \N__16407\,
            in3 => \N__16549\,
            lcout => \Lab_UT.nine\,
            ltout => \Lab_UT.nine_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNI84NN1_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17551\,
            in1 => \N__16160\,
            in2 => \N__13114\,
            in3 => \N__16711\,
            lcout => \Lab_UT.didp.q_RNI84NN1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment2.segment_i_1_1_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__16710\,
            in1 => \N__17550\,
            in2 => \N__16172\,
            in3 => \N__14207\,
            lcout => OPEN,
            ltout => \Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13873\,
            in2 => \N__13867\,
            in3 => \_gnd_net_\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__17791\
        );

    \Lab_UT.didp.countrce1.q_1_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001100"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__16554\,
            in2 => \N__16671\,
            in3 => \N__16467\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__16466\,
            in1 => \N__17143\,
            in2 => \_gnd_net_\,
            in3 => \N__16663\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment1.un1_num_5_2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16553\,
            in2 => \_gnd_net_\,
            in3 => \N__16465\,
            lcout => OPEN,
            ltout => \Lab_UT.three_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__16667\,
            in1 => \N__17146\,
            in2 => \N__13855\,
            in3 => \N__16617\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__16341\,
            in1 => \N__16180\,
            in2 => \N__15855\,
            in3 => \N__16162\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__16340\,
            in1 => \N__16087\,
            in2 => \N__17560\,
            in3 => \N__15851\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15847\,
            in1 => \N__16339\,
            in2 => \_gnd_net_\,
            in3 => \N__16239\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__13852\,
            in1 => \N__17144\,
            in2 => \N__16672\,
            in3 => \N__16397\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18045\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_set_0_1_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14006\,
            in2 => \_gnd_net_\,
            in3 => \N__14040\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNILGF17_3_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__14547\,
            in1 => \N__14751\,
            in2 => \N__14059\,
            in3 => \N__14056\,
            lcout => \Lab_UT.dictrl.next_state_set_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m34_ns_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011101010"
        )
    port map (
            in0 => \N__14601\,
            in1 => \N__14635\,
            in2 => \N__14548\,
            in3 => \N__14050\,
            lcout => \Lab_UT.m34_ns\,
            ltout => \Lab_UT.m34_ns_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIM00A3_3_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__14041\,
            in1 => \N__14546\,
            in2 => \N__14020\,
            in3 => \N__14007\,
            lcout => \Lab_UT.dictrl.next_state_set_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011000000110"
        )
    port map (
            in0 => \N__17219\,
            in1 => \N__14917\,
            in2 => \N__17365\,
            in3 => \N__13990\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__14918\,
            in1 => \N__17335\,
            in2 => \N__13954\,
            in3 => \N__17292\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13951\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18038\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__14496\,
            in1 => \N__15593\,
            in2 => \N__15640\,
            in3 => \N__15565\,
            lcout => \Lab_UT.dictrl.next_state_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18032\,
            ce => \N__14388\,
            sr => \N__13906\
        );

    \Lab_UT.didp.m41_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__14529\,
            in1 => \N__14630\,
            in2 => \_gnd_net_\,
            in3 => \N__16780\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.N_164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m42_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__16781\,
            in1 => \N__14597\,
            in2 => \N__13897\,
            in3 => \N__17015\,
            lcout => \Lab_UT.m42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__15488\,
            in1 => \N__14914\,
            in2 => \_gnd_net_\,
            in3 => \N__17214\,
            lcout => \Lab_UT.didp.countrce4.N_88_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_RNICI8U_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__17016\,
            in1 => \N__14631\,
            in2 => \N__14605\,
            in3 => \N__16782\,
            lcout => \Lab_UT.LdMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__15489\,
            in1 => \N__14343\,
            in2 => \_gnd_net_\,
            in3 => \N__17215\,
            lcout => \Lab_UT.didp.un31_reset_i_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__14418\,
            in1 => \N__16897\,
            in2 => \N__14470\,
            in3 => \N__14449\,
            lcout => \Lab_UT.state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_0_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__14448\,
            in1 => \N__14465\,
            in2 => \N__16912\,
            in3 => \N__14417\,
            lcout => \Lab_UT.state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_ret_3_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010001111110011"
        )
    port map (
            in0 => \N__14263\,
            in1 => \N__14286\,
            in2 => \N__16913\,
            in3 => \N__14310\,
            lcout => \Lab_UT.dictrl.state_i_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_0_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__14309\,
            in1 => \N__16901\,
            in2 => \N__14287\,
            in3 => \N__14262\,
            lcout => \Lab_UT.state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17041\,
            in1 => \N__16755\,
            in2 => \_gnd_net_\,
            in3 => \N__17162\,
            lcout => \Lab_UT.Run\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14086\,
            in2 => \_gnd_net_\,
            in3 => \N__14074\,
            lcout => \Lab_UT.dictrl.dicRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_0_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__16896\,
            in1 => \N__15570\,
            in2 => \N__15600\,
            in3 => \N__15638\,
            lcout => \Lab_UT.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18027\,
            ce => 'H',
            sr => \N__17812\
        );

    \Lab_UT.dictrl.state_ret_3_RNI2T7U_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14627\,
            in2 => \_gnd_net_\,
            in3 => \N__17042\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_state_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNITFCD1_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__17080\,
            in2 => \N__14644\,
            in3 => \N__17019\,
            lcout => \Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m37_ns_1_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111110"
        )
    port map (
            in0 => \N__14583\,
            in1 => \N__14629\,
            in2 => \N__14542\,
            in3 => \N__16759\,
            lcout => \Lab_UT.didp.m37_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_RNI0P1V_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111011111"
        )
    port map (
            in0 => \N__14628\,
            in1 => \N__14582\,
            in2 => \N__14541\,
            in3 => \N__17163\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.un1_state_24_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_RNIRB6E1_1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000001111"
        )
    port map (
            in0 => \N__17020\,
            in1 => \N__17079\,
            in2 => \N__14500\,
            in3 => \N__16761\,
            lcout => \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16914\,
            in2 => \_gnd_net_\,
            in3 => \N__17853\,
            lcout => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0\,
            ltout => \Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__14469\,
            in1 => \N__14447\,
            in2 => \N__14422\,
            in3 => \N__14419\,
            lcout => \Lab_UT.dictrl.next_state_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18023\,
            ce => \N__14387\,
            sr => \N__14755\
        );

    \Lab_UT.dispString.dOut_5_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011000100"
        )
    port map (
            in0 => \N__15375\,
            in1 => \N__15163\,
            in2 => \N__18277\,
            in3 => \N__15270\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m28_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__15371\,
            in1 => \N__15155\,
            in2 => \_gnd_net_\,
            in3 => \N__15266\,
            lcout => \Lab_UT.un29_dOutP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011111000111"
        )
    port map (
            in0 => \N__15268\,
            in1 => \N__15373\,
            in2 => \N__15173\,
            in3 => \N__16174\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000001000000"
        )
    port map (
            in0 => \N__15028\,
            in1 => \N__15412\,
            in2 => \N__14710\,
            in3 => \N__16646\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__17659\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14831\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000100"
        )
    port map (
            in0 => \N__15374\,
            in1 => \N__15162\,
            in2 => \N__16723\,
            in3 => \N__15269\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111101111"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__15372\,
            in2 => \N__15172\,
            in3 => \N__15813\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__15402\,
            in1 => \N__16419\,
            in2 => \N__15030\,
            in3 => \N__17493\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.G_64_a0_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14845\,
            in1 => \N__17404\,
            in2 => \N__15487\,
            in3 => \N__15073\,
            lcout => \Lab_UT.alarmMatch\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100101"
        )
    port map (
            in0 => \N__15242\,
            in1 => \N__14761\,
            in2 => \N__15178\,
            in3 => \N__15726\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15401\,
            in2 => \N__15040\,
            in3 => \N__17230\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__15403\,
            in1 => \N__16576\,
            in2 => \N__15031\,
            in3 => \N__14942\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15004\,
            in2 => \N__14998\,
            in3 => \N__14953\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18075\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__16321\,
            in1 => \N__14838\,
            in2 => \N__15087\,
            in3 => \N__14814\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.G_64_a0_1_0_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14919\,
            in1 => \N__16320\,
            in2 => \N__16173\,
            in3 => \N__16250\,
            lcout => \Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110001"
        )
    port map (
            in0 => \N__14839\,
            in1 => \N__14815\,
            in2 => \N__15088\,
            in3 => \N__17559\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__14806\,
            in1 => \_gnd_net_\,
            in2 => \N__14797\,
            in3 => \N__15832\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18262\,
            lcout => \Lab_UT.alarmcharZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18261\,
            in2 => \_gnd_net_\,
            in3 => \N__18317\,
            lcout => OPEN,
            ltout => \Lab_UT.alarmchar9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_2_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15091\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmcharZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_1_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18127\,
            in2 => \_gnd_net_\,
            in3 => \N__18318\,
            lcout => \Lab_UT.alarmcharZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18069\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment3.un1_num_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15943\,
            in1 => \N__15774\,
            in2 => \N__16047\,
            in3 => \N__15698\,
            lcout => \Lab_UT.zero\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__15699\,
            in1 => \N__16026\,
            in2 => \N__15794\,
            in3 => \N__15945\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.qPone_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__16698\,
            in1 => \N__16031\,
            in2 => \N__15064\,
            in3 => \N__15057\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__15701\,
            in1 => \N__15058\,
            in2 => \N__15795\,
            in3 => \N__16699\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101010101"
        )
    port map (
            in0 => \N__15944\,
            in1 => \N__15778\,
            in2 => \_gnd_net_\,
            in3 => \N__15700\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.N_79_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100000100"
        )
    port map (
            in0 => \N__15056\,
            in1 => \N__16697\,
            in2 => \N__15061\,
            in3 => \N__15946\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16696\,
            in1 => \N__15055\,
            in2 => \_gnd_net_\,
            in3 => \N__15702\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__15265\,
            in1 => \N__15147\,
            in2 => \N__15376\,
            in3 => \N__16025\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNI36SS_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15773\,
            in2 => \_gnd_net_\,
            in3 => \N__15692\,
            lcout => \Lab_UT.N_207\,
            ltout => \Lab_UT.N_207_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIIKFH3_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15879\,
            in1 => \N__16027\,
            in2 => \N__15658\,
            in3 => \N__15953\,
            lcout => \Lab_UT.didp.q_RNIIKFH3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000110110101111"
        )
    port map (
            in0 => \N__16886\,
            in1 => \N__15639\,
            in2 => \N__15604\,
            in3 => \N__15574\,
            lcout => \Lab_UT.state_i_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18057\,
            ce => 'H',
            sr => \N__17809\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110011"
        )
    port map (
            in0 => \N__15541\,
            in1 => \N__15245\,
            in2 => \N__15985\,
            in3 => \N__15121\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001010000"
        )
    port map (
            in0 => \N__15393\,
            in1 => \_gnd_net_\,
            in2 => \N__15532\,
            in3 => \N__15525\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.m29_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__15339\,
            in1 => \N__15120\,
            in2 => \_gnd_net_\,
            in3 => \N__15244\,
            lcout => \Lab_UT.un3_dOutP\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15247\,
            in1 => \N__15312\,
            in2 => \N__15148\,
            in3 => \N__15340\,
            lcout => \Lab_UT.cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18057\,
            ce => 'H',
            sr => \N__17809\
        );

    \Lab_UT.dispString.cnt_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__15311\,
            in1 => \N__15122\,
            in2 => \_gnd_net_\,
            in3 => \N__15246\,
            lcout => \Lab_UT.cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18057\,
            ce => 'H',
            sr => \N__17809\
        );

    \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16312\,
            in2 => \_gnd_net_\,
            in3 => \N__16229\,
            lcout => \Lab_UT.N_204\,
            ltout => \Lab_UT.N_204_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_2_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16681\,
            in1 => \N__16171\,
            in2 => \N__16702\,
            in3 => \N__17558\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18051\,
            ce => 'H',
            sr => \N__17127\
        );

    \Lab_UT.didp.reset_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16680\,
            in2 => \_gnd_net_\,
            in3 => \N__17856\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18051\,
            ce => 'H',
            sr => \N__17127\
        );

    \Lab_UT.didp.ce_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16618\,
            in1 => \N__16558\,
            in2 => \N__16482\,
            in3 => \N__16398\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18051\,
            ce => 'H',
            sr => \N__17127\
        );

    \Lab_UT.didp.countrce2.q_RNI1S78_0_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16313\,
            in2 => \_gnd_net_\,
            in3 => \N__16230\,
            lcout => \Lab_UT.didp.countrce2.three_2\,
            ltout => \Lab_UT.didp.countrce2.three_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__16161\,
            in1 => \_gnd_net_\,
            in2 => \N__16090\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.countrce2.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_3_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__16048\,
            in1 => \N__15968\,
            in2 => \N__15880\,
            in3 => \N__15894\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18051\,
            ce => 'H',
            sr => \N__17127\
        );

    \Lab_UT.didp.reset_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17857\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15875\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18051\,
            ce => 'H',
            sr => \N__17127\
        );

    \Lab_UT.bcd2segment4.G_64_a0_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__17547\,
            in1 => \N__17471\,
            in2 => \_gnd_net_\,
            in3 => \N__17201\,
            lcout => \Lab_UT.bcd2segment4.G_64_a0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__17395\,
            in1 => \N__17202\,
            in2 => \_gnd_net_\,
            in3 => \N__17364\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__17203\,
            in1 => \N__17340\,
            in2 => \N__17296\,
            in3 => \N__17275\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18046\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17044\,
            in1 => \N__16783\,
            in2 => \_gnd_net_\,
            in3 => \N__17164\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18039\,
            ce => 'H',
            sr => \N__17128\
        );

    \Lab_UT.dictrl.state_ret_3_RNIDH8U_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__17078\,
            in1 => \N__17043\,
            in2 => \N__17017\,
            in3 => \N__16772\,
            lcout => \Lab_UT.dictrl.state_ret_3_RNIDH8UZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__16963\,
            in1 => \N__16932\,
            in2 => \N__16918\,
            in3 => \N__16810\,
            lcout => \Lab_UT.state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18028\,
            ce => 'H',
            sr => \N__17813\
        );

    \Lab_UT.alarmchar_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18373\,
            lcout => \Lab_UT.alarmcharZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18126\,
            in2 => \_gnd_net_\,
            in3 => \N__18316\,
            lcout => OPEN,
            ltout => \Lab_UT.alarmchar_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.alarmchar_6_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17662\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmcharZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000101"
        )
    port map (
            in0 => \N__18330\,
            in1 => \N__18217\,
            in2 => \N__18190\,
            in3 => \N__18353\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1\,
            ltout => \Lab_UT.dictrl.next_alarmstate_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_3_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__17646\,
            in1 => \_gnd_net_\,
            in2 => \N__17650\,
            in3 => \N__17587\,
            lcout => \Lab_UT.un1_next_alarmstate21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.G_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__18305\,
            in1 => \N__18354\,
            in2 => \N__18232\,
            in3 => \N__17645\,
            lcout => OPEN,
            ltout => \Lab_UT.G_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_0_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__17581\,
            in1 => \_gnd_net_\,
            in2 => \N__17593\,
            in3 => \N__18216\,
            lcout => \Lab_UT.dictrl.next_alarmstate_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18086\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__17566\,
            in1 => \N__18352\,
            in2 => \N__18260\,
            in3 => \N__17580\,
            lcout => \Lab_UT.dictrl.next_alarmstate_1_0\,
            ltout => \Lab_UT.dictrl.next_alarmstate_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18215\,
            in2 => \N__17590\,
            in3 => \N__18181\,
            lcout => \Lab_UT.dictrl.next_alarmstateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__18304\,
            in1 => \N__18119\,
            in2 => \_gnd_net_\,
            in3 => \N__17579\,
            lcout => \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18118\,
            in2 => \_gnd_net_\,
            in3 => \N__18303\,
            lcout => \Lab_UT.dictrl.idle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_1_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__18188\,
            in1 => \N__18146\,
            in2 => \_gnd_net_\,
            in3 => \N__18363\,
            lcout => \Lab_UT.alarmchar10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18077\,
            ce => 'H',
            sr => \N__17810\
        );

    \Lab_UT.dictrl.alarmstate_ret_2_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__18364\,
            in1 => \N__18189\,
            in2 => \_gnd_net_\,
            in3 => \N__18148\,
            lcout => \Lab_UT.alarmchar10_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18077\,
            ce => 'H',
            sr => \N__17810\
        );

    \Lab_UT.dictrl.alarmstate_0_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__18218\,
            in1 => \N__18185\,
            in2 => \_gnd_net_\,
            in3 => \N__18145\,
            lcout => \Lab_UT.alarmstate_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18077\,
            ce => 'H',
            sr => \N__17810\
        );

    \Lab_UT.dictrl.alarmstate_0_1_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__18187\,
            in1 => \N__18355\,
            in2 => \N__18223\,
            in3 => \N__18331\,
            lcout => \Lab_UT.alarmstate_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18077\,
            ce => 'H',
            sr => \N__17810\
        );

    \Lab_UT.alarmchar_5_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18283\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.alarmcharZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18070\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.bcd2segment4.G_1_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18180\,
            in2 => \_gnd_net_\,
            in3 => \N__18253\,
            lcout => \Lab_UT.bcd2segment4.GZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_ret_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__18222\,
            in1 => \N__18186\,
            in2 => \_gnd_net_\,
            in3 => \N__18147\,
            lcout => \Lab_UT.dictrl.alarmstate_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18087\,
            ce => 'H',
            sr => \N__17811\
        );
end \INTERFACE\;
