-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     May 20 2019 23:10:54

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "latticehx1k" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of latticehx1k
entity latticehx1k is
port (
    led : out std_logic_vector(4 downto 0);
    o_serial_data : out std_logic;
    to_ir : out std_logic;
    sd : out std_logic;
    from_pc : in std_logic;
    clk_in : in std_logic);
end latticehx1k;

-- Architecture of latticehx1k
-- View name is \INTERFACE\
architecture \INTERFACE\ of latticehx1k is

signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26840\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26824\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26822\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26813\ : std_logic;
signal \N__26806\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26804\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26795\ : std_logic;
signal \N__26788\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26786\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26777\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26738\ : std_logic;
signal \N__26735\ : std_logic;
signal \N__26732\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26725\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26722\ : std_logic;
signal \N__26719\ : std_logic;
signal \N__26716\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26693\ : std_logic;
signal \N__26690\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26687\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26681\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26639\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26623\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26617\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26594\ : std_logic;
signal \N__26591\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26572\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26566\ : std_logic;
signal \N__26563\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26537\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26531\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26521\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26497\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26489\ : std_logic;
signal \N__26486\ : std_logic;
signal \N__26483\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26459\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26456\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26432\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26417\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26395\ : std_logic;
signal \N__26392\ : std_logic;
signal \N__26391\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26371\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26359\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26350\ : std_logic;
signal \N__26349\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26309\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26294\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26282\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26267\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26256\ : std_logic;
signal \N__26253\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26243\ : std_logic;
signal \N__26238\ : std_logic;
signal \N__26235\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26231\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26228\ : std_logic;
signal \N__26223\ : std_logic;
signal \N__26216\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26205\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26201\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26198\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26196\ : std_logic;
signal \N__26195\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26193\ : std_logic;
signal \N__26192\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26190\ : std_logic;
signal \N__26189\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26180\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26177\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26174\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26171\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26168\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26165\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26162\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26159\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26156\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26154\ : std_logic;
signal \N__26153\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26151\ : std_logic;
signal \N__26150\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26146\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26144\ : std_logic;
signal \N__26143\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26141\ : std_logic;
signal \N__26140\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26138\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26135\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26132\ : std_logic;
signal \N__26131\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26129\ : std_logic;
signal \N__26128\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26126\ : std_logic;
signal \N__26125\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26123\ : std_logic;
signal \N__26122\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26120\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26117\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25903\ : std_logic;
signal \N__25900\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25891\ : std_logic;
signal \N__25888\ : std_logic;
signal \N__25881\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25878\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25875\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25849\ : std_logic;
signal \N__25846\ : std_logic;
signal \N__25843\ : std_logic;
signal \N__25842\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25836\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25833\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25830\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25827\ : std_logic;
signal \N__25826\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25823\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25820\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25818\ : std_logic;
signal \N__25817\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25815\ : std_logic;
signal \N__25814\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25811\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25806\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25801\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25790\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25776\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25772\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25767\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25611\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25599\ : std_logic;
signal \N__25598\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25589\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25586\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25580\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25559\ : std_logic;
signal \N__25558\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25556\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25553\ : std_logic;
signal \N__25550\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25521\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25513\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25502\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25494\ : std_logic;
signal \N__25493\ : std_logic;
signal \N__25490\ : std_logic;
signal \N__25485\ : std_logic;
signal \N__25482\ : std_logic;
signal \N__25481\ : std_logic;
signal \N__25478\ : std_logic;
signal \N__25475\ : std_logic;
signal \N__25470\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25439\ : std_logic;
signal \N__25434\ : std_logic;
signal \N__25431\ : std_logic;
signal \N__25426\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25409\ : std_logic;
signal \N__25408\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25394\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25365\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25338\ : std_logic;
signal \N__25335\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25272\ : std_logic;
signal \N__25269\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25257\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25206\ : std_logic;
signal \N__25203\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25188\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25183\ : std_logic;
signal \N__25176\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25170\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25167\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25131\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25116\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25104\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25089\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25079\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25061\ : std_logic;
signal \N__25058\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25043\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25031\ : std_logic;
signal \N__25030\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24960\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24933\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24927\ : std_logic;
signal \N__24924\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24918\ : std_logic;
signal \N__24909\ : std_logic;
signal \N__24906\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24897\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24890\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24878\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24872\ : std_logic;
signal \N__24869\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24824\ : std_logic;
signal \N__24821\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24751\ : std_logic;
signal \N__24748\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24720\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24703\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24695\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24692\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24673\ : std_logic;
signal \N__24670\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24652\ : std_logic;
signal \N__24649\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24622\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24591\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24578\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24528\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24481\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24466\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24460\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24458\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24401\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24383\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24368\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24362\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24348\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24341\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24321\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24313\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24308\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24305\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24272\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24254\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24243\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24087\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24062\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24053\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24051\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24035\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24015\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24008\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23997\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23981\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23972\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23925\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23909\ : std_logic;
signal \N__23906\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23669\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23642\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23616\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23580\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23562\ : std_logic;
signal \N__23555\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23534\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23502\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23435\ : std_logic;
signal \N__23432\ : std_logic;
signal \N__23429\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23411\ : std_logic;
signal \N__23408\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23329\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23291\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23123\ : std_logic;
signal \N__23120\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23066\ : std_logic;
signal \N__23063\ : std_logic;
signal \N__23060\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23036\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23013\ : std_logic;
signal \N__23010\ : std_logic;
signal \N__23007\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22967\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22940\ : std_logic;
signal \N__22937\ : std_logic;
signal \N__22934\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22907\ : std_logic;
signal \N__22904\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22878\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22851\ : std_logic;
signal \N__22848\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22817\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22814\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22781\ : std_logic;
signal \N__22778\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22766\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22742\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22718\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22686\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22647\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22618\ : std_logic;
signal \N__22615\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22508\ : std_logic;
signal \N__22505\ : std_logic;
signal \N__22502\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22473\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22379\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22370\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22304\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22268\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22245\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22213\ : std_logic;
signal \N__22210\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22185\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22157\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22148\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22145\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22065\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22059\ : std_logic;
signal \N__22056\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21971\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21961\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21906\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21876\ : std_logic;
signal \N__21873\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21858\ : std_logic;
signal \N__21855\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21783\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21740\ : std_logic;
signal \N__21737\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21714\ : std_logic;
signal \N__21711\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21690\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21651\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21624\ : std_logic;
signal \N__21621\ : std_logic;
signal \N__21620\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21588\ : std_logic;
signal \N__21585\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21543\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21531\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21525\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21504\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21498\ : std_logic;
signal \N__21495\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21422\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21410\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21384\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21375\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21333\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21255\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21249\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21222\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21162\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21133\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21031\ : std_logic;
signal \N__21028\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21015\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21012\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20921\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20904\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20888\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20882\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20868\ : std_logic;
signal \N__20865\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20859\ : std_logic;
signal \N__20854\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20844\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20823\ : std_logic;
signal \N__20820\ : std_logic;
signal \N__20817\ : std_logic;
signal \N__20814\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20799\ : std_logic;
signal \N__20796\ : std_logic;
signal \N__20793\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20789\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20775\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20763\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20760\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20756\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20754\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20744\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20717\ : std_logic;
signal \N__20714\ : std_logic;
signal \N__20711\ : std_logic;
signal \N__20706\ : std_logic;
signal \N__20691\ : std_logic;
signal \N__20688\ : std_logic;
signal \N__20685\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20664\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20604\ : std_logic;
signal \N__20601\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20532\ : std_logic;
signal \N__20529\ : std_logic;
signal \N__20526\ : std_logic;
signal \N__20523\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20499\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20489\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20481\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20442\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20433\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20423\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20408\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20402\ : std_logic;
signal \N__20399\ : std_logic;
signal \N__20396\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20387\ : std_logic;
signal \N__20384\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20375\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20360\ : std_logic;
signal \N__20357\ : std_logic;
signal \N__20354\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20345\ : std_logic;
signal \N__20342\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20324\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20321\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20318\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20269\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20246\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20207\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20183\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20123\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20092\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20090\ : std_logic;
signal \N__20087\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20078\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20075\ : std_logic;
signal \N__20072\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20015\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20009\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19961\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19958\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19914\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19845\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19832\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19805\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19778\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19711\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19688\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19665\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19655\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19619\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19590\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19554\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19538\ : std_logic;
signal \N__19535\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19485\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19464\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19455\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19449\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19446\ : std_logic;
signal \N__19445\ : std_logic;
signal \N__19440\ : std_logic;
signal \N__19439\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19425\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19385\ : std_logic;
signal \N__19380\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19305\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19295\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19194\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19164\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19091\ : std_logic;
signal \N__19088\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19041\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19020\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__18999\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18945\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18935\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18910\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18877\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18875\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18869\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18850\ : std_logic;
signal \N__18847\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18731\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18725\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18716\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18689\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18676\ : std_logic;
signal \N__18673\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18650\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18641\ : std_logic;
signal \N__18638\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18617\ : std_logic;
signal \N__18614\ : std_logic;
signal \N__18611\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18605\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18586\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18560\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18548\ : std_logic;
signal \N__18545\ : std_logic;
signal \N__18542\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18506\ : std_logic;
signal \N__18503\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18425\ : std_logic;
signal \N__18422\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18395\ : std_logic;
signal \N__18392\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18368\ : std_logic;
signal \N__18365\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18353\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18347\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18323\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18297\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18272\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18254\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18233\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18221\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18182\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18164\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18152\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18137\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18079\ : std_logic;
signal \N__18076\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18032\ : std_logic;
signal \N__18029\ : std_logic;
signal \N__18026\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18014\ : std_logic;
signal \N__18011\ : std_logic;
signal \N__18008\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17999\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17964\ : std_logic;
signal \N__17961\ : std_logic;
signal \N__17958\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17939\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17936\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17904\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17901\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17874\ : std_logic;
signal \N__17871\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17864\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17825\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17799\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17772\ : std_logic;
signal \N__17769\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17751\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17739\ : std_logic;
signal \N__17736\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17727\ : std_logic;
signal \N__17724\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17718\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17682\ : std_logic;
signal \N__17679\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17664\ : std_logic;
signal \N__17661\ : std_logic;
signal \N__17658\ : std_logic;
signal \N__17655\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17634\ : std_logic;
signal \N__17631\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17580\ : std_logic;
signal \N__17577\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17552\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17540\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17484\ : std_logic;
signal \N__17481\ : std_logic;
signal \N__17478\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17465\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17439\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17421\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17393\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17385\ : std_logic;
signal \N__17382\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17345\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17339\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17295\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17286\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17147\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17046\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17042\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17012\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16835\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16832\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16829\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16796\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16767\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16733\ : std_logic;
signal \N__16730\ : std_logic;
signal \N__16727\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16656\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16652\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16643\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16616\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16586\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16517\ : std_logic;
signal \N__16514\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16481\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16434\ : std_logic;
signal \N__16431\ : std_logic;
signal \N__16428\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16424\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16379\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16376\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16337\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16328\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16307\ : std_logic;
signal \N__16304\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16253\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16250\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16241\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16238\ : std_logic;
signal \N__16235\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16226\ : std_logic;
signal \N__16223\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16130\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16109\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16103\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16094\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15999\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15989\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15962\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15935\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15926\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15851\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15805\ : std_logic;
signal \N__15802\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15772\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15750\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15729\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15723\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15717\ : std_logic;
signal \N__15714\ : std_logic;
signal \N__15711\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15702\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15666\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15632\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15584\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15374\ : std_logic;
signal \N__15371\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15317\ : std_logic;
signal \N__15314\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15197\ : std_logic;
signal \N__15194\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15130\ : std_logic;
signal \N__15125\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15077\ : std_logic;
signal \N__15074\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15068\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14952\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14719\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14712\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14691\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14427\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14369\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14258\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14137\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14045\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13931\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13916\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13886\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13703\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13688\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13329\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13084\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12833\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12173\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal clk_in_c : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \uu0.l_precountZ0Z_3\ : std_logic;
signal \uu0.l_precountZ0Z_1\ : std_logic;
signal \uu0.l_precountZ0Z_2\ : std_logic;
signal \uu0.l_precountZ0Z_0\ : std_logic;
signal \uu0.un4_l_count_14_cascade_\ : std_logic;
signal \uu0.un154_ci_9_cascade_\ : std_logic;
signal \uu0.un187_ci_1_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_14\ : std_logic;
signal \uu0.l_countZ0Z_15\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.un2_counter_cry_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_6\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_tx.Z_baudgen.ser_clk_4\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_tx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \resetGen_reset_count_2_2_cascade_\ : std_logic;
signal \resetGen_reset_count_2\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2_THRU_CO\ : std_logic;
signal \buart.Z_rx.bitcount_cry_2\ : std_logic;
signal \buart.Z_rx.bitcount_cry_3\ : std_logic;
signal \Lab_UT_dispString_m103_ns_1_cascade_\ : std_logic;
signal \buart.Z_rx.bitcount_cry_0_THRU_CO\ : std_logic;
signal \buart__rx_N_27_0_i_cascade_\ : std_logic;
signal \N_179\ : std_logic;
signal \uart_RXD\ : std_logic;
signal \Lab_UT.dispString.N_115_mux\ : std_logic;
signal \Lab_UT.dispString.N_115_mux_cascade_\ : std_logic;
signal \buart__rx_bitcount_1\ : std_logic;
signal \buart__rx_bitcount_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_177\ : std_logic;
signal \buart__rx_ser_clk_cascade_\ : std_logic;
signal \buart__rx_bitcount_0\ : std_logic;
signal \buart__rx_sample\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_0\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_1\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_3\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_2\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_3\ : std_logic;
signal \buart__rx_ser_clk\ : std_logic;
signal \buart.Z_rx.Z_baudgen.un5_counter_cry_4\ : std_logic;
signal \buart.Z_rx.Z_baudgen.counterZ0Z_5\ : std_logic;
signal \uu2.r_data_wire_0\ : std_logic;
signal \uu2.r_data_wire_1\ : std_logic;
signal \uu2.r_data_wire_2\ : std_logic;
signal \uu2.r_data_wire_3\ : std_logic;
signal \uu2.r_data_wire_4\ : std_logic;
signal \uu2.r_data_wire_5\ : std_logic;
signal \uu2.r_data_wire_6\ : std_logic;
signal \uu2.r_data_wire_7\ : std_logic;
signal \INVuu2.r_data_reg_0C_net\ : std_logic;
signal vbuf_tx_data_0 : std_logic;
signal \buart.Z_tx.shifterZ0Z_1\ : std_logic;
signal \buart.Z_tx.shifterZ0Z_0\ : std_logic;
signal o_serial_data_c : std_logic;
signal vbuf_tx_data_1 : std_logic;
signal \buart.Z_tx.shifterZ0Z_2\ : std_logic;
signal vbuf_tx_data_2 : std_logic;
signal \buart.Z_tx.shifterZ0Z_3\ : std_logic;
signal vbuf_tx_data_3 : std_logic;
signal \buart.Z_tx.shifterZ0Z_4\ : std_logic;
signal vbuf_tx_data_4 : std_logic;
signal \buart.Z_tx.shifterZ0Z_5\ : std_logic;
signal \uu0.un44_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_0\ : std_logic;
signal \uu0.l_countZ0Z_1\ : std_logic;
signal \uu0.un66_ci_cascade_\ : std_logic;
signal \uu0.un110_ci_cascade_\ : std_logic;
signal \uu0.l_countZ0Z_10\ : std_logic;
signal \uu0.l_countZ0Z_8\ : std_logic;
signal \uu0.l_countZ0Z_9\ : std_logic;
signal \uu0.l_countZ0Z_17\ : std_logic;
signal \uu0.un198_ci_2\ : std_logic;
signal \uu0.l_countZ0Z_16\ : std_logic;
signal \uu0.un44_ci\ : std_logic;
signal \uu0.l_countZ0Z_2\ : std_logic;
signal \uu0.l_countZ0Z_3\ : std_logic;
signal \uu0.un66_ci\ : std_logic;
signal \uu0.l_countZ0Z_7\ : std_logic;
signal \uu0.un220_ci\ : std_logic;
signal \uu0.un143_ci_0\ : std_logic;
signal \uu0.l_countZ0Z_11\ : std_logic;
signal \uu0.l_countZ0Z_18\ : std_logic;
signal \uu0.un4_l_count_11\ : std_logic;
signal \uu0.un4_l_count_12\ : std_logic;
signal \uu0.un4_l_count_13\ : std_logic;
signal \uu0.un4_l_count_16_cascade_\ : std_logic;
signal \uu0.un4_l_count_18\ : std_logic;
signal \uu0.un110_ci\ : std_logic;
signal \uu0.un4_l_count_0_cascade_\ : std_logic;
signal \uu0.un11_l_count_i_g\ : std_logic;
signal vbuf_tx_data_5 : std_logic;
signal \buart.Z_tx.shifterZ0Z_6\ : std_logic;
signal vbuf_tx_data_6 : std_logic;
signal \buart.Z_tx.shifterZ0Z_7\ : std_logic;
signal vbuf_tx_data_7 : std_logic;
signal \buart.Z_tx.shifterZ0Z_8\ : std_logic;
signal \buart.Z_tx.un1_uart_wr_i_0_i\ : std_logic;
signal \uu0.l_countZ0Z_13\ : std_logic;
signal \uu0.un4_l_count_0_8\ : std_logic;
signal \uu0.un154_ci_9\ : std_logic;
signal \uu0.l_countZ0Z_12\ : std_logic;
signal \uu0.un165_ci_0\ : std_logic;
signal \resetGen_reset_count_1\ : std_logic;
signal \N_107\ : std_logic;
signal \m72_cascade_\ : std_logic;
signal \N_105\ : std_logic;
signal \resetGen.reset_countZ0Z_3\ : std_logic;
signal \resetGen_reset_count_4\ : std_logic;
signal \resetGen_reset_count_0\ : std_logic;
signal \buart__rx_hh_0\ : std_logic;
signal \Lab_UT.dictrl.g0_69_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_0_3_1\ : std_logic;
signal \Lab_UT.dictrl.g1_5_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_61_1\ : std_logic;
signal \Lab_UT.dictrl.g1_7_0\ : std_logic;
signal \Lab_UT.dictrl.N_1792_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1451_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a5_2_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a5_2_5\ : std_logic;
signal \Lab_UT.dictrl.g0_5_3\ : std_logic;
signal \Lab_UT.dictrl.g0_5_4\ : std_logic;
signal \Lab_UT.dictrl.g1_6_0\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3\ : std_logic;
signal \uu2.vbuf_raddr.un426_ci_3_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_8\ : std_logic;
signal \uu2.r_addrZ0Z_7\ : std_logic;
signal \uu2.vbuf_raddr.un448_ci_0\ : std_logic;
signal \uu2.un404_ci_0_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_6\ : std_logic;
signal \uu2.r_addrZ0Z_3\ : std_logic;
signal \uu2.r_addrZ0Z_2\ : std_logic;
signal \uu2.r_addrZ0Z_1\ : std_logic;
signal \uu2.trig_rd_is_det_0\ : std_logic;
signal \uu2.trig_rd_is_det_cascade_\ : std_logic;
signal \uu2.r_addrZ0Z_0\ : std_logic;
signal \uu2.trig_rd_detZ0Z_1\ : std_logic;
signal \uu2.trig_rd_detZ0Z_0\ : std_logic;
signal \uu2.un1_l_count_1_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_0_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_3\ : std_logic;
signal \uu2.l_countZ0Z_3\ : std_logic;
signal \uu2.l_countZ0Z_2\ : std_logic;
signal \uu2.un306_ci_cascade_\ : std_logic;
signal \uu2.un1_l_count_1_2_0\ : std_logic;
signal \uu2.l_countZ0Z_5\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3_cascade_\ : std_logic;
signal \uu2.un1_l_count_2_0\ : std_logic;
signal \uu2.un350_ci_cascade_\ : std_logic;
signal \uu2.l_countZ0Z_4\ : std_logic;
signal \uu2.l_countZ0Z_9\ : std_logic;
signal \uu2.un1_l_count_2_2\ : std_logic;
signal \uu2.un306_ci\ : std_logic;
signal \uu2.vbuf_count.un328_ci_3\ : std_logic;
signal \uu2.l_countZ0Z_6\ : std_logic;
signal \uu2.l_countZ0Z_7\ : std_logic;
signal \uu2.un350_ci\ : std_logic;
signal \uu2.l_countZ0Z_8\ : std_logic;
signal \uu0.un4_l_count_0\ : std_logic;
signal \uu0.un11_l_count_i\ : std_logic;
signal \uu0.delay_lineZ0Z_0\ : std_logic;
signal \uu0.delay_lineZ0Z_1\ : std_logic;
signal \buart.Z_tx.un1_bitcount_c3_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_3\ : std_logic;
signal \buart.Z_tx.uart_busy_0_0\ : std_logic;
signal \buart.Z_tx.ser_clk\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_1\ : std_logic;
signal \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\ : std_logic;
signal \buart.Z_tx.bitcountZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g0_12_o6_2_2\ : std_logic;
signal \Lab_UT.dictrl.N_13_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_10Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.m34_4Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_\ : std_logic;
signal \buart__rx_hh_1\ : std_logic;
signal \Lab_UT.dictrl.m40Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_10_3\ : std_logic;
signal \Lab_UT.dictrl.N_5_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_9Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.g1_4\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_2435_0\ : std_logic;
signal \Lab_UT.dictrl.g1_5_0\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_0\ : std_logic;
signal \Lab_UT.dictrl.g0_16_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_2446_1\ : std_logic;
signal \uu2.mem0.w_addr_0\ : std_logic;
signal clk : std_logic;
signal \uu2.vram_wr_en_0_iZ0\ : std_logic;
signal \uu2.mem0.w_addr_1\ : std_logic;
signal \uu2.mem0.w_addr_2\ : std_logic;
signal \INVuu2.w_addr_user_1C_net\ : std_logic;
signal \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\ : std_logic;
signal \uu2.w_addr_userZ0Z_0\ : std_logic;
signal \uu2.un426_ci_3_cascade_\ : std_logic;
signal \INVuu2.w_addr_user_nesr_8C_net\ : std_logic;
signal \uu2.r_addrZ0Z_4\ : std_logic;
signal \uu2.un404_ci_0\ : std_logic;
signal \uu2.trig_rd_is_det\ : std_logic;
signal \uu2.r_addrZ0Z_5\ : std_logic;
signal \uu0.l_countZ0Z_5\ : std_logic;
signal \uu0.l_countZ0Z_4\ : std_logic;
signal \uu2.un284_ci\ : std_logic;
signal \uu2.l_countZ0Z_1\ : std_logic;
signal \uu2.l_countZ0Z_0\ : std_logic;
signal \uu2.un28_w_addr_user_i_0\ : std_logic;
signal \uu2.un1_l_count_1_0\ : std_logic;
signal vbuf_tx_data_rdy : std_logic;
signal \uu0.un88_ci_3\ : std_logic;
signal \uu0.l_countZ0Z_6\ : std_logic;
signal \uu0.un99_ci_0\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_2_tz_1\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_1_1_1\ : std_logic;
signal \Lab_UT.dispString.m74_ns_1\ : std_logic;
signal \Lab_UT.dispString.m77_ns_1\ : std_logic;
signal \Lab_UT.dispString.N_30_i\ : std_logic;
signal \Lab_UT.dispString.dOutP_0_iv_0_1\ : std_logic;
signal \uu0.sec_clkDZ0\ : std_logic;
signal \Lab_UT.alarmstate_1_0_i_1_cascade_\ : std_logic;
signal \G_215_cascade_\ : std_logic;
signal \G_214\ : std_logic;
signal \G_216\ : std_logic;
signal \G_214_cascade_\ : std_logic;
signal \Lab_UT.m57\ : std_logic;
signal \G_213\ : std_logic;
signal \G_215\ : std_logic;
signal \G_213_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m71Z0Z_0\ : std_logic;
signal \N_105_mux\ : std_logic;
signal \Lab_UT.dispString.N_186\ : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_3Z0Z_7\ : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_3_8_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_16\ : std_logic;
signal \N_10_2\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.g0_10_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m63_d_0_ns_1_1\ : std_logic;
signal \Lab_UT.dispString.N_112_mux\ : std_logic;
signal \Lab_UT.dictrl.m27_d_1\ : std_logic;
signal \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_17_i_a5_0_0\ : std_logic;
signal \buart.Z_rx.G_17_i_a5_2_5\ : std_logic;
signal \buart.Z_rx.G_17_i_a5_2_4\ : std_logic;
signal \G_17_i_a5_2_6_cascade_\ : std_logic;
signal bu_rx_data_fast_1 : std_logic;
signal bu_rx_data_fast_2 : std_logic;
signal \Lab_UT.dictrl.g2_0_3_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_0\ : std_logic;
signal bu_rx_data_1_rep1 : std_logic;
signal bu_rx_data_2_rep1 : std_logic;
signal \Lab_UT.dispString.m107_eZ0Z_3\ : std_logic;
signal bu_rx_data_fast_5 : std_logic;
signal \Lab_UT.dictrl.N_10_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_17_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_\ : std_logic;
signal \N_22\ : std_logic;
signal \Lab_UT.dictrl.N_1105_0\ : std_logic;
signal bu_rx_data_fast_7 : std_logic;
signal \Lab_UT.dictrl.N_10_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_1_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_1_a6_3_2\ : std_logic;
signal bu_rx_data_fast_3 : std_logic;
signal \Lab_UT.dictrl.N_7_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.G_17_i_a5_1\ : std_logic;
signal \uu2.mem0.N_66_i\ : std_logic;
signal \uu2.mem0.N_56_i\ : std_logic;
signal \uu2.N_95_mux\ : std_logic;
signal \uu2.N_96_mux_cascade_\ : std_logic;
signal \uu2.mem0.N_63_i\ : std_logic;
signal \uu2.mem0.N_69_i\ : std_logic;
signal \uu2.N_96_mux\ : std_logic;
signal \uu2.mem0.N_71_i\ : std_logic;
signal \uu2.mem0.N_91_mux\ : std_logic;
signal \uu2.mem0.N_50_i\ : std_logic;
signal \uu2.w_addr_userZ0Z_3\ : std_logic;
signal \uu2.mem0.w_addr_3\ : std_logic;
signal \uu2.mem0.w_addr_4\ : std_logic;
signal \uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_4C_net\ : std_logic;
signal \uu2.un1_w_user_lf_0_cascade_\ : std_logic;
signal \uu2.un1_w_user_lfZ0Z_4\ : std_logic;
signal \uu2.un1_w_user_lf_0\ : std_logic;
signal \L3_tx_data_5\ : std_logic;
signal \L3_tx_data_1\ : std_logic;
signal \L3_tx_data_4\ : std_logic;
signal \uu2.m35Z0Z_4_cascade_\ : std_logic;
signal \uu2.un1_w_user_cr_0_cascade_\ : std_logic;
signal \uu2.mem0.w_data_2\ : std_logic;
signal \Lab_UT.dispString.N_145\ : std_logic;
signal \Lab_UT.dispString.N_146_cascade_\ : std_logic;
signal \L3_tx_data_2\ : std_logic;
signal \L3_tx_data_0\ : std_logic;
signal \L3_tx_data_6\ : std_logic;
signal \Lab_UT.dispString.m82_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_156_cascade_\ : std_logic;
signal \L3_tx_data_3\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_2\ : std_logic;
signal \Lab_UT.dispString.b1_m_1\ : std_logic;
signal \Lab_UT.dispString.m67_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_143\ : std_logic;
signal \Lab_UT.dispString.N_23_0\ : std_logic;
signal \Lab_UT.dispString.N_158\ : std_logic;
signal \Lab_UT.dispString.m90_ns_1_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_164\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_0\ : std_logic;
signal \Lab_UT.dispString.cntZ0Z_1\ : std_logic;
signal \Lab_UT.dispString.N_166\ : std_logic;
signal \Lab_UT.dispString.N_167\ : std_logic;
signal \Lab_UT_dictrl_g1_0_3\ : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_3_6\ : std_logic;
signal \Lab_UT.dictrl.N_10\ : std_logic;
signal \Lab_UT.dictrl.g0_12_1\ : std_logic;
signal \Lab_UT.dictrl.m15Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_8_0\ : std_logic;
signal \Lab_UT.dictrl.N_93_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_10_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_0_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_0_3\ : std_logic;
signal \Lab_UT.dictrl.m15Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_88_mux\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m53_d_1_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_45_cascade_\ : std_logic;
signal bu_rx_data_1_rep2 : std_logic;
signal \Lab_UT.dictrl.g2_0_3_1\ : std_logic;
signal bu_rx_data_2_rep2 : std_logic;
signal \Lab_UT_dictrl_m59_1\ : std_logic;
signal \Lab_UT.dictrl.m59_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_3_4\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_3_2\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_0_3\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_cascade_\ : std_logic;
signal bu_rx_data_fast_0 : std_logic;
signal bu_rx_data_fast_4 : std_logic;
signal bu_rx_data_3_rep1 : std_logic;
signal \Lab_UT.dictrl.g2_0_3_3\ : std_logic;
signal \Lab_UT.dictrl.g2_0_4_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m12Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_11_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0\ : std_logic;
signal \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_\ : std_logic;
signal bu_rx_data_fast_6 : std_logic;
signal \buart.Z_rx.sample_g\ : std_logic;
signal \Lab_UT.dictrl.N_100\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_8Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m63_d_0_ns_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_3Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.m67_am_1_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\ : std_logic;
signal \Lab_UT.dictrl.G_17_i_a5_0\ : std_logic;
signal \Lab_UT.dictrl.N_65\ : std_logic;
signal \Lab_UT.dictrl.N_65_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_101\ : std_logic;
signal \uu2.mem0.w_addr_5\ : std_logic;
signal \uu2.mem0.w_addr_6\ : std_logic;
signal \uu2.w_addr_userZ0Z_7\ : std_logic;
signal \uu2.mem0.w_addr_7\ : std_logic;
signal \uu2.N_91\ : std_logic;
signal \uu2.N_28_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_26_i_m2_1_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_20\ : std_logic;
signal \uu2.N_55_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_i7_mux_0\ : std_logic;
signal \uu2.N_406_cascade_\ : std_logic;
signal \uu2.bitmap_pmux\ : std_logic;
signal \uu2.bitmapZ0Z_40\ : std_logic;
signal \uu2.bitmapZ0Z_296\ : std_logic;
signal \uu2.N_207\ : std_logic;
signal \uu2.bitmapZ0Z_168\ : std_logic;
signal \uu2.N_195\ : std_logic;
signal \INVuu2.bitmap_296C_net\ : std_logic;
signal \uu2.bitmapZ0Z_66\ : std_logic;
signal \uu2.bitmapZ0Z_162\ : std_logic;
signal \uu2.bitmap_pmux_15_ns_1\ : std_logic;
signal \INVuu2.bitmap_66C_net\ : std_logic;
signal \o_One_Sec_Pulse\ : std_logic;
signal \uu2.bitmapZ0Z_111\ : std_logic;
signal \uu2.vram_rd_clkZ0\ : std_logic;
signal \uu2.bitmapZ0Z_194\ : std_logic;
signal \uu2.bitmapZ0Z_34\ : std_logic;
signal \uu2.bitmapZ0Z_290\ : std_logic;
signal \INVuu2.bitmap_111C_net\ : std_logic;
signal \Lab_UT.didp.regrce4.LdAMtens_0\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.di_AMtens_3\ : std_logic;
signal \Lab_UT.didp.countrce4.un20_qPone\ : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_0_1\ : std_logic;
signal \Lab_UT.dictrl.state_2_rep1\ : std_logic;
signal \Lab_UT.dictrl.N_62_1\ : std_logic;
signal \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.N_79\ : std_logic;
signal \Lab_UT.dictrl.state_i_4_1\ : std_logic;
signal \Lab_UT.dictrl.N_99\ : std_logic;
signal \buart__rx_bitcount_3\ : std_logic;
signal \buart__rx_valid_3\ : std_logic;
signal \Lab_UT.dictrl.g0_0_2_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1_0\ : std_logic;
signal \Lab_UT.dictrl.g0_0_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m27_1\ : std_logic;
signal \Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83\ : std_logic;
signal \Lab_UT.dictrl.N_61\ : std_logic;
signal \Lab_UT.dictrl.N_62_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_9_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.state_fast_1\ : std_logic;
signal \Lab_UT.dictrl.N_1110_1\ : std_logic;
signal \Lab_UT.dictrl.N_1459_1\ : std_logic;
signal \Lab_UT.dictrl.N_40_8\ : std_logic;
signal \Lab_UT.dictrl.N_40_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1102_2\ : std_logic;
signal \Lab_UT.dictrl.g2_1_2\ : std_logic;
signal \Lab_UT.dictrl.N_1462_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3\ : std_logic;
signal \Lab_UT.dictrl.N_11_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0\ : std_logic;
signal \Lab_UT.dictrl.N_8\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_20_0\ : std_logic;
signal \Lab_UT.dictrl.N_18_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_fast_3\ : std_logic;
signal \Lab_UT.dictrl.state_fast_2\ : std_logic;
signal \Lab_UT.dictrl.state_1_rep1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_3_2\ : std_logic;
signal \Lab_UT.dictrl.N_11_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_4_6\ : std_logic;
signal \Lab_UT.dictrl.N_22_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_4_7\ : std_logic;
signal \Lab_UT.dictrl.m53_d_1_3\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_40\ : std_logic;
signal \Lab_UT.dictrl.N_62\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_1Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNO_0Z0Z_2\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep1\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_RNINV3PZ0Z_2\ : std_logic;
signal \Lab_UT.min2_3\ : std_logic;
signal \uu2.bitmapZ0Z_203\ : std_logic;
signal \uu2.bitmapZ0Z_200\ : std_logic;
signal \INVuu2.bitmap_203C_net\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_65\ : std_logic;
signal \uu2.N_54\ : std_logic;
signal \uu2.N_53\ : std_logic;
signal \uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_\ : std_logic;
signal \INVuu2.w_addr_displaying_1C_net\ : std_logic;
signal \Lab_UT.min1_2\ : std_logic;
signal \Lab_UT.min1_1\ : std_logic;
signal \Lab_UT.min1_3\ : std_logic;
signal \Lab_UT.min1_0\ : std_logic;
signal \uu2.bitmapZ0Z_69\ : std_logic;
signal \uu2.bitmapZ0Z_197\ : std_logic;
signal \uu2.un4_w_user_data_rdyZ0Z_0\ : std_logic;
signal \INVuu2.bitmap_197C_net\ : std_logic;
signal \buart__rx_startbit\ : std_logic;
signal \buart__rx_N_27_0_i\ : std_logic;
signal \buart.Z_rx.bitcount_cry_1_THRU_CO\ : std_logic;
signal \buart__rx_bitcount_2\ : std_logic;
signal \buart.Z_rx.bitcounte_0_0\ : std_logic;
signal \uu2.bitmapZ0Z_75\ : std_logic;
signal \uu2.bitmapZ0Z_72\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_1\ : std_logic;
signal \uu2.vram_rd_clk_detZ0Z_0\ : std_logic;
signal \uu2.vram_rd_clk_det_RNI95711Z0Z_1\ : std_logic;
signal \Lab_UT.di_ASones_3\ : std_logic;
signal \Lab_UT.min2_1\ : std_logic;
signal \Lab_UT.min2_2\ : std_logic;
signal \Lab_UT.di_AStens_3\ : std_logic;
signal \Lab_UT.didp.regrce2.LdAStens_0\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.di_AMtens_2\ : std_logic;
signal \Lab_UT.di_AMtens_1\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_0\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_1\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.loadalarm_0_cascade_\ : std_logic;
signal \Lab_UT.min2_0\ : std_logic;
signal \Lab_UT.di_AMones_0\ : std_logic;
signal \Lab_UT.di_AMtens_0\ : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_1_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_18\ : std_logic;
signal \Lab_UT.dictrl.m35_0\ : std_logic;
signal \Lab_UT.didp.countrce4.un13_qPone\ : std_logic;
signal \Lab_UT.LdAMtens\ : std_logic;
signal \Lab_UT.LdAMones\ : std_logic;
signal \Lab_UT.LdAStens\ : std_logic;
signal \Lab_UT.dictrl.N_1460_2\ : std_logic;
signal \Lab_UT.dictrl.state_fast_0\ : std_logic;
signal \Lab_UT.dictrl.N_23_1\ : std_logic;
signal \G_17_i_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_latmux_2_1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_3\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.G_17_i_a5_1_1\ : std_logic;
signal \Lab_UT.dictrl.state_1_rep2\ : std_logic;
signal \Lab_UT.dictrl.N_15_0\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_2\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_0_2_cascade_\ : std_logic;
signal rst : std_logic;
signal \Lab_UT.dictrl.g0_12_a6_2_2\ : std_logic;
signal \Lab_UT.dictrl.N_19\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3\ : std_logic;
signal \Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1792_0_0_0\ : std_logic;
signal \Lab_UT.dictrl.m53_d_1_5\ : std_logic;
signal bu_rx_data_4_rep1 : std_logic;
signal \Lab_UT.dictrl.N_40_0\ : std_logic;
signal \Lab_UT.dictrl.N_6\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_i_1\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a5_0_2\ : std_logic;
signal \Lab_UT.dictrl.g2_2\ : std_logic;
signal \Lab_UT.dictrl.g2_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_3_1\ : std_logic;
signal \Lab_UT.dictrl.g1_1\ : std_logic;
signal \Lab_UT.dictrl.N_5\ : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_9\ : std_logic;
signal \Lab_UT.dictrl.g2_1_3\ : std_logic;
signal \Lab_UT.dictrl.N_1462_3_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1102_3\ : std_logic;
signal \Lab_UT.dictrl.N_1460_3\ : std_logic;
signal \Lab_UT.dictrl.m53_d_1_1\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_3_cascade_\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_42\ : std_logic;
signal \uu2.w_addr_userZ0Z_1\ : std_logic;
signal \uu2.w_addr_userZ0Z_2\ : std_logic;
signal \uu2.un3_w_addr_user_4_cascade_\ : std_logic;
signal \uu2.un3_w_addr_user_5\ : std_logic;
signal \uu2.un3_w_addr_user\ : std_logic;
signal \INVuu2.w_addr_displaying_nesr_5C_net\ : std_logic;
signal \uu2.un21_w_addr_displaying_0_0\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33\ : std_logic;
signal \uu2.w_addr_displayingZ1Z_4\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_33_cascade_\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_2\ : std_logic;
signal \uu2.bitmap_pmux_sn_m15_0_1\ : std_logic;
signal \uu2.w_addr_displaying_0_rep1_RNIDASJZ0\ : std_logic;
signal \uu2.w_addr_displaying_RNIR2PLZ0Z_8\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1\ : std_logic;
signal \uu2.bitmap_pmux_29_0\ : std_logic;
signal \uu2.N_24_0\ : std_logic;
signal \uu2.w_addr_displaying_RNIU1AF7Z0Z_0\ : std_logic;
signal \INVuu2.w_addr_displaying_3C_net\ : std_logic;
signal \Lab_UT.dictrl.m12Z0Z_2\ : std_logic;
signal \INVuu2.bitmap_215C_net\ : std_logic;
signal \uu2.bitmapZ0Z_215\ : std_logic;
signal \uu2.N_198_cascade_\ : std_logic;
signal \uu2.N_199\ : std_logic;
signal \uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_\ : std_logic;
signal \uu2.N_196\ : std_logic;
signal \uu2.bitmap_pmux_27_i_m2_ns_1\ : std_logic;
signal \INVuu2.bitmap_93C_net\ : std_logic;
signal \uu2.w_addr_displaying_0_repZ0Z1\ : std_logic;
signal \uu2.N_15\ : std_logic;
signal \uu2.N_17\ : std_logic;
signal \uu2.bitmap_pmux_25_i_m2_ns_1_cascade_\ : std_logic;
signal \uu2.N_49\ : std_logic;
signal \uu2.bitmapZ0Z_221\ : std_logic;
signal \uu2.bitmapZ0Z_93\ : std_logic;
signal \uu2.N_13\ : std_logic;
signal \Lab_UT.didp.countrce1.un20_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.di_Sones_3\ : std_logic;
signal \Lab_UT.didp.countrce1.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.di_Sones_2\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_12\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_4_cascade_\ : std_logic;
signal \Lab_UT.dispString.N_128_mux\ : std_logic;
signal \Lab_UT.di_AStens_2\ : std_logic;
signal \Lab_UT.di_ASones_2\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_1\ : std_logic;
signal \Lab_UT.LdASones\ : std_logic;
signal \Lab_UT.didp.regrce1.LdASones_0\ : std_logic;
signal \Lab_UT.di_ASones_0\ : std_logic;
signal \Lab_UT.dispString.N_180\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_7\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_11\ : std_logic;
signal \Lab_UT.didp.countrce1.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.di_Sones_0\ : std_logic;
signal \Lab_UT.LdMtens_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.LdMtens\ : std_logic;
signal \Lab_UT.didp.countrce4.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMtens_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_rep1\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0\ : std_logic;
signal \Lab_UT.state_i_4_0\ : std_logic;
signal \Lab_UT.dicRun_2\ : std_logic;
signal bu_rx_data_7 : std_logic;
signal bu_rx_data_6 : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_1_5\ : std_logic;
signal \Lab_UT.dictrl.g0_i_a4_1_4_cascade_\ : std_logic;
signal bu_rx_data_5 : std_logic;
signal \Lab_UT.dictrl.N_12\ : std_logic;
signal \Lab_UT.dictrl.N_4\ : std_logic;
signal bu_rx_data_4 : std_logic;
signal \Lab_UT.dictrl.N_7\ : std_logic;
signal bu_rx_data_3_rep2 : std_logic;
signal \Lab_UT.N_115\ : std_logic;
signal \Lab_UT.dictrl.N_39\ : std_logic;
signal bu_rx_data_6_rep1 : std_logic;
signal \Lab_UT.dictrl.m53_d_1_0\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1\ : std_logic;
signal \Lab_UT.dictrl.N_1462_0\ : std_logic;
signal \Lab_UT.dictrl.N_1102_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_7\ : std_logic;
signal \Lab_UT.dictrl.N_1106_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g1_1_1_0\ : std_logic;
signal bu_rx_data_7_rep1 : std_logic;
signal \Lab_UT.dictrl.N_59\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux\ : std_logic;
signal \Lab_UT.dictrl.N_59_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_0_rep2\ : std_logic;
signal \Lab_UT.dictrl.N_40_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_40_4\ : std_logic;
signal \Lab_UT.dictrl.N_40_2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.m23_aZ0Z0\ : std_logic;
signal \Lab_UT.dictrl.N_40_7\ : std_logic;
signal \Lab_UT.dictrl.N_40_7_cascade_\ : std_logic;
signal \Lab_UT.dictrl.g2_1_5\ : std_logic;
signal \Lab_UT.dictrl.N_1462_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1102_5\ : std_logic;
signal bu_rx_data_0_rep1 : std_logic;
signal bu_rx_data_5_rep1 : std_logic;
signal bu_rx_data_4_rep2 : std_logic;
signal \Lab_UT.dictrl.g0_i_m2_0_a7_4_8\ : std_logic;
signal \Lab_UT.dictrl.N_19_0\ : std_logic;
signal bu_rx_data_6_rep2 : std_logic;
signal \Lab_UT.dictrl.m40Z0Z_1\ : std_logic;
signal \Lab_UT.dictrl.m53_d_1_4\ : std_logic;
signal \Lab_UT.dictrl.state_2_rep2\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_6_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_3_rep2\ : std_logic;
signal \Lab_UT.dictrl.g2_1_4\ : std_logic;
signal \Lab_UT.dictrl.N_1462_4\ : std_logic;
signal \Lab_UT.dictrl.N_1102_4_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_6_0\ : std_logic;
signal \Lab_UT.dictrl.next_state_2_1\ : std_logic;
signal \Lab_UT.dictrl.g0_i_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_5\ : std_logic;
signal \uu2.w_addr_userZ0Z_4\ : std_logic;
signal \uu2.un28_w_addr_user_i\ : std_logic;
signal \uu2.un404_ci\ : std_logic;
signal \uu2.un426_ci_3\ : std_logic;
signal \uu2.w_addr_userZ0Z_6\ : std_logic;
signal \INVuu2.w_addr_user_5C_net\ : std_logic;
signal \uu2.w_addr_user_RNI43E87Z0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_\ : std_logic;
signal \uu2.N_397\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_1\ : std_logic;
signal \uu2.w_addr_displayingZ1Z_3\ : std_logic;
signal \uu2.bitmap_pmux_sn_N_11\ : std_logic;
signal \uu2.N_32\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_3\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_2\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2\ : std_logic;
signal \INVuu2.bitmap_314C_net\ : std_logic;
signal \uu2.bitmapZ0Z_218\ : std_logic;
signal \uu2.bitmapZ0Z_90\ : std_logic;
signal \uu2.N_20\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_7\ : std_logic;
signal \uu2.bitmap_RNIE7RKZ0Z_58_cascade_\ : std_logic;
signal \uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7\ : std_logic;
signal \uu2.bitmapZ0Z_314\ : std_logic;
signal \uu2.bitmap_RNI020QZ0Z_186\ : std_logic;
signal \uu2.bitmapZ0Z_186\ : std_logic;
signal \Lab_UT.sec2_1\ : std_logic;
signal \Lab_UT.sec2_3\ : std_logic;
signal \Lab_UT.sec2_2\ : std_logic;
signal \Lab_UT.sec2_0\ : std_logic;
signal \uu2.bitmapZ0Z_58\ : std_logic;
signal \INVuu2.bitmap_87C_net\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_0_cascade_\ : std_logic;
signal \Lab_UT.di_AStens_0\ : std_logic;
signal \Lab_UT.loadalarm_0\ : std_logic;
signal \Lab_UT.di_Sones_1\ : std_logic;
signal \Lab_UT.di_AStens_1\ : std_logic;
signal \Lab_UT.di_ASones_1\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_5\ : std_logic;
signal \Lab_UT.di_AMones_3\ : std_logic;
signal \Lab_UT.didp.regrce3.LdAMones_0\ : std_logic;
signal bu_rx_data_0 : std_logic;
signal \Lab_UT.didp.countrce3.q_5_0\ : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_1\ : std_logic;
signal \Lab_UT.di_AMones_2\ : std_logic;
signal \Lab_UT.di_AMones_1\ : std_logic;
signal \Lab_UT.dispString.m49Z0Z_2\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_2\ : std_logic;
signal \Lab_UT.didp.un24_ce_2\ : std_logic;
signal \Lab_UT.di_Mtens_1\ : std_logic;
signal \Lab_UT.didp.ce_12_3_cascade_\ : std_logic;
signal \Lab_UT.di_Mtens_3\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_3\ : std_logic;
signal \Lab_UT.didp.un18_ce\ : std_logic;
signal \oneSecStrb\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_0\ : std_logic;
signal \Lab_UT.di_Mtens_0\ : std_logic;
signal \Lab_UT.di_Mtens_2\ : std_logic;
signal \Lab_UT.didp.reset_12_1_3\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_1\ : std_logic;
signal \Lab_UT.LdStens_i_4\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.N_1460_4\ : std_logic;
signal \Lab_UT.dictrl.g2_4\ : std_logic;
signal \Lab_UT.dictrl.next_state_4_1_cascade_\ : std_logic;
signal \Lab_UT.didp.ceZ0Z_0\ : std_logic;
signal \Lab_UT.LdSones_i_4\ : std_logic;
signal \Lab_UT.didp.un1_dicLdSones_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_2\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_3\ : std_logic;
signal \Lab_UT.LdSones\ : std_logic;
signal bu_rx_data_rdy_0_g : std_logic;
signal \Lab_UT.dictrl.g2_5\ : std_logic;
signal \Lab_UT.dictrl.g1_3\ : std_logic;
signal \Lab_UT.dictrl.g2_5_cascade_\ : std_logic;
signal \Lab_UT.dictrl.N_1460_5\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12and_0_ns_sn\ : std_logic;
signal \Lab_UT.dictrl.state_ret_12and_0_ns_rn_0\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g2_0_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_2_0_1\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_1\ : std_logic;
signal \Lab_UT.dictrl.N_1460_0\ : std_logic;
signal \Lab_UT.dictrl.g2_cascade_\ : std_logic;
signal \Lab_UT.dictrl.next_state_0_1\ : std_logic;
signal \Lab_UT.dictrl.N_40_3\ : std_logic;
signal \Lab_UT.dictrl.N_1105_1_cascade_\ : std_logic;
signal \Lab_UT.dictrl.state_i_3_2\ : std_logic;
signal \Lab_UT.dictrl.N_79_0\ : std_logic;
signal \Lab_UT.dictrl.N_40_5\ : std_logic;
signal \Lab_UT.dictrl.g1_2\ : std_logic;
signal \Lab_UT.dictrl.N_40_2\ : std_logic;
signal \Lab_UT.dictrl.g1_0\ : std_logic;
signal \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0\ : std_logic;
signal \Lab_UT.state_3\ : std_logic;
signal \Lab_UT.dictrl.N_40_1\ : std_logic;
signal \Lab_UT.dictrl.g1\ : std_logic;
signal \Lab_UT.dictrl.N_97_mux_4\ : std_logic;
signal \Lab_UT.dictrl.stateZ0Z_0\ : std_logic;
signal \Lab_UT.dictrl.g1_1_1\ : std_logic;
signal \Lab_UT.dictrl.m34_4\ : std_logic;
signal \Lab_UT.dictrl.N_1106_0\ : std_logic;
signal \Lab_UT.dictrl.N_1462_1\ : std_logic;
signal \Lab_UT.dictrl.N_1102_1\ : std_logic;
signal \Lab_UT.dictrl.g2_1_1\ : std_logic;
signal \Lab_UT.dictrl.un1_next_state66_0\ : std_logic;
signal \Lab_UT.dictrl.N_1460_1\ : std_logic;
signal \L3_tx_data_rdy\ : std_logic;
signal \uu2.un1_w_user_cr_0\ : std_logic;
signal \uu2.w_addr_userZ0Z_8\ : std_logic;
signal \uu2.mem0.w_addr_8\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_1\ : std_logic;
signal \uu2.N_75_mux\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_0\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_5\ : std_logic;
signal \uu2.N_14_i_cascade_\ : std_logic;
signal \uu2.N_15_i\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_8\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_7\ : std_logic;
signal \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\ : std_logic;
signal \uu2.N_33_cascade_\ : std_logic;
signal \uu2.N_14_i\ : std_logic;
signal \uu2.w_addr_displayingZ0Z_6\ : std_logic;
signal \INVuu2.w_addr_displaying_0C_net\ : std_logic;
signal \uu2.bitmapZ0Z_212\ : std_logic;
signal \uu2.bitmapZ0Z_180\ : std_logic;
signal \INVuu2.bitmap_212C_net\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_8\ : std_logic;
signal \uu2.bitmapZ0Z_52\ : std_logic;
signal \uu2.bitmapZ0Z_308\ : std_logic;
signal \uu2.N_194\ : std_logic;
signal \uu2.bitmapZ0Z_87\ : std_logic;
signal \uu2.w_addr_displaying_fastZ0Z_0\ : std_logic;
signal \uu2.N_197\ : std_logic;
signal \Lab_UT.sec1_2\ : std_logic;
signal \Lab_UT.sec1_1\ : std_logic;
signal \Lab_UT.sec1_3\ : std_logic;
signal \Lab_UT.sec1_0\ : std_logic;
signal \uu2.bitmapZ0Z_84\ : std_logic;
signal \INVuu2.bitmap_84C_net\ : std_logic;
signal \Lab_UT.didp.countrce2.un13_qPone_cascade_\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.di_Stens_2\ : std_logic;
signal \Lab_UT.di_Stens_0\ : std_logic;
signal bu_rx_data_1 : std_logic;
signal \Lab_UT.didp.un1_dicLdStens_0\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_1_cascade_\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_1\ : std_logic;
signal \Lab_UT.di_Stens_1\ : std_logic;
signal \Lab_UT.didp.countrce2.un20_qPone\ : std_logic;
signal \Lab_UT.LdStens\ : std_logic;
signal \Lab_UT.di_Stens_3\ : std_logic;
signal \Lab_UT.didp.countrce2.q_5_3\ : std_logic;
signal \Lab_UT.didp.countrce3.ce_12_2_3\ : std_logic;
signal \Lab_UT.didp.countrce3.un13_qPone_cascade_\ : std_logic;
signal bu_rx_data_2 : std_logic;
signal \Lab_UT.didp.countrce3.q_5_2_cascade_\ : std_logic;
signal \Lab_UT.di_Mones_1\ : std_logic;
signal \Lab_UT.di_Mones_0\ : std_logic;
signal \Lab_UT.di_Mones_2\ : std_logic;
signal \Lab_UT.LdMones\ : std_logic;
signal \Lab_UT.didp.countrce3.un20_qPone_cascade_\ : std_logic;
signal bu_rx_data_3 : std_logic;
signal \Lab_UT.didp.un1_dicLdMones_0\ : std_logic;
signal \Lab_UT.didp.resetZ0Z_2\ : std_logic;
signal \Lab_UT.didp.countrce3.q_5_3_cascade_\ : std_logic;
signal \Lab_UT.di_Mones_3\ : std_logic;
signal clk_g : std_logic;
signal bu_rx_data_rdy : std_logic;
signal rst_g : std_logic;
signal bu_rx_data_rdy_0 : std_logic;
signal \_gnd_net_\ : std_logic;

signal led_wire : std_logic_vector(4 downto 0);
signal from_pc_wire : std_logic;
signal clk_in_wire : std_logic;
signal to_ir_wire : std_logic;
signal o_serial_data_wire : std_logic;
signal sd_wire : std_logic;
signal \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    led <= led_wire;
    from_pc_wire <= from_pc;
    clk_in_wire <= clk_in;
    to_ir <= to_ir_wire;
    o_serial_data <= o_serial_data_wire;
    sd <= sd_wire;
    \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    \uu2.r_data_wire_7\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(14);
    \uu2.r_data_wire_6\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(12);
    \uu2.r_data_wire_5\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(10);
    \uu2.r_data_wire_4\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(8);
    \uu2.r_data_wire_3\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(6);
    \uu2.r_data_wire_2\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(4);
    \uu2.r_data_wire_1\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(2);
    \uu2.r_data_wire_0\ <= \uu2.mem0.ram512X8_inst_physical_RDATA_wire\(0);
    \uu2.mem0.ram512X8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__11040\&\N__11025\&\N__11220\&\N__11937\&\N__12015\&\N__11199\&\N__11175\&\N__11148\&\N__11109\;
    \uu2.mem0.ram512X8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__23511\&\N__14397\&\N__14439\&\N__14451\&\N__13041\&\N__13059\&\N__11811\&\N__11823\&\N__11874\;
    \uu2.mem0.ram512X8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uu2.mem0.ram512X8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__13101\&'0'&\N__12942\&'0'&\N__12915\&'0'&\N__12951\&'0'&\N__13320\&'0'&\N__13137\&'0'&\N__13119\;

    \latticehx1k_pll_inst.latticehx1k_pll_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "110",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            SCLK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => clk,
            REFERENCECLK => \N__9504\,
            RESETB => \N__16951\,
            BYPASS => \GNDG0\,
            SDI => \GNDG0\,
            DYNAMICDELAY => \latticehx1k_pll_inst.latticehx1k_pll_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \uu2.mem0.ram512X8_inst_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_F => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_E => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_D => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_C => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_B => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_A => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_9 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_8 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_7 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_6 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_5 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_4 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_3 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_2 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000",
            INIT_1 => "0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000"
        )
    port map (
            RDATA => \uu2.mem0.ram512X8_inst_physical_RDATA_wire\,
            RADDR => \uu2.mem0.ram512X8_inst_physical_RADDR_wire\,
            WADDR => \uu2.mem0.ram512X8_inst_physical_WADDR_wire\,
            MASK => \uu2.mem0.ram512X8_inst_physical_MASK_wire\,
            WDATA => \uu2.mem0.ram512X8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__26198\,
            RE => \N__16944\,
            WCLKE => \N__11840\,
            WCLK => \N__26197\,
            WE => \N__11844\
        );

    \led_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26842\,
            DIN => \N__26841\,
            DOUT => \N__26840\,
            PACKAGEPIN => led_wire(3)
        );

    \led_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__26842\,
            PADOUT => \N__26841\,
            PADIN => \N__26840\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26833\,
            DIN => \N__26832\,
            DOUT => \N__26831\,
            PACKAGEPIN => led_wire(4)
        );

    \led_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__26833\,
            PADOUT => \N__26832\,
            PADIN => \N__26831\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \Z_rcxd.Z_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26824\,
            DIN => \N__26823\,
            DOUT => \N__26822\,
            PACKAGEPIN => from_pc_wire
        );

    \Z_rcxd.Z_io_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000000",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__26824\,
            PADOUT => \N__26823\,
            PADIN => \N__26822\,
            CLOCKENABLE => 'H',
            DOUT1 => \GNDG0\,
            OUTPUTENABLE => '0',
            DIN0 => \uart_RXD\,
            DOUT0 => \GNDG0\,
            INPUTCLK => \N__26142\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_in_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26815\,
            DIN => \N__26814\,
            DOUT => \N__26813\,
            PACKAGEPIN => clk_in_wire
        );

    \clk_in_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__26815\,
            PADOUT => \N__26814\,
            PADIN => \N__26813\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_in_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26806\,
            DIN => \N__26805\,
            DOUT => \N__26804\,
            PACKAGEPIN => led_wire(1)
        );

    \led_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__26806\,
            PADOUT => \N__26805\,
            PADIN => \N__26804\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26797\,
            DIN => \N__26796\,
            DOUT => \N__26795\,
            PACKAGEPIN => led_wire(2)
        );

    \led_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__26797\,
            PADOUT => \N__26796\,
            PADIN => \N__26795\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \to_ir_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26788\,
            DIN => \N__26787\,
            DOUT => \N__26786\,
            PACKAGEPIN => to_ir_wire
        );

    \to_ir_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26788\,
            PADOUT => \N__26787\,
            PADIN => \N__26786\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_serial_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26779\,
            DIN => \N__26778\,
            DOUT => \N__26777\,
            PACKAGEPIN => o_serial_data_wire
        );

    \o_serial_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26779\,
            PADOUT => \N__26778\,
            PADIN => \N__26777\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sd_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26770\,
            DIN => \N__26769\,
            DOUT => \N__26768\,
            PACKAGEPIN => sd_wire
        );

    \sd_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__26770\,
            PADOUT => \N__26769\,
            PADIN => \N__26768\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__26761\,
            DIN => \N__26760\,
            DOUT => \N__26759\,
            PACKAGEPIN => led_wire(0)
        );

    \led_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__26761\,
            PADOUT => \N__26760\,
            PADIN => \N__26759\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6553\ : CascadeMux
    port map (
            O => \N__26742\,
            I => \Lab_UT.didp.countrce3.un13_qPone_cascade_\
        );

    \I__6552\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26735\
        );

    \I__6551\ : InMux
    port map (
            O => \N__26738\,
            I => \N__26732\
        );

    \I__6550\ : LocalMux
    port map (
            O => \N__26735\,
            I => \N__26725\
        );

    \I__6549\ : LocalMux
    port map (
            O => \N__26732\,
            I => \N__26725\
        );

    \I__6548\ : InMux
    port map (
            O => \N__26731\,
            I => \N__26719\
        );

    \I__6547\ : InMux
    port map (
            O => \N__26730\,
            I => \N__26716\
        );

    \I__6546\ : Span4Mux_v
    port map (
            O => \N__26725\,
            I => \N__26712\
        );

    \I__6545\ : InMux
    port map (
            O => \N__26724\,
            I => \N__26709\
        );

    \I__6544\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26706\
        );

    \I__6543\ : InMux
    port map (
            O => \N__26722\,
            I => \N__26703\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__26719\,
            I => \N__26700\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__26716\,
            I => \N__26697\
        );

    \I__6540\ : InMux
    port map (
            O => \N__26715\,
            I => \N__26694\
        );

    \I__6539\ : IoSpan4Mux
    port map (
            O => \N__26712\,
            I => \N__26690\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__26709\,
            I => \N__26681\
        );

    \I__6537\ : LocalMux
    port map (
            O => \N__26706\,
            I => \N__26681\
        );

    \I__6536\ : LocalMux
    port map (
            O => \N__26703\,
            I => \N__26672\
        );

    \I__6535\ : Span4Mux_s2_h
    port map (
            O => \N__26700\,
            I => \N__26672\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__26697\,
            I => \N__26672\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__26694\,
            I => \N__26672\
        );

    \I__6532\ : InMux
    port map (
            O => \N__26693\,
            I => \N__26669\
        );

    \I__6531\ : IoSpan4Mux
    port map (
            O => \N__26690\,
            I => \N__26664\
        );

    \I__6530\ : InMux
    port map (
            O => \N__26689\,
            I => \N__26655\
        );

    \I__6529\ : InMux
    port map (
            O => \N__26688\,
            I => \N__26655\
        );

    \I__6528\ : InMux
    port map (
            O => \N__26687\,
            I => \N__26655\
        );

    \I__6527\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26655\
        );

    \I__6526\ : Span4Mux_v
    port map (
            O => \N__26681\,
            I => \N__26652\
        );

    \I__6525\ : Span4Mux_h
    port map (
            O => \N__26672\,
            I => \N__26644\
        );

    \I__6524\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26644\
        );

    \I__6523\ : InMux
    port map (
            O => \N__26668\,
            I => \N__26639\
        );

    \I__6522\ : InMux
    port map (
            O => \N__26667\,
            I => \N__26639\
        );

    \I__6521\ : Span4Mux_s2_h
    port map (
            O => \N__26664\,
            I => \N__26634\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__26655\,
            I => \N__26634\
        );

    \I__6519\ : Sp12to4
    port map (
            O => \N__26652\,
            I => \N__26631\
        );

    \I__6518\ : InMux
    port map (
            O => \N__26651\,
            I => \N__26628\
        );

    \I__6517\ : InMux
    port map (
            O => \N__26650\,
            I => \N__26623\
        );

    \I__6516\ : InMux
    port map (
            O => \N__26649\,
            I => \N__26623\
        );

    \I__6515\ : Span4Mux_v
    port map (
            O => \N__26644\,
            I => \N__26618\
        );

    \I__6514\ : LocalMux
    port map (
            O => \N__26639\,
            I => \N__26618\
        );

    \I__6513\ : Span4Mux_h
    port map (
            O => \N__26634\,
            I => \N__26612\
        );

    \I__6512\ : Span12Mux_s10_h
    port map (
            O => \N__26631\,
            I => \N__26607\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__26628\,
            I => \N__26607\
        );

    \I__6510\ : LocalMux
    port map (
            O => \N__26623\,
            I => \N__26604\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__26618\,
            I => \N__26601\
        );

    \I__6508\ : InMux
    port map (
            O => \N__26617\,
            I => \N__26594\
        );

    \I__6507\ : InMux
    port map (
            O => \N__26616\,
            I => \N__26594\
        );

    \I__6506\ : InMux
    port map (
            O => \N__26615\,
            I => \N__26594\
        );

    \I__6505\ : Span4Mux_h
    port map (
            O => \N__26612\,
            I => \N__26591\
        );

    \I__6504\ : Odrv12
    port map (
            O => \N__26607\,
            I => bu_rx_data_2
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__26604\,
            I => bu_rx_data_2
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__26601\,
            I => bu_rx_data_2
        );

    \I__6501\ : LocalMux
    port map (
            O => \N__26594\,
            I => bu_rx_data_2
        );

    \I__6500\ : Odrv4
    port map (
            O => \N__26591\,
            I => bu_rx_data_2
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__26580\,
            I => \Lab_UT.didp.countrce3.q_5_2_cascade_\
        );

    \I__6498\ : InMux
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__26574\,
            I => \N__26567\
        );

    \I__6496\ : CascadeMux
    port map (
            O => \N__26573\,
            I => \N__26563\
        );

    \I__6495\ : InMux
    port map (
            O => \N__26572\,
            I => \N__26555\
        );

    \I__6494\ : InMux
    port map (
            O => \N__26571\,
            I => \N__26555\
        );

    \I__6493\ : InMux
    port map (
            O => \N__26570\,
            I => \N__26555\
        );

    \I__6492\ : Span4Mux_v
    port map (
            O => \N__26567\,
            I => \N__26552\
        );

    \I__6491\ : InMux
    port map (
            O => \N__26566\,
            I => \N__26545\
        );

    \I__6490\ : InMux
    port map (
            O => \N__26563\,
            I => \N__26545\
        );

    \I__6489\ : InMux
    port map (
            O => \N__26562\,
            I => \N__26545\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__26555\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__6487\ : Odrv4
    port map (
            O => \N__26552\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__26545\,
            I => \Lab_UT.di_Mones_1\
        );

    \I__6485\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26532\
        );

    \I__6484\ : InMux
    port map (
            O => \N__26537\,
            I => \N__26532\
        );

    \I__6483\ : LocalMux
    port map (
            O => \N__26532\,
            I => \N__26524\
        );

    \I__6482\ : InMux
    port map (
            O => \N__26531\,
            I => \N__26521\
        );

    \I__6481\ : InMux
    port map (
            O => \N__26530\,
            I => \N__26518\
        );

    \I__6480\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26511\
        );

    \I__6479\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26511\
        );

    \I__6478\ : InMux
    port map (
            O => \N__26527\,
            I => \N__26511\
        );

    \I__6477\ : Span4Mux_h
    port map (
            O => \N__26524\,
            I => \N__26508\
        );

    \I__6476\ : LocalMux
    port map (
            O => \N__26521\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__26518\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__6474\ : LocalMux
    port map (
            O => \N__26511\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__6473\ : Odrv4
    port map (
            O => \N__26508\,
            I => \Lab_UT.di_Mones_0\
        );

    \I__6472\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26494\
        );

    \I__6471\ : CascadeMux
    port map (
            O => \N__26498\,
            I => \N__26489\
        );

    \I__6470\ : CascadeMux
    port map (
            O => \N__26497\,
            I => \N__26486\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26483\
        );

    \I__6468\ : InMux
    port map (
            O => \N__26493\,
            I => \N__26473\
        );

    \I__6467\ : InMux
    port map (
            O => \N__26492\,
            I => \N__26473\
        );

    \I__6466\ : InMux
    port map (
            O => \N__26489\,
            I => \N__26473\
        );

    \I__6465\ : InMux
    port map (
            O => \N__26486\,
            I => \N__26473\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__26483\,
            I => \N__26470\
        );

    \I__6463\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26467\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__26473\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__6461\ : Odrv4
    port map (
            O => \N__26470\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__26467\,
            I => \Lab_UT.di_Mones_2\
        );

    \I__6459\ : InMux
    port map (
            O => \N__26460\,
            I => \N__26452\
        );

    \I__6458\ : InMux
    port map (
            O => \N__26459\,
            I => \N__26449\
        );

    \I__6457\ : InMux
    port map (
            O => \N__26458\,
            I => \N__26440\
        );

    \I__6456\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26440\
        );

    \I__6455\ : InMux
    port map (
            O => \N__26456\,
            I => \N__26440\
        );

    \I__6454\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26440\
        );

    \I__6453\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26435\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__26449\,
            I => \N__26435\
        );

    \I__6451\ : LocalMux
    port map (
            O => \N__26440\,
            I => \N__26432\
        );

    \I__6450\ : Odrv4
    port map (
            O => \N__26435\,
            I => \Lab_UT.LdMones\
        );

    \I__6449\ : Odrv4
    port map (
            O => \N__26432\,
            I => \Lab_UT.LdMones\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__26427\,
            I => \Lab_UT.didp.countrce3.un20_qPone_cascade_\
        );

    \I__6447\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26417\
        );

    \I__6446\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26414\
        );

    \I__6445\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26409\
        );

    \I__6444\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26406\
        );

    \I__6443\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26403\
        );

    \I__6442\ : LocalMux
    port map (
            O => \N__26417\,
            I => \N__26398\
        );

    \I__6441\ : LocalMux
    port map (
            O => \N__26414\,
            I => \N__26398\
        );

    \I__6440\ : InMux
    port map (
            O => \N__26413\,
            I => \N__26395\
        );

    \I__6439\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26392\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26381\
        );

    \I__6437\ : LocalMux
    port map (
            O => \N__26406\,
            I => \N__26381\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26381\
        );

    \I__6435\ : Span4Mux_v
    port map (
            O => \N__26398\,
            I => \N__26378\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__26395\,
            I => \N__26373\
        );

    \I__6433\ : LocalMux
    port map (
            O => \N__26392\,
            I => \N__26373\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__26391\,
            I => \N__26367\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__26390\,
            I => \N__26364\
        );

    \I__6430\ : InMux
    port map (
            O => \N__26389\,
            I => \N__26361\
        );

    \I__6429\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26355\
        );

    \I__6428\ : Span4Mux_v
    port map (
            O => \N__26381\,
            I => \N__26350\
        );

    \I__6427\ : Span4Mux_h
    port map (
            O => \N__26378\,
            I => \N__26350\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__26373\,
            I => \N__26345\
        );

    \I__6425\ : InMux
    port map (
            O => \N__26372\,
            I => \N__26342\
        );

    \I__6424\ : InMux
    port map (
            O => \N__26371\,
            I => \N__26339\
        );

    \I__6423\ : InMux
    port map (
            O => \N__26370\,
            I => \N__26332\
        );

    \I__6422\ : InMux
    port map (
            O => \N__26367\,
            I => \N__26332\
        );

    \I__6421\ : InMux
    port map (
            O => \N__26364\,
            I => \N__26332\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__26361\,
            I => \N__26327\
        );

    \I__6419\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26320\
        );

    \I__6418\ : InMux
    port map (
            O => \N__26359\,
            I => \N__26320\
        );

    \I__6417\ : InMux
    port map (
            O => \N__26358\,
            I => \N__26320\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__26355\,
            I => \N__26317\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__26350\,
            I => \N__26314\
        );

    \I__6414\ : InMux
    port map (
            O => \N__26349\,
            I => \N__26309\
        );

    \I__6413\ : InMux
    port map (
            O => \N__26348\,
            I => \N__26309\
        );

    \I__6412\ : Span4Mux_h
    port map (
            O => \N__26345\,
            I => \N__26302\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__26342\,
            I => \N__26302\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__26339\,
            I => \N__26302\
        );

    \I__6409\ : LocalMux
    port map (
            O => \N__26332\,
            I => \N__26299\
        );

    \I__6408\ : InMux
    port map (
            O => \N__26331\,
            I => \N__26294\
        );

    \I__6407\ : InMux
    port map (
            O => \N__26330\,
            I => \N__26294\
        );

    \I__6406\ : Span4Mux_v
    port map (
            O => \N__26327\,
            I => \N__26289\
        );

    \I__6405\ : LocalMux
    port map (
            O => \N__26320\,
            I => \N__26289\
        );

    \I__6404\ : Span12Mux_s8_h
    port map (
            O => \N__26317\,
            I => \N__26282\
        );

    \I__6403\ : Sp12to4
    port map (
            O => \N__26314\,
            I => \N__26282\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__26309\,
            I => \N__26282\
        );

    \I__6401\ : Span4Mux_v
    port map (
            O => \N__26302\,
            I => \N__26277\
        );

    \I__6400\ : Span4Mux_h
    port map (
            O => \N__26299\,
            I => \N__26277\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__26294\,
            I => bu_rx_data_3
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__26289\,
            I => bu_rx_data_3
        );

    \I__6397\ : Odrv12
    port map (
            O => \N__26282\,
            I => bu_rx_data_3
        );

    \I__6396\ : Odrv4
    port map (
            O => \N__26277\,
            I => bu_rx_data_3
        );

    \I__6395\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26262\
        );

    \I__6394\ : InMux
    port map (
            O => \N__26267\,
            I => \N__26262\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__26262\,
            I => \Lab_UT.didp.un1_dicLdMones_0\
        );

    \I__6392\ : CascadeMux
    port map (
            O => \N__26259\,
            I => \N__26253\
        );

    \I__6391\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26248\
        );

    \I__6390\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26248\
        );

    \I__6389\ : InMux
    port map (
            O => \N__26256\,
            I => \N__26243\
        );

    \I__6388\ : InMux
    port map (
            O => \N__26253\,
            I => \N__26243\
        );

    \I__6387\ : LocalMux
    port map (
            O => \N__26248\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__6386\ : LocalMux
    port map (
            O => \N__26243\,
            I => \Lab_UT.didp.resetZ0Z_2\
        );

    \I__6385\ : CascadeMux
    port map (
            O => \N__26238\,
            I => \Lab_UT.didp.countrce3.q_5_3_cascade_\
        );

    \I__6384\ : CascadeMux
    port map (
            O => \N__26235\,
            I => \N__26232\
        );

    \I__6383\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26223\
        );

    \I__6382\ : InMux
    port map (
            O => \N__26231\,
            I => \N__26223\
        );

    \I__6381\ : InMux
    port map (
            O => \N__26230\,
            I => \N__26216\
        );

    \I__6380\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26216\
        );

    \I__6379\ : InMux
    port map (
            O => \N__26228\,
            I => \N__26216\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__26223\,
            I => \N__26213\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__26216\,
            I => \N__26208\
        );

    \I__6376\ : Span4Mux_h
    port map (
            O => \N__26213\,
            I => \N__26208\
        );

    \I__6375\ : Odrv4
    port map (
            O => \N__26208\,
            I => \Lab_UT.di_Mones_3\
        );

    \I__6374\ : ClkMux
    port map (
            O => \N__26205\,
            I => \N__25932\
        );

    \I__6373\ : ClkMux
    port map (
            O => \N__26204\,
            I => \N__25932\
        );

    \I__6372\ : ClkMux
    port map (
            O => \N__26203\,
            I => \N__25932\
        );

    \I__6371\ : ClkMux
    port map (
            O => \N__26202\,
            I => \N__25932\
        );

    \I__6370\ : ClkMux
    port map (
            O => \N__26201\,
            I => \N__25932\
        );

    \I__6369\ : ClkMux
    port map (
            O => \N__26200\,
            I => \N__25932\
        );

    \I__6368\ : ClkMux
    port map (
            O => \N__26199\,
            I => \N__25932\
        );

    \I__6367\ : ClkMux
    port map (
            O => \N__26198\,
            I => \N__25932\
        );

    \I__6366\ : ClkMux
    port map (
            O => \N__26197\,
            I => \N__25932\
        );

    \I__6365\ : ClkMux
    port map (
            O => \N__26196\,
            I => \N__25932\
        );

    \I__6364\ : ClkMux
    port map (
            O => \N__26195\,
            I => \N__25932\
        );

    \I__6363\ : ClkMux
    port map (
            O => \N__26194\,
            I => \N__25932\
        );

    \I__6362\ : ClkMux
    port map (
            O => \N__26193\,
            I => \N__25932\
        );

    \I__6361\ : ClkMux
    port map (
            O => \N__26192\,
            I => \N__25932\
        );

    \I__6360\ : ClkMux
    port map (
            O => \N__26191\,
            I => \N__25932\
        );

    \I__6359\ : ClkMux
    port map (
            O => \N__26190\,
            I => \N__25932\
        );

    \I__6358\ : ClkMux
    port map (
            O => \N__26189\,
            I => \N__25932\
        );

    \I__6357\ : ClkMux
    port map (
            O => \N__26188\,
            I => \N__25932\
        );

    \I__6356\ : ClkMux
    port map (
            O => \N__26187\,
            I => \N__25932\
        );

    \I__6355\ : ClkMux
    port map (
            O => \N__26186\,
            I => \N__25932\
        );

    \I__6354\ : ClkMux
    port map (
            O => \N__26185\,
            I => \N__25932\
        );

    \I__6353\ : ClkMux
    port map (
            O => \N__26184\,
            I => \N__25932\
        );

    \I__6352\ : ClkMux
    port map (
            O => \N__26183\,
            I => \N__25932\
        );

    \I__6351\ : ClkMux
    port map (
            O => \N__26182\,
            I => \N__25932\
        );

    \I__6350\ : ClkMux
    port map (
            O => \N__26181\,
            I => \N__25932\
        );

    \I__6349\ : ClkMux
    port map (
            O => \N__26180\,
            I => \N__25932\
        );

    \I__6348\ : ClkMux
    port map (
            O => \N__26179\,
            I => \N__25932\
        );

    \I__6347\ : ClkMux
    port map (
            O => \N__26178\,
            I => \N__25932\
        );

    \I__6346\ : ClkMux
    port map (
            O => \N__26177\,
            I => \N__25932\
        );

    \I__6345\ : ClkMux
    port map (
            O => \N__26176\,
            I => \N__25932\
        );

    \I__6344\ : ClkMux
    port map (
            O => \N__26175\,
            I => \N__25932\
        );

    \I__6343\ : ClkMux
    port map (
            O => \N__26174\,
            I => \N__25932\
        );

    \I__6342\ : ClkMux
    port map (
            O => \N__26173\,
            I => \N__25932\
        );

    \I__6341\ : ClkMux
    port map (
            O => \N__26172\,
            I => \N__25932\
        );

    \I__6340\ : ClkMux
    port map (
            O => \N__26171\,
            I => \N__25932\
        );

    \I__6339\ : ClkMux
    port map (
            O => \N__26170\,
            I => \N__25932\
        );

    \I__6338\ : ClkMux
    port map (
            O => \N__26169\,
            I => \N__25932\
        );

    \I__6337\ : ClkMux
    port map (
            O => \N__26168\,
            I => \N__25932\
        );

    \I__6336\ : ClkMux
    port map (
            O => \N__26167\,
            I => \N__25932\
        );

    \I__6335\ : ClkMux
    port map (
            O => \N__26166\,
            I => \N__25932\
        );

    \I__6334\ : ClkMux
    port map (
            O => \N__26165\,
            I => \N__25932\
        );

    \I__6333\ : ClkMux
    port map (
            O => \N__26164\,
            I => \N__25932\
        );

    \I__6332\ : ClkMux
    port map (
            O => \N__26163\,
            I => \N__25932\
        );

    \I__6331\ : ClkMux
    port map (
            O => \N__26162\,
            I => \N__25932\
        );

    \I__6330\ : ClkMux
    port map (
            O => \N__26161\,
            I => \N__25932\
        );

    \I__6329\ : ClkMux
    port map (
            O => \N__26160\,
            I => \N__25932\
        );

    \I__6328\ : ClkMux
    port map (
            O => \N__26159\,
            I => \N__25932\
        );

    \I__6327\ : ClkMux
    port map (
            O => \N__26158\,
            I => \N__25932\
        );

    \I__6326\ : ClkMux
    port map (
            O => \N__26157\,
            I => \N__25932\
        );

    \I__6325\ : ClkMux
    port map (
            O => \N__26156\,
            I => \N__25932\
        );

    \I__6324\ : ClkMux
    port map (
            O => \N__26155\,
            I => \N__25932\
        );

    \I__6323\ : ClkMux
    port map (
            O => \N__26154\,
            I => \N__25932\
        );

    \I__6322\ : ClkMux
    port map (
            O => \N__26153\,
            I => \N__25932\
        );

    \I__6321\ : ClkMux
    port map (
            O => \N__26152\,
            I => \N__25932\
        );

    \I__6320\ : ClkMux
    port map (
            O => \N__26151\,
            I => \N__25932\
        );

    \I__6319\ : ClkMux
    port map (
            O => \N__26150\,
            I => \N__25932\
        );

    \I__6318\ : ClkMux
    port map (
            O => \N__26149\,
            I => \N__25932\
        );

    \I__6317\ : ClkMux
    port map (
            O => \N__26148\,
            I => \N__25932\
        );

    \I__6316\ : ClkMux
    port map (
            O => \N__26147\,
            I => \N__25932\
        );

    \I__6315\ : ClkMux
    port map (
            O => \N__26146\,
            I => \N__25932\
        );

    \I__6314\ : ClkMux
    port map (
            O => \N__26145\,
            I => \N__25932\
        );

    \I__6313\ : ClkMux
    port map (
            O => \N__26144\,
            I => \N__25932\
        );

    \I__6312\ : ClkMux
    port map (
            O => \N__26143\,
            I => \N__25932\
        );

    \I__6311\ : ClkMux
    port map (
            O => \N__26142\,
            I => \N__25932\
        );

    \I__6310\ : ClkMux
    port map (
            O => \N__26141\,
            I => \N__25932\
        );

    \I__6309\ : ClkMux
    port map (
            O => \N__26140\,
            I => \N__25932\
        );

    \I__6308\ : ClkMux
    port map (
            O => \N__26139\,
            I => \N__25932\
        );

    \I__6307\ : ClkMux
    port map (
            O => \N__26138\,
            I => \N__25932\
        );

    \I__6306\ : ClkMux
    port map (
            O => \N__26137\,
            I => \N__25932\
        );

    \I__6305\ : ClkMux
    port map (
            O => \N__26136\,
            I => \N__25932\
        );

    \I__6304\ : ClkMux
    port map (
            O => \N__26135\,
            I => \N__25932\
        );

    \I__6303\ : ClkMux
    port map (
            O => \N__26134\,
            I => \N__25932\
        );

    \I__6302\ : ClkMux
    port map (
            O => \N__26133\,
            I => \N__25932\
        );

    \I__6301\ : ClkMux
    port map (
            O => \N__26132\,
            I => \N__25932\
        );

    \I__6300\ : ClkMux
    port map (
            O => \N__26131\,
            I => \N__25932\
        );

    \I__6299\ : ClkMux
    port map (
            O => \N__26130\,
            I => \N__25932\
        );

    \I__6298\ : ClkMux
    port map (
            O => \N__26129\,
            I => \N__25932\
        );

    \I__6297\ : ClkMux
    port map (
            O => \N__26128\,
            I => \N__25932\
        );

    \I__6296\ : ClkMux
    port map (
            O => \N__26127\,
            I => \N__25932\
        );

    \I__6295\ : ClkMux
    port map (
            O => \N__26126\,
            I => \N__25932\
        );

    \I__6294\ : ClkMux
    port map (
            O => \N__26125\,
            I => \N__25932\
        );

    \I__6293\ : ClkMux
    port map (
            O => \N__26124\,
            I => \N__25932\
        );

    \I__6292\ : ClkMux
    port map (
            O => \N__26123\,
            I => \N__25932\
        );

    \I__6291\ : ClkMux
    port map (
            O => \N__26122\,
            I => \N__25932\
        );

    \I__6290\ : ClkMux
    port map (
            O => \N__26121\,
            I => \N__25932\
        );

    \I__6289\ : ClkMux
    port map (
            O => \N__26120\,
            I => \N__25932\
        );

    \I__6288\ : ClkMux
    port map (
            O => \N__26119\,
            I => \N__25932\
        );

    \I__6287\ : ClkMux
    port map (
            O => \N__26118\,
            I => \N__25932\
        );

    \I__6286\ : ClkMux
    port map (
            O => \N__26117\,
            I => \N__25932\
        );

    \I__6285\ : ClkMux
    port map (
            O => \N__26116\,
            I => \N__25932\
        );

    \I__6284\ : ClkMux
    port map (
            O => \N__26115\,
            I => \N__25932\
        );

    \I__6283\ : GlobalMux
    port map (
            O => \N__25932\,
            I => \N__25929\
        );

    \I__6282\ : gio2CtrlBuf
    port map (
            O => \N__25929\,
            I => clk_g
        );

    \I__6281\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25919\
        );

    \I__6280\ : InMux
    port map (
            O => \N__25925\,
            I => \N__25919\
        );

    \I__6279\ : InMux
    port map (
            O => \N__25924\,
            I => \N__25915\
        );

    \I__6278\ : LocalMux
    port map (
            O => \N__25919\,
            I => \N__25912\
        );

    \I__6277\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25909\
        );

    \I__6276\ : LocalMux
    port map (
            O => \N__25915\,
            I => \N__25906\
        );

    \I__6275\ : Span4Mux_v
    port map (
            O => \N__25912\,
            I => \N__25903\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__25909\,
            I => \N__25900\
        );

    \I__6273\ : Span4Mux_s3_h
    port map (
            O => \N__25906\,
            I => \N__25896\
        );

    \I__6272\ : Sp12to4
    port map (
            O => \N__25903\,
            I => \N__25891\
        );

    \I__6271\ : Span12Mux_s1_h
    port map (
            O => \N__25900\,
            I => \N__25891\
        );

    \I__6270\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25888\
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__25896\,
            I => bu_rx_data_rdy
        );

    \I__6268\ : Odrv12
    port map (
            O => \N__25891\,
            I => bu_rx_data_rdy
        );

    \I__6267\ : LocalMux
    port map (
            O => \N__25888\,
            I => bu_rx_data_rdy
        );

    \I__6266\ : InMux
    port map (
            O => \N__25881\,
            I => \N__25869\
        );

    \I__6265\ : InMux
    port map (
            O => \N__25880\,
            I => \N__25866\
        );

    \I__6264\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25863\
        );

    \I__6263\ : InMux
    port map (
            O => \N__25878\,
            I => \N__25860\
        );

    \I__6262\ : InMux
    port map (
            O => \N__25877\,
            I => \N__25855\
        );

    \I__6261\ : InMux
    port map (
            O => \N__25876\,
            I => \N__25855\
        );

    \I__6260\ : InMux
    port map (
            O => \N__25875\,
            I => \N__25852\
        );

    \I__6259\ : InMux
    port map (
            O => \N__25874\,
            I => \N__25849\
        );

    \I__6258\ : InMux
    port map (
            O => \N__25873\,
            I => \N__25846\
        );

    \I__6257\ : InMux
    port map (
            O => \N__25872\,
            I => \N__25843\
        );

    \I__6256\ : LocalMux
    port map (
            O => \N__25869\,
            I => \N__25796\
        );

    \I__6255\ : LocalMux
    port map (
            O => \N__25866\,
            I => \N__25793\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__25863\,
            I => \N__25790\
        );

    \I__6253\ : LocalMux
    port map (
            O => \N__25860\,
            I => \N__25787\
        );

    \I__6252\ : LocalMux
    port map (
            O => \N__25855\,
            I => \N__25784\
        );

    \I__6251\ : LocalMux
    port map (
            O => \N__25852\,
            I => \N__25781\
        );

    \I__6250\ : LocalMux
    port map (
            O => \N__25849\,
            I => \N__25762\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__25846\,
            I => \N__25759\
        );

    \I__6248\ : LocalMux
    port map (
            O => \N__25843\,
            I => \N__25756\
        );

    \I__6247\ : SRMux
    port map (
            O => \N__25842\,
            I => \N__25617\
        );

    \I__6246\ : SRMux
    port map (
            O => \N__25841\,
            I => \N__25617\
        );

    \I__6245\ : SRMux
    port map (
            O => \N__25840\,
            I => \N__25617\
        );

    \I__6244\ : SRMux
    port map (
            O => \N__25839\,
            I => \N__25617\
        );

    \I__6243\ : SRMux
    port map (
            O => \N__25838\,
            I => \N__25617\
        );

    \I__6242\ : SRMux
    port map (
            O => \N__25837\,
            I => \N__25617\
        );

    \I__6241\ : SRMux
    port map (
            O => \N__25836\,
            I => \N__25617\
        );

    \I__6240\ : SRMux
    port map (
            O => \N__25835\,
            I => \N__25617\
        );

    \I__6239\ : SRMux
    port map (
            O => \N__25834\,
            I => \N__25617\
        );

    \I__6238\ : SRMux
    port map (
            O => \N__25833\,
            I => \N__25617\
        );

    \I__6237\ : SRMux
    port map (
            O => \N__25832\,
            I => \N__25617\
        );

    \I__6236\ : SRMux
    port map (
            O => \N__25831\,
            I => \N__25617\
        );

    \I__6235\ : SRMux
    port map (
            O => \N__25830\,
            I => \N__25617\
        );

    \I__6234\ : SRMux
    port map (
            O => \N__25829\,
            I => \N__25617\
        );

    \I__6233\ : SRMux
    port map (
            O => \N__25828\,
            I => \N__25617\
        );

    \I__6232\ : SRMux
    port map (
            O => \N__25827\,
            I => \N__25617\
        );

    \I__6231\ : SRMux
    port map (
            O => \N__25826\,
            I => \N__25617\
        );

    \I__6230\ : SRMux
    port map (
            O => \N__25825\,
            I => \N__25617\
        );

    \I__6229\ : SRMux
    port map (
            O => \N__25824\,
            I => \N__25617\
        );

    \I__6228\ : SRMux
    port map (
            O => \N__25823\,
            I => \N__25617\
        );

    \I__6227\ : SRMux
    port map (
            O => \N__25822\,
            I => \N__25617\
        );

    \I__6226\ : SRMux
    port map (
            O => \N__25821\,
            I => \N__25617\
        );

    \I__6225\ : SRMux
    port map (
            O => \N__25820\,
            I => \N__25617\
        );

    \I__6224\ : SRMux
    port map (
            O => \N__25819\,
            I => \N__25617\
        );

    \I__6223\ : SRMux
    port map (
            O => \N__25818\,
            I => \N__25617\
        );

    \I__6222\ : SRMux
    port map (
            O => \N__25817\,
            I => \N__25617\
        );

    \I__6221\ : SRMux
    port map (
            O => \N__25816\,
            I => \N__25617\
        );

    \I__6220\ : SRMux
    port map (
            O => \N__25815\,
            I => \N__25617\
        );

    \I__6219\ : SRMux
    port map (
            O => \N__25814\,
            I => \N__25617\
        );

    \I__6218\ : SRMux
    port map (
            O => \N__25813\,
            I => \N__25617\
        );

    \I__6217\ : SRMux
    port map (
            O => \N__25812\,
            I => \N__25617\
        );

    \I__6216\ : SRMux
    port map (
            O => \N__25811\,
            I => \N__25617\
        );

    \I__6215\ : SRMux
    port map (
            O => \N__25810\,
            I => \N__25617\
        );

    \I__6214\ : SRMux
    port map (
            O => \N__25809\,
            I => \N__25617\
        );

    \I__6213\ : SRMux
    port map (
            O => \N__25808\,
            I => \N__25617\
        );

    \I__6212\ : SRMux
    port map (
            O => \N__25807\,
            I => \N__25617\
        );

    \I__6211\ : SRMux
    port map (
            O => \N__25806\,
            I => \N__25617\
        );

    \I__6210\ : SRMux
    port map (
            O => \N__25805\,
            I => \N__25617\
        );

    \I__6209\ : SRMux
    port map (
            O => \N__25804\,
            I => \N__25617\
        );

    \I__6208\ : SRMux
    port map (
            O => \N__25803\,
            I => \N__25617\
        );

    \I__6207\ : SRMux
    port map (
            O => \N__25802\,
            I => \N__25617\
        );

    \I__6206\ : SRMux
    port map (
            O => \N__25801\,
            I => \N__25617\
        );

    \I__6205\ : SRMux
    port map (
            O => \N__25800\,
            I => \N__25617\
        );

    \I__6204\ : SRMux
    port map (
            O => \N__25799\,
            I => \N__25617\
        );

    \I__6203\ : Glb2LocalMux
    port map (
            O => \N__25796\,
            I => \N__25617\
        );

    \I__6202\ : Glb2LocalMux
    port map (
            O => \N__25793\,
            I => \N__25617\
        );

    \I__6201\ : Glb2LocalMux
    port map (
            O => \N__25790\,
            I => \N__25617\
        );

    \I__6200\ : Glb2LocalMux
    port map (
            O => \N__25787\,
            I => \N__25617\
        );

    \I__6199\ : Glb2LocalMux
    port map (
            O => \N__25784\,
            I => \N__25617\
        );

    \I__6198\ : Glb2LocalMux
    port map (
            O => \N__25781\,
            I => \N__25617\
        );

    \I__6197\ : SRMux
    port map (
            O => \N__25780\,
            I => \N__25617\
        );

    \I__6196\ : SRMux
    port map (
            O => \N__25779\,
            I => \N__25617\
        );

    \I__6195\ : SRMux
    port map (
            O => \N__25778\,
            I => \N__25617\
        );

    \I__6194\ : SRMux
    port map (
            O => \N__25777\,
            I => \N__25617\
        );

    \I__6193\ : SRMux
    port map (
            O => \N__25776\,
            I => \N__25617\
        );

    \I__6192\ : SRMux
    port map (
            O => \N__25775\,
            I => \N__25617\
        );

    \I__6191\ : SRMux
    port map (
            O => \N__25774\,
            I => \N__25617\
        );

    \I__6190\ : SRMux
    port map (
            O => \N__25773\,
            I => \N__25617\
        );

    \I__6189\ : SRMux
    port map (
            O => \N__25772\,
            I => \N__25617\
        );

    \I__6188\ : SRMux
    port map (
            O => \N__25771\,
            I => \N__25617\
        );

    \I__6187\ : SRMux
    port map (
            O => \N__25770\,
            I => \N__25617\
        );

    \I__6186\ : SRMux
    port map (
            O => \N__25769\,
            I => \N__25617\
        );

    \I__6185\ : SRMux
    port map (
            O => \N__25768\,
            I => \N__25617\
        );

    \I__6184\ : SRMux
    port map (
            O => \N__25767\,
            I => \N__25617\
        );

    \I__6183\ : SRMux
    port map (
            O => \N__25766\,
            I => \N__25617\
        );

    \I__6182\ : SRMux
    port map (
            O => \N__25765\,
            I => \N__25617\
        );

    \I__6181\ : Glb2LocalMux
    port map (
            O => \N__25762\,
            I => \N__25617\
        );

    \I__6180\ : Glb2LocalMux
    port map (
            O => \N__25759\,
            I => \N__25617\
        );

    \I__6179\ : Glb2LocalMux
    port map (
            O => \N__25756\,
            I => \N__25617\
        );

    \I__6178\ : GlobalMux
    port map (
            O => \N__25617\,
            I => \N__25614\
        );

    \I__6177\ : gio2CtrlBuf
    port map (
            O => \N__25614\,
            I => rst_g
        );

    \I__6176\ : IoInMux
    port map (
            O => \N__25611\,
            I => \N__25608\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__25608\,
            I => bu_rx_data_rdy_0
        );

    \I__6174\ : CascadeMux
    port map (
            O => \N__25605\,
            I => \Lab_UT.didp.countrce2.un13_qPone_cascade_\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__25602\,
            I => \Lab_UT.didp.countrce2.q_5_2_cascade_\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__25599\,
            I => \N__25595\
        );

    \I__6171\ : InMux
    port map (
            O => \N__25598\,
            I => \N__25590\
        );

    \I__6170\ : InMux
    port map (
            O => \N__25595\,
            I => \N__25590\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__25590\,
            I => \N__25583\
        );

    \I__6168\ : InMux
    port map (
            O => \N__25589\,
            I => \N__25580\
        );

    \I__6167\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25577\
        );

    \I__6166\ : InMux
    port map (
            O => \N__25587\,
            I => \N__25572\
        );

    \I__6165\ : InMux
    port map (
            O => \N__25586\,
            I => \N__25572\
        );

    \I__6164\ : Span4Mux_h
    port map (
            O => \N__25583\,
            I => \N__25569\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__25580\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__6162\ : LocalMux
    port map (
            O => \N__25577\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__25572\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__6160\ : Odrv4
    port map (
            O => \N__25569\,
            I => \Lab_UT.di_Stens_2\
        );

    \I__6159\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25550\
        );

    \I__6158\ : InMux
    port map (
            O => \N__25559\,
            I => \N__25543\
        );

    \I__6157\ : InMux
    port map (
            O => \N__25558\,
            I => \N__25543\
        );

    \I__6156\ : InMux
    port map (
            O => \N__25557\,
            I => \N__25543\
        );

    \I__6155\ : InMux
    port map (
            O => \N__25556\,
            I => \N__25534\
        );

    \I__6154\ : InMux
    port map (
            O => \N__25555\,
            I => \N__25534\
        );

    \I__6153\ : InMux
    port map (
            O => \N__25554\,
            I => \N__25534\
        );

    \I__6152\ : InMux
    port map (
            O => \N__25553\,
            I => \N__25534\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__25550\,
            I => \N__25531\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__25543\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__25534\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__6148\ : Odrv4
    port map (
            O => \N__25531\,
            I => \Lab_UT.di_Stens_0\
        );

    \I__6147\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25516\
        );

    \I__6146\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25513\
        );

    \I__6145\ : InMux
    port map (
            O => \N__25522\,
            I => \N__25510\
        );

    \I__6144\ : InMux
    port map (
            O => \N__25521\,
            I => \N__25507\
        );

    \I__6143\ : InMux
    port map (
            O => \N__25520\,
            I => \N__25504\
        );

    \I__6142\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25498\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__25516\,
            I => \N__25490\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__25513\,
            I => \N__25485\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25485\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__25507\,
            I => \N__25482\
        );

    \I__6137\ : LocalMux
    port map (
            O => \N__25504\,
            I => \N__25478\
        );

    \I__6136\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25475\
        );

    \I__6135\ : InMux
    port map (
            O => \N__25502\,
            I => \N__25470\
        );

    \I__6134\ : InMux
    port map (
            O => \N__25501\,
            I => \N__25470\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__25498\,
            I => \N__25467\
        );

    \I__6132\ : InMux
    port map (
            O => \N__25497\,
            I => \N__25458\
        );

    \I__6131\ : InMux
    port map (
            O => \N__25496\,
            I => \N__25458\
        );

    \I__6130\ : InMux
    port map (
            O => \N__25495\,
            I => \N__25458\
        );

    \I__6129\ : InMux
    port map (
            O => \N__25494\,
            I => \N__25458\
        );

    \I__6128\ : InMux
    port map (
            O => \N__25493\,
            I => \N__25453\
        );

    \I__6127\ : Span4Mux_v
    port map (
            O => \N__25490\,
            I => \N__25450\
        );

    \I__6126\ : Span4Mux_v
    port map (
            O => \N__25485\,
            I => \N__25447\
        );

    \I__6125\ : Span4Mux_v
    port map (
            O => \N__25482\,
            I => \N__25444\
        );

    \I__6124\ : InMux
    port map (
            O => \N__25481\,
            I => \N__25441\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__25478\,
            I => \N__25434\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__25475\,
            I => \N__25434\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__25470\,
            I => \N__25431\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__25467\,
            I => \N__25426\
        );

    \I__6119\ : LocalMux
    port map (
            O => \N__25458\,
            I => \N__25426\
        );

    \I__6118\ : InMux
    port map (
            O => \N__25457\,
            I => \N__25421\
        );

    \I__6117\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25421\
        );

    \I__6116\ : LocalMux
    port map (
            O => \N__25453\,
            I => \N__25418\
        );

    \I__6115\ : Sp12to4
    port map (
            O => \N__25450\,
            I => \N__25409\
        );

    \I__6114\ : Sp12to4
    port map (
            O => \N__25447\,
            I => \N__25409\
        );

    \I__6113\ : Sp12to4
    port map (
            O => \N__25444\,
            I => \N__25409\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__25441\,
            I => \N__25409\
        );

    \I__6111\ : CascadeMux
    port map (
            O => \N__25440\,
            I => \N__25405\
        );

    \I__6110\ : CascadeMux
    port map (
            O => \N__25439\,
            I => \N__25402\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__25434\,
            I => \N__25399\
        );

    \I__6108\ : Span4Mux_v
    port map (
            O => \N__25431\,
            I => \N__25394\
        );

    \I__6107\ : Span4Mux_h
    port map (
            O => \N__25426\,
            I => \N__25394\
        );

    \I__6106\ : LocalMux
    port map (
            O => \N__25421\,
            I => \N__25389\
        );

    \I__6105\ : Span12Mux_v
    port map (
            O => \N__25418\,
            I => \N__25389\
        );

    \I__6104\ : Span12Mux_s10_h
    port map (
            O => \N__25409\,
            I => \N__25386\
        );

    \I__6103\ : InMux
    port map (
            O => \N__25408\,
            I => \N__25379\
        );

    \I__6102\ : InMux
    port map (
            O => \N__25405\,
            I => \N__25379\
        );

    \I__6101\ : InMux
    port map (
            O => \N__25402\,
            I => \N__25379\
        );

    \I__6100\ : Span4Mux_v
    port map (
            O => \N__25399\,
            I => \N__25374\
        );

    \I__6099\ : Span4Mux_h
    port map (
            O => \N__25394\,
            I => \N__25374\
        );

    \I__6098\ : Odrv12
    port map (
            O => \N__25389\,
            I => bu_rx_data_1
        );

    \I__6097\ : Odrv12
    port map (
            O => \N__25386\,
            I => bu_rx_data_1
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__25379\,
            I => bu_rx_data_1
        );

    \I__6095\ : Odrv4
    port map (
            O => \N__25374\,
            I => bu_rx_data_1
        );

    \I__6094\ : InMux
    port map (
            O => \N__25365\,
            I => \N__25357\
        );

    \I__6093\ : InMux
    port map (
            O => \N__25364\,
            I => \N__25357\
        );

    \I__6092\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25354\
        );

    \I__6091\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25351\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__25357\,
            I => \N__25344\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__25354\,
            I => \N__25344\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__25351\,
            I => \N__25344\
        );

    \I__6087\ : Span4Mux_s1_h
    port map (
            O => \N__25344\,
            I => \N__25341\
        );

    \I__6086\ : Odrv4
    port map (
            O => \N__25341\,
            I => \Lab_UT.didp.un1_dicLdStens_0\
        );

    \I__6085\ : CascadeMux
    port map (
            O => \N__25338\,
            I => \Lab_UT.didp.countrce2.q_5_1_cascade_\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__25335\,
            I => \N__25332\
        );

    \I__6083\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25324\
        );

    \I__6082\ : InMux
    port map (
            O => \N__25331\,
            I => \N__25324\
        );

    \I__6081\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25321\
        );

    \I__6080\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25318\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__25324\,
            I => \N__25313\
        );

    \I__6078\ : LocalMux
    port map (
            O => \N__25321\,
            I => \N__25313\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__25318\,
            I => \N__25310\
        );

    \I__6076\ : Span4Mux_s1_h
    port map (
            O => \N__25313\,
            I => \N__25307\
        );

    \I__6075\ : Odrv4
    port map (
            O => \N__25310\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__25307\,
            I => \Lab_UT.didp.resetZ0Z_1\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__25302\,
            I => \N__25293\
        );

    \I__6072\ : InMux
    port map (
            O => \N__25301\,
            I => \N__25284\
        );

    \I__6071\ : InMux
    port map (
            O => \N__25300\,
            I => \N__25284\
        );

    \I__6070\ : InMux
    port map (
            O => \N__25299\,
            I => \N__25284\
        );

    \I__6069\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25284\
        );

    \I__6068\ : InMux
    port map (
            O => \N__25297\,
            I => \N__25277\
        );

    \I__6067\ : InMux
    port map (
            O => \N__25296\,
            I => \N__25277\
        );

    \I__6066\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25277\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__25284\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__25277\,
            I => \Lab_UT.di_Stens_1\
        );

    \I__6063\ : InMux
    port map (
            O => \N__25272\,
            I => \N__25269\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__25269\,
            I => \Lab_UT.didp.countrce2.un20_qPone\
        );

    \I__6061\ : CascadeMux
    port map (
            O => \N__25266\,
            I => \N__25261\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__25265\,
            I => \N__25257\
        );

    \I__6059\ : InMux
    port map (
            O => \N__25264\,
            I => \N__25252\
        );

    \I__6058\ : InMux
    port map (
            O => \N__25261\,
            I => \N__25252\
        );

    \I__6057\ : InMux
    port map (
            O => \N__25260\,
            I => \N__25249\
        );

    \I__6056\ : InMux
    port map (
            O => \N__25257\,
            I => \N__25246\
        );

    \I__6055\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25241\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__25249\,
            I => \N__25241\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__25246\,
            I => \N__25238\
        );

    \I__6052\ : Span4Mux_v
    port map (
            O => \N__25241\,
            I => \N__25235\
        );

    \I__6051\ : Span4Mux_s0_h
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__6050\ : Odrv4
    port map (
            O => \N__25235\,
            I => \Lab_UT.LdStens\
        );

    \I__6049\ : Odrv4
    port map (
            O => \N__25232\,
            I => \Lab_UT.LdStens\
        );

    \I__6048\ : CascadeMux
    port map (
            O => \N__25227\,
            I => \N__25223\
        );

    \I__6047\ : CascadeMux
    port map (
            O => \N__25226\,
            I => \N__25217\
        );

    \I__6046\ : InMux
    port map (
            O => \N__25223\,
            I => \N__25212\
        );

    \I__6045\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25212\
        );

    \I__6044\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25209\
        );

    \I__6043\ : InMux
    port map (
            O => \N__25220\,
            I => \N__25206\
        );

    \I__6042\ : InMux
    port map (
            O => \N__25217\,
            I => \N__25203\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__25212\,
            I => \N__25200\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__25209\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__25206\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__25203\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__6037\ : Odrv12
    port map (
            O => \N__25200\,
            I => \Lab_UT.di_Stens_3\
        );

    \I__6036\ : InMux
    port map (
            O => \N__25191\,
            I => \N__25188\
        );

    \I__6035\ : LocalMux
    port map (
            O => \N__25188\,
            I => \Lab_UT.didp.countrce2.q_5_3\
        );

    \I__6034\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25176\
        );

    \I__6033\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25176\
        );

    \I__6032\ : InMux
    port map (
            O => \N__25183\,
            I => \N__25176\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__25176\,
            I => \Lab_UT.didp.countrce3.ce_12_2_3\
        );

    \I__6030\ : CascadeMux
    port map (
            O => \N__25173\,
            I => \N__25164\
        );

    \I__6029\ : InMux
    port map (
            O => \N__25172\,
            I => \N__25157\
        );

    \I__6028\ : InMux
    port map (
            O => \N__25171\,
            I => \N__25157\
        );

    \I__6027\ : InMux
    port map (
            O => \N__25170\,
            I => \N__25154\
        );

    \I__6026\ : CascadeMux
    port map (
            O => \N__25169\,
            I => \N__25151\
        );

    \I__6025\ : CascadeMux
    port map (
            O => \N__25168\,
            I => \N__25148\
        );

    \I__6024\ : InMux
    port map (
            O => \N__25167\,
            I => \N__25143\
        );

    \I__6023\ : InMux
    port map (
            O => \N__25164\,
            I => \N__25143\
        );

    \I__6022\ : CascadeMux
    port map (
            O => \N__25163\,
            I => \N__25140\
        );

    \I__6021\ : CascadeMux
    port map (
            O => \N__25162\,
            I => \N__25137\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__25157\,
            I => \N__25131\
        );

    \I__6019\ : LocalMux
    port map (
            O => \N__25154\,
            I => \N__25131\
        );

    \I__6018\ : InMux
    port map (
            O => \N__25151\,
            I => \N__25126\
        );

    \I__6017\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25126\
        );

    \I__6016\ : LocalMux
    port map (
            O => \N__25143\,
            I => \N__25123\
        );

    \I__6015\ : InMux
    port map (
            O => \N__25140\,
            I => \N__25116\
        );

    \I__6014\ : InMux
    port map (
            O => \N__25137\,
            I => \N__25116\
        );

    \I__6013\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25116\
        );

    \I__6012\ : Span4Mux_s3_h
    port map (
            O => \N__25131\,
            I => \N__25113\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__25126\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__6010\ : Odrv4
    port map (
            O => \N__25123\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__6009\ : LocalMux
    port map (
            O => \N__25116\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__25113\,
            I => \uu2.w_addr_displayingZ0Z_8\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__25104\,
            I => \N__25097\
        );

    \I__6006\ : InMux
    port map (
            O => \N__25103\,
            I => \N__25094\
        );

    \I__6005\ : InMux
    port map (
            O => \N__25102\,
            I => \N__25091\
        );

    \I__6004\ : InMux
    port map (
            O => \N__25101\,
            I => \N__25080\
        );

    \I__6003\ : InMux
    port map (
            O => \N__25100\,
            I => \N__25080\
        );

    \I__6002\ : InMux
    port map (
            O => \N__25097\,
            I => \N__25080\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__25094\,
            I => \N__25071\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__25091\,
            I => \N__25071\
        );

    \I__5999\ : InMux
    port map (
            O => \N__25090\,
            I => \N__25068\
        );

    \I__5998\ : InMux
    port map (
            O => \N__25089\,
            I => \N__25061\
        );

    \I__5997\ : InMux
    port map (
            O => \N__25088\,
            I => \N__25061\
        );

    \I__5996\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25061\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__25080\,
            I => \N__25058\
        );

    \I__5994\ : InMux
    port map (
            O => \N__25079\,
            I => \N__25053\
        );

    \I__5993\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25053\
        );

    \I__5992\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25048\
        );

    \I__5991\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25048\
        );

    \I__5990\ : Span4Mux_s3_h
    port map (
            O => \N__25071\,
            I => \N__25043\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__25068\,
            I => \N__25043\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__25061\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__5987\ : Odrv4
    port map (
            O => \N__25058\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__25053\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__25048\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__25043\,
            I => \uu2.w_addr_displayingZ0Z_7\
        );

    \I__5983\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25021\
        );

    \I__5982\ : InMux
    port map (
            O => \N__25031\,
            I => \N__25021\
        );

    \I__5981\ : InMux
    port map (
            O => \N__25030\,
            I => \N__25021\
        );

    \I__5980\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25014\
        );

    \I__5979\ : InMux
    port map (
            O => \N__25028\,
            I => \N__25014\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__25021\,
            I => \N__25011\
        );

    \I__5977\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25008\
        );

    \I__5976\ : InMux
    port map (
            O => \N__25019\,
            I => \N__25005\
        );

    \I__5975\ : LocalMux
    port map (
            O => \N__25014\,
            I => \N__25002\
        );

    \I__5974\ : Span4Mux_s3_h
    port map (
            O => \N__25011\,
            I => \N__24995\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__25008\,
            I => \N__24992\
        );

    \I__5972\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24989\
        );

    \I__5971\ : Span4Mux_s2_v
    port map (
            O => \N__25002\,
            I => \N__24986\
        );

    \I__5970\ : InMux
    port map (
            O => \N__25001\,
            I => \N__24977\
        );

    \I__5969\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24977\
        );

    \I__5968\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24977\
        );

    \I__5967\ : InMux
    port map (
            O => \N__24998\,
            I => \N__24977\
        );

    \I__5966\ : Odrv4
    port map (
            O => \N__24995\,
            I => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\
        );

    \I__5965\ : Odrv4
    port map (
            O => \N__24992\,
            I => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\
        );

    \I__5964\ : Odrv4
    port map (
            O => \N__24989\,
            I => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__24986\,
            I => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__24977\,
            I => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\
        );

    \I__5961\ : CascadeMux
    port map (
            O => \N__24966\,
            I => \uu2.N_33_cascade_\
        );

    \I__5960\ : InMux
    port map (
            O => \N__24963\,
            I => \N__24960\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__24960\,
            I => \uu2.N_14_i\
        );

    \I__5958\ : InMux
    port map (
            O => \N__24957\,
            I => \N__24947\
        );

    \I__5957\ : InMux
    port map (
            O => \N__24956\,
            I => \N__24947\
        );

    \I__5956\ : InMux
    port map (
            O => \N__24955\,
            I => \N__24947\
        );

    \I__5955\ : CascadeMux
    port map (
            O => \N__24954\,
            I => \N__24944\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__24947\,
            I => \N__24941\
        );

    \I__5953\ : InMux
    port map (
            O => \N__24944\,
            I => \N__24938\
        );

    \I__5952\ : Span4Mux_s0_v
    port map (
            O => \N__24941\,
            I => \N__24933\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__24938\,
            I => \N__24930\
        );

    \I__5950\ : InMux
    port map (
            O => \N__24937\,
            I => \N__24927\
        );

    \I__5949\ : InMux
    port map (
            O => \N__24936\,
            I => \N__24924\
        );

    \I__5948\ : Span4Mux_h
    port map (
            O => \N__24933\,
            I => \N__24921\
        );

    \I__5947\ : Span4Mux_s1_v
    port map (
            O => \N__24930\,
            I => \N__24918\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__24927\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__24924\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__5944\ : Odrv4
    port map (
            O => \N__24921\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__5943\ : Odrv4
    port map (
            O => \N__24918\,
            I => \uu2.w_addr_displayingZ0Z_6\
        );

    \I__5942\ : InMux
    port map (
            O => \N__24909\,
            I => \N__24906\
        );

    \I__5941\ : LocalMux
    port map (
            O => \N__24906\,
            I => \N__24903\
        );

    \I__5940\ : Odrv12
    port map (
            O => \N__24903\,
            I => \uu2.bitmapZ0Z_212\
        );

    \I__5939\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24897\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__24897\,
            I => \uu2.bitmapZ0Z_180\
        );

    \I__5937\ : InMux
    port map (
            O => \N__24894\,
            I => \N__24886\
        );

    \I__5936\ : InMux
    port map (
            O => \N__24893\,
            I => \N__24883\
        );

    \I__5935\ : InMux
    port map (
            O => \N__24892\,
            I => \N__24878\
        );

    \I__5934\ : InMux
    port map (
            O => \N__24891\,
            I => \N__24878\
        );

    \I__5933\ : InMux
    port map (
            O => \N__24890\,
            I => \N__24875\
        );

    \I__5932\ : InMux
    port map (
            O => \N__24889\,
            I => \N__24872\
        );

    \I__5931\ : LocalMux
    port map (
            O => \N__24886\,
            I => \N__24869\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N__24864\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__24878\,
            I => \N__24864\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__24875\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__24872\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__5926\ : Odrv4
    port map (
            O => \N__24869\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__5925\ : Odrv12
    port map (
            O => \N__24864\,
            I => \uu2.w_addr_displaying_fastZ0Z_8\
        );

    \I__5924\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__24852\,
            I => \uu2.bitmapZ0Z_52\
        );

    \I__5922\ : InMux
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__5921\ : LocalMux
    port map (
            O => \N__24846\,
            I => \uu2.bitmapZ0Z_308\
        );

    \I__5920\ : InMux
    port map (
            O => \N__24843\,
            I => \N__24840\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__24840\,
            I => \uu2.N_194\
        );

    \I__5918\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24834\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24831\
        );

    \I__5916\ : Odrv4
    port map (
            O => \N__24831\,
            I => \uu2.bitmapZ0Z_87\
        );

    \I__5915\ : InMux
    port map (
            O => \N__24828\,
            I => \N__24825\
        );

    \I__5914\ : LocalMux
    port map (
            O => \N__24825\,
            I => \N__24821\
        );

    \I__5913\ : InMux
    port map (
            O => \N__24824\,
            I => \N__24817\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__24821\,
            I => \N__24814\
        );

    \I__5911\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24811\
        );

    \I__5910\ : LocalMux
    port map (
            O => \N__24817\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__5909\ : Odrv4
    port map (
            O => \N__24814\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__24811\,
            I => \uu2.w_addr_displaying_fastZ0Z_0\
        );

    \I__5907\ : InMux
    port map (
            O => \N__24804\,
            I => \N__24801\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__24801\,
            I => \N__24798\
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__24798\,
            I => \uu2.N_197\
        );

    \I__5904\ : CascadeMux
    port map (
            O => \N__24795\,
            I => \N__24791\
        );

    \I__5903\ : CascadeMux
    port map (
            O => \N__24794\,
            I => \N__24788\
        );

    \I__5902\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24779\
        );

    \I__5901\ : InMux
    port map (
            O => \N__24788\,
            I => \N__24779\
        );

    \I__5900\ : InMux
    port map (
            O => \N__24787\,
            I => \N__24776\
        );

    \I__5899\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24769\
        );

    \I__5898\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24769\
        );

    \I__5897\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24769\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__24779\,
            I => \N__24765\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24760\
        );

    \I__5894\ : LocalMux
    port map (
            O => \N__24769\,
            I => \N__24760\
        );

    \I__5893\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24757\
        );

    \I__5892\ : Span4Mux_s2_h
    port map (
            O => \N__24765\,
            I => \N__24754\
        );

    \I__5891\ : Span4Mux_s2_h
    port map (
            O => \N__24760\,
            I => \N__24751\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__24757\,
            I => \N__24748\
        );

    \I__5889\ : Odrv4
    port map (
            O => \N__24754\,
            I => \Lab_UT.sec1_2\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__24751\,
            I => \Lab_UT.sec1_2\
        );

    \I__5887\ : Odrv12
    port map (
            O => \N__24748\,
            I => \Lab_UT.sec1_2\
        );

    \I__5886\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24736\
        );

    \I__5885\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24731\
        );

    \I__5884\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24731\
        );

    \I__5883\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24727\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__24731\,
            I => \N__24724\
        );

    \I__5881\ : CascadeMux
    port map (
            O => \N__24730\,
            I => \N__24720\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__24727\,
            I => \N__24713\
        );

    \I__5879\ : Span4Mux_s0_h
    port map (
            O => \N__24724\,
            I => \N__24713\
        );

    \I__5878\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24710\
        );

    \I__5877\ : InMux
    port map (
            O => \N__24720\,
            I => \N__24703\
        );

    \I__5876\ : InMux
    port map (
            O => \N__24719\,
            I => \N__24703\
        );

    \I__5875\ : InMux
    port map (
            O => \N__24718\,
            I => \N__24703\
        );

    \I__5874\ : Odrv4
    port map (
            O => \N__24713\,
            I => \Lab_UT.sec1_1\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__24710\,
            I => \Lab_UT.sec1_1\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__24703\,
            I => \Lab_UT.sec1_1\
        );

    \I__5871\ : CascadeMux
    port map (
            O => \N__24696\,
            I => \N__24688\
        );

    \I__5870\ : CascadeMux
    port map (
            O => \N__24695\,
            I => \N__24684\
        );

    \I__5869\ : CascadeMux
    port map (
            O => \N__24694\,
            I => \N__24681\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__24693\,
            I => \N__24678\
        );

    \I__5867\ : InMux
    port map (
            O => \N__24692\,
            I => \N__24673\
        );

    \I__5866\ : InMux
    port map (
            O => \N__24691\,
            I => \N__24673\
        );

    \I__5865\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24670\
        );

    \I__5864\ : InMux
    port map (
            O => \N__24687\,
            I => \N__24663\
        );

    \I__5863\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24663\
        );

    \I__5862\ : InMux
    port map (
            O => \N__24681\,
            I => \N__24663\
        );

    \I__5861\ : InMux
    port map (
            O => \N__24678\,
            I => \N__24660\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__24673\,
            I => \N__24657\
        );

    \I__5859\ : LocalMux
    port map (
            O => \N__24670\,
            I => \N__24652\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__24663\,
            I => \N__24652\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__24660\,
            I => \N__24649\
        );

    \I__5856\ : Span12Mux_s4_h
    port map (
            O => \N__24657\,
            I => \N__24646\
        );

    \I__5855\ : Span4Mux_s3_h
    port map (
            O => \N__24652\,
            I => \N__24641\
        );

    \I__5854\ : Span4Mux_s3_v
    port map (
            O => \N__24649\,
            I => \N__24641\
        );

    \I__5853\ : Odrv12
    port map (
            O => \N__24646\,
            I => \Lab_UT.sec1_3\
        );

    \I__5852\ : Odrv4
    port map (
            O => \N__24641\,
            I => \Lab_UT.sec1_3\
        );

    \I__5851\ : InMux
    port map (
            O => \N__24636\,
            I => \N__24633\
        );

    \I__5850\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24628\
        );

    \I__5849\ : InMux
    port map (
            O => \N__24632\,
            I => \N__24623\
        );

    \I__5848\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24623\
        );

    \I__5847\ : Span4Mux_v
    port map (
            O => \N__24628\,
            I => \N__24616\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__24623\,
            I => \N__24613\
        );

    \I__5845\ : InMux
    port map (
            O => \N__24622\,
            I => \N__24610\
        );

    \I__5844\ : InMux
    port map (
            O => \N__24621\,
            I => \N__24603\
        );

    \I__5843\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24603\
        );

    \I__5842\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24603\
        );

    \I__5841\ : Odrv4
    port map (
            O => \N__24616\,
            I => \Lab_UT.sec1_0\
        );

    \I__5840\ : Odrv4
    port map (
            O => \N__24613\,
            I => \Lab_UT.sec1_0\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__24610\,
            I => \Lab_UT.sec1_0\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__24603\,
            I => \Lab_UT.sec1_0\
        );

    \I__5837\ : InMux
    port map (
            O => \N__24594\,
            I => \N__24591\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__24591\,
            I => \uu2.bitmapZ0Z_84\
        );

    \I__5835\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24579\
        );

    \I__5833\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24571\
        );

    \I__5832\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24571\
        );

    \I__5831\ : InMux
    port map (
            O => \N__24582\,
            I => \N__24571\
        );

    \I__5830\ : Span4Mux_s3_v
    port map (
            O => \N__24579\,
            I => \N__24568\
        );

    \I__5829\ : InMux
    port map (
            O => \N__24578\,
            I => \N__24565\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__24571\,
            I => \N__24562\
        );

    \I__5827\ : Odrv4
    port map (
            O => \N__24568\,
            I => \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__24565\,
            I => \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0\
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__24562\,
            I => \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0\
        );

    \I__5824\ : CascadeMux
    port map (
            O => \N__24555\,
            I => \N__24548\
        );

    \I__5823\ : CascadeMux
    port map (
            O => \N__24554\,
            I => \N__24540\
        );

    \I__5822\ : CascadeMux
    port map (
            O => \N__24553\,
            I => \N__24537\
        );

    \I__5821\ : InMux
    port map (
            O => \N__24552\,
            I => \N__24528\
        );

    \I__5820\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24528\
        );

    \I__5819\ : InMux
    port map (
            O => \N__24548\,
            I => \N__24525\
        );

    \I__5818\ : CascadeMux
    port map (
            O => \N__24547\,
            I => \N__24518\
        );

    \I__5817\ : InMux
    port map (
            O => \N__24546\,
            I => \N__24515\
        );

    \I__5816\ : InMux
    port map (
            O => \N__24545\,
            I => \N__24512\
        );

    \I__5815\ : InMux
    port map (
            O => \N__24544\,
            I => \N__24509\
        );

    \I__5814\ : InMux
    port map (
            O => \N__24543\,
            I => \N__24504\
        );

    \I__5813\ : InMux
    port map (
            O => \N__24540\,
            I => \N__24504\
        );

    \I__5812\ : InMux
    port map (
            O => \N__24537\,
            I => \N__24501\
        );

    \I__5811\ : InMux
    port map (
            O => \N__24536\,
            I => \N__24498\
        );

    \I__5810\ : InMux
    port map (
            O => \N__24535\,
            I => \N__24495\
        );

    \I__5809\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24492\
        );

    \I__5808\ : CascadeMux
    port map (
            O => \N__24533\,
            I => \N__24486\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__24528\,
            I => \N__24481\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__24525\,
            I => \N__24478\
        );

    \I__5805\ : InMux
    port map (
            O => \N__24524\,
            I => \N__24469\
        );

    \I__5804\ : InMux
    port map (
            O => \N__24523\,
            I => \N__24469\
        );

    \I__5803\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24469\
        );

    \I__5802\ : InMux
    port map (
            O => \N__24521\,
            I => \N__24469\
        );

    \I__5801\ : InMux
    port map (
            O => \N__24518\,
            I => \N__24466\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24463\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__24512\,
            I => \N__24460\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24451\
        );

    \I__5797\ : LocalMux
    port map (
            O => \N__24504\,
            I => \N__24451\
        );

    \I__5796\ : LocalMux
    port map (
            O => \N__24501\,
            I => \N__24451\
        );

    \I__5795\ : LocalMux
    port map (
            O => \N__24498\,
            I => \N__24446\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__24495\,
            I => \N__24446\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__24492\,
            I => \N__24443\
        );

    \I__5792\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24438\
        );

    \I__5791\ : InMux
    port map (
            O => \N__24490\,
            I => \N__24438\
        );

    \I__5790\ : InMux
    port map (
            O => \N__24489\,
            I => \N__24433\
        );

    \I__5789\ : InMux
    port map (
            O => \N__24486\,
            I => \N__24433\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24485\,
            I => \N__24430\
        );

    \I__5787\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24427\
        );

    \I__5786\ : Span4Mux_s2_v
    port map (
            O => \N__24481\,
            I => \N__24420\
        );

    \I__5785\ : Span4Mux_h
    port map (
            O => \N__24478\,
            I => \N__24420\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__24469\,
            I => \N__24420\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__24466\,
            I => \N__24417\
        );

    \I__5782\ : Span4Mux_s2_v
    port map (
            O => \N__24463\,
            I => \N__24414\
        );

    \I__5781\ : Span4Mux_h
    port map (
            O => \N__24460\,
            I => \N__24411\
        );

    \I__5780\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24406\
        );

    \I__5779\ : InMux
    port map (
            O => \N__24458\,
            I => \N__24406\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__24451\,
            I => \N__24401\
        );

    \I__5777\ : Span4Mux_h
    port map (
            O => \N__24446\,
            I => \N__24401\
        );

    \I__5776\ : Span4Mux_s3_v
    port map (
            O => \N__24443\,
            I => \N__24394\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__24438\,
            I => \N__24394\
        );

    \I__5774\ : LocalMux
    port map (
            O => \N__24433\,
            I => \N__24394\
        );

    \I__5773\ : LocalMux
    port map (
            O => \N__24430\,
            I => \N__24383\
        );

    \I__5772\ : LocalMux
    port map (
            O => \N__24427\,
            I => \N__24383\
        );

    \I__5771\ : Span4Mux_v
    port map (
            O => \N__24420\,
            I => \N__24383\
        );

    \I__5770\ : Span4Mux_v
    port map (
            O => \N__24417\,
            I => \N__24383\
        );

    \I__5769\ : Span4Mux_v
    port map (
            O => \N__24414\,
            I => \N__24383\
        );

    \I__5768\ : Odrv4
    port map (
            O => \N__24411\,
            I => \Lab_UT.state_3\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__24406\,
            I => \Lab_UT.state_3\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__24401\,
            I => \Lab_UT.state_3\
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__24394\,
            I => \Lab_UT.state_3\
        );

    \I__5764\ : Odrv4
    port map (
            O => \N__24383\,
            I => \Lab_UT.state_3\
        );

    \I__5763\ : InMux
    port map (
            O => \N__24372\,
            I => \N__24369\
        );

    \I__5762\ : LocalMux
    port map (
            O => \N__24369\,
            I => \N__24365\
        );

    \I__5761\ : InMux
    port map (
            O => \N__24368\,
            I => \N__24362\
        );

    \I__5760\ : Span4Mux_v
    port map (
            O => \N__24365\,
            I => \N__24357\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__24362\,
            I => \N__24357\
        );

    \I__5758\ : Span4Mux_h
    port map (
            O => \N__24357\,
            I => \N__24354\
        );

    \I__5757\ : Odrv4
    port map (
            O => \N__24354\,
            I => \Lab_UT.dictrl.N_40_1\
        );

    \I__5756\ : InMux
    port map (
            O => \N__24351\,
            I => \N__24348\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__24348\,
            I => \Lab_UT.dictrl.g1\
        );

    \I__5754\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24342\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__24342\,
            I => \N__24338\
        );

    \I__5752\ : InMux
    port map (
            O => \N__24341\,
            I => \N__24335\
        );

    \I__5751\ : Span4Mux_h
    port map (
            O => \N__24338\,
            I => \N__24332\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24329\
        );

    \I__5749\ : Odrv4
    port map (
            O => \N__24332\,
            I => \Lab_UT.dictrl.N_97_mux_4\
        );

    \I__5748\ : Odrv4
    port map (
            O => \N__24329\,
            I => \Lab_UT.dictrl.N_97_mux_4\
        );

    \I__5747\ : InMux
    port map (
            O => \N__24324\,
            I => \N__24313\
        );

    \I__5746\ : CascadeMux
    port map (
            O => \N__24323\,
            I => \N__24310\
        );

    \I__5745\ : InMux
    port map (
            O => \N__24322\,
            I => \N__24300\
        );

    \I__5744\ : InMux
    port map (
            O => \N__24321\,
            I => \N__24295\
        );

    \I__5743\ : InMux
    port map (
            O => \N__24320\,
            I => \N__24295\
        );

    \I__5742\ : InMux
    port map (
            O => \N__24319\,
            I => \N__24283\
        );

    \I__5741\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24283\
        );

    \I__5740\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24283\
        );

    \I__5739\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24283\
        );

    \I__5738\ : LocalMux
    port map (
            O => \N__24313\,
            I => \N__24280\
        );

    \I__5737\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24272\
        );

    \I__5736\ : InMux
    port map (
            O => \N__24309\,
            I => \N__24272\
        );

    \I__5735\ : InMux
    port map (
            O => \N__24308\,
            I => \N__24268\
        );

    \I__5734\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24265\
        );

    \I__5733\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24262\
        );

    \I__5732\ : InMux
    port map (
            O => \N__24305\,
            I => \N__24259\
        );

    \I__5731\ : InMux
    port map (
            O => \N__24304\,
            I => \N__24254\
        );

    \I__5730\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24254\
        );

    \I__5729\ : LocalMux
    port map (
            O => \N__24300\,
            I => \N__24249\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__24295\,
            I => \N__24249\
        );

    \I__5727\ : InMux
    port map (
            O => \N__24294\,
            I => \N__24246\
        );

    \I__5726\ : InMux
    port map (
            O => \N__24293\,
            I => \N__24243\
        );

    \I__5725\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24240\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24237\
        );

    \I__5723\ : Span4Mux_s2_v
    port map (
            O => \N__24280\,
            I => \N__24234\
        );

    \I__5722\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24229\
        );

    \I__5721\ : InMux
    port map (
            O => \N__24278\,
            I => \N__24229\
        );

    \I__5720\ : InMux
    port map (
            O => \N__24277\,
            I => \N__24226\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__24272\,
            I => \N__24223\
        );

    \I__5718\ : InMux
    port map (
            O => \N__24271\,
            I => \N__24220\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__24268\,
            I => \N__24217\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N__24210\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__24262\,
            I => \N__24210\
        );

    \I__5714\ : LocalMux
    port map (
            O => \N__24259\,
            I => \N__24210\
        );

    \I__5713\ : LocalMux
    port map (
            O => \N__24254\,
            I => \N__24201\
        );

    \I__5712\ : Span4Mux_h
    port map (
            O => \N__24249\,
            I => \N__24201\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__24246\,
            I => \N__24201\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__24243\,
            I => \N__24201\
        );

    \I__5709\ : LocalMux
    port map (
            O => \N__24240\,
            I => \N__24196\
        );

    \I__5708\ : Span4Mux_s3_h
    port map (
            O => \N__24237\,
            I => \N__24196\
        );

    \I__5707\ : Span4Mux_v
    port map (
            O => \N__24234\,
            I => \N__24191\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24191\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__24226\,
            I => \N__24186\
        );

    \I__5704\ : Span4Mux_s3_h
    port map (
            O => \N__24223\,
            I => \N__24186\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__24220\,
            I => \N__24183\
        );

    \I__5702\ : Span4Mux_v
    port map (
            O => \N__24217\,
            I => \N__24178\
        );

    \I__5701\ : Span4Mux_v
    port map (
            O => \N__24210\,
            I => \N__24178\
        );

    \I__5700\ : Span4Mux_v
    port map (
            O => \N__24201\,
            I => \N__24173\
        );

    \I__5699\ : Span4Mux_h
    port map (
            O => \N__24196\,
            I => \N__24173\
        );

    \I__5698\ : Odrv4
    port map (
            O => \N__24191\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5697\ : Odrv4
    port map (
            O => \N__24186\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5696\ : Odrv12
    port map (
            O => \N__24183\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5695\ : Odrv4
    port map (
            O => \N__24178\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5694\ : Odrv4
    port map (
            O => \N__24173\,
            I => \Lab_UT.dictrl.stateZ0Z_0\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__24162\,
            I => \N__24159\
        );

    \I__5692\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24156\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__24156\,
            I => \N__24153\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__24153\,
            I => \N__24150\
        );

    \I__5689\ : Odrv4
    port map (
            O => \N__24150\,
            I => \Lab_UT.dictrl.g1_1_1\
        );

    \I__5688\ : InMux
    port map (
            O => \N__24147\,
            I => \N__24141\
        );

    \I__5687\ : InMux
    port map (
            O => \N__24146\,
            I => \N__24136\
        );

    \I__5686\ : InMux
    port map (
            O => \N__24145\,
            I => \N__24136\
        );

    \I__5685\ : InMux
    port map (
            O => \N__24144\,
            I => \N__24133\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__24141\,
            I => \N__24130\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__24136\,
            I => \N__24127\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__24133\,
            I => \N__24122\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__24130\,
            I => \N__24122\
        );

    \I__5680\ : Span4Mux_s3_h
    port map (
            O => \N__24127\,
            I => \N__24119\
        );

    \I__5679\ : Span4Mux_h
    port map (
            O => \N__24122\,
            I => \N__24116\
        );

    \I__5678\ : Span4Mux_h
    port map (
            O => \N__24119\,
            I => \N__24113\
        );

    \I__5677\ : Odrv4
    port map (
            O => \N__24116\,
            I => \Lab_UT.dictrl.m34_4\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__24113\,
            I => \Lab_UT.dictrl.m34_4\
        );

    \I__5675\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24105\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24102\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__24102\,
            I => \Lab_UT.dictrl.N_1106_0\
        );

    \I__5672\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24096\
        );

    \I__5671\ : LocalMux
    port map (
            O => \N__24096\,
            I => \N__24093\
        );

    \I__5670\ : Span4Mux_s2_v
    port map (
            O => \N__24093\,
            I => \N__24090\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__24090\,
            I => \Lab_UT.dictrl.N_1462_1\
        );

    \I__5668\ : InMux
    port map (
            O => \N__24087\,
            I => \N__24084\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__24084\,
            I => \N__24081\
        );

    \I__5666\ : Span4Mux_s3_h
    port map (
            O => \N__24081\,
            I => \N__24078\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__24078\,
            I => \Lab_UT.dictrl.N_1102_1\
        );

    \I__5664\ : CascadeMux
    port map (
            O => \N__24075\,
            I => \N__24072\
        );

    \I__5663\ : InMux
    port map (
            O => \N__24072\,
            I => \N__24069\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__24069\,
            I => \N__24066\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__24066\,
            I => \Lab_UT.dictrl.g2_1_1\
        );

    \I__5660\ : InMux
    port map (
            O => \N__24063\,
            I => \N__24059\
        );

    \I__5659\ : InMux
    port map (
            O => \N__24062\,
            I => \N__24045\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__24059\,
            I => \N__24042\
        );

    \I__5657\ : CascadeMux
    port map (
            O => \N__24058\,
            I => \N__24027\
        );

    \I__5656\ : CascadeMux
    port map (
            O => \N__24057\,
            I => \N__24024\
        );

    \I__5655\ : InMux
    port map (
            O => \N__24056\,
            I => \N__24021\
        );

    \I__5654\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24018\
        );

    \I__5653\ : CascadeMux
    port map (
            O => \N__24054\,
            I => \N__24008\
        );

    \I__5652\ : CascadeMux
    port map (
            O => \N__24053\,
            I => \N__24005\
        );

    \I__5651\ : CascadeMux
    port map (
            O => \N__24052\,
            I => \N__23994\
        );

    \I__5650\ : CascadeMux
    port map (
            O => \N__24051\,
            I => \N__23991\
        );

    \I__5649\ : CascadeMux
    port map (
            O => \N__24050\,
            I => \N__23988\
        );

    \I__5648\ : CascadeMux
    port map (
            O => \N__24049\,
            I => \N__23985\
        );

    \I__5647\ : InMux
    port map (
            O => \N__24048\,
            I => \N__23978\
        );

    \I__5646\ : LocalMux
    port map (
            O => \N__24045\,
            I => \N__23975\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__24042\,
            I => \N__23972\
        );

    \I__5644\ : InMux
    port map (
            O => \N__24041\,
            I => \N__23969\
        );

    \I__5643\ : InMux
    port map (
            O => \N__24040\,
            I => \N__23959\
        );

    \I__5642\ : InMux
    port map (
            O => \N__24039\,
            I => \N__23955\
        );

    \I__5641\ : InMux
    port map (
            O => \N__24038\,
            I => \N__23940\
        );

    \I__5640\ : InMux
    port map (
            O => \N__24037\,
            I => \N__23940\
        );

    \I__5639\ : InMux
    port map (
            O => \N__24036\,
            I => \N__23940\
        );

    \I__5638\ : InMux
    port map (
            O => \N__24035\,
            I => \N__23940\
        );

    \I__5637\ : InMux
    port map (
            O => \N__24034\,
            I => \N__23940\
        );

    \I__5636\ : InMux
    port map (
            O => \N__24033\,
            I => \N__23940\
        );

    \I__5635\ : InMux
    port map (
            O => \N__24032\,
            I => \N__23940\
        );

    \I__5634\ : InMux
    port map (
            O => \N__24031\,
            I => \N__23935\
        );

    \I__5633\ : InMux
    port map (
            O => \N__24030\,
            I => \N__23935\
        );

    \I__5632\ : InMux
    port map (
            O => \N__24027\,
            I => \N__23930\
        );

    \I__5631\ : InMux
    port map (
            O => \N__24024\,
            I => \N__23930\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__24021\,
            I => \N__23925\
        );

    \I__5629\ : LocalMux
    port map (
            O => \N__24018\,
            I => \N__23925\
        );

    \I__5628\ : InMux
    port map (
            O => \N__24017\,
            I => \N__23922\
        );

    \I__5627\ : InMux
    port map (
            O => \N__24016\,
            I => \N__23919\
        );

    \I__5626\ : InMux
    port map (
            O => \N__24015\,
            I => \N__23912\
        );

    \I__5625\ : InMux
    port map (
            O => \N__24014\,
            I => \N__23912\
        );

    \I__5624\ : InMux
    port map (
            O => \N__24013\,
            I => \N__23912\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__24012\,
            I => \N__23906\
        );

    \I__5622\ : InMux
    port map (
            O => \N__24011\,
            I => \N__23902\
        );

    \I__5621\ : InMux
    port map (
            O => \N__24008\,
            I => \N__23893\
        );

    \I__5620\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23893\
        );

    \I__5619\ : InMux
    port map (
            O => \N__24004\,
            I => \N__23893\
        );

    \I__5618\ : InMux
    port map (
            O => \N__24003\,
            I => \N__23893\
        );

    \I__5617\ : InMux
    port map (
            O => \N__24002\,
            I => \N__23890\
        );

    \I__5616\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23883\
        );

    \I__5615\ : InMux
    port map (
            O => \N__24000\,
            I => \N__23883\
        );

    \I__5614\ : InMux
    port map (
            O => \N__23999\,
            I => \N__23883\
        );

    \I__5613\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23876\
        );

    \I__5612\ : InMux
    port map (
            O => \N__23997\,
            I => \N__23876\
        );

    \I__5611\ : InMux
    port map (
            O => \N__23994\,
            I => \N__23876\
        );

    \I__5610\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23869\
        );

    \I__5609\ : InMux
    port map (
            O => \N__23988\,
            I => \N__23869\
        );

    \I__5608\ : InMux
    port map (
            O => \N__23985\,
            I => \N__23869\
        );

    \I__5607\ : InMux
    port map (
            O => \N__23984\,
            I => \N__23866\
        );

    \I__5606\ : InMux
    port map (
            O => \N__23983\,
            I => \N__23859\
        );

    \I__5605\ : InMux
    port map (
            O => \N__23982\,
            I => \N__23859\
        );

    \I__5604\ : InMux
    port map (
            O => \N__23981\,
            I => \N__23859\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23978\,
            I => \N__23854\
        );

    \I__5602\ : Span4Mux_v
    port map (
            O => \N__23975\,
            I => \N__23854\
        );

    \I__5601\ : IoSpan4Mux
    port map (
            O => \N__23972\,
            I => \N__23849\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__23969\,
            I => \N__23849\
        );

    \I__5599\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23840\
        );

    \I__5598\ : InMux
    port map (
            O => \N__23967\,
            I => \N__23840\
        );

    \I__5597\ : InMux
    port map (
            O => \N__23966\,
            I => \N__23840\
        );

    \I__5596\ : InMux
    port map (
            O => \N__23965\,
            I => \N__23840\
        );

    \I__5595\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23833\
        );

    \I__5594\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23833\
        );

    \I__5593\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23833\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23830\
        );

    \I__5591\ : InMux
    port map (
            O => \N__23958\,
            I => \N__23824\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__23955\,
            I => \N__23821\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__23940\,
            I => \N__23818\
        );

    \I__5588\ : LocalMux
    port map (
            O => \N__23935\,
            I => \N__23805\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__23930\,
            I => \N__23805\
        );

    \I__5586\ : Span4Mux_h
    port map (
            O => \N__23925\,
            I => \N__23805\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23922\,
            I => \N__23805\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__23919\,
            I => \N__23805\
        );

    \I__5583\ : LocalMux
    port map (
            O => \N__23912\,
            I => \N__23805\
        );

    \I__5582\ : InMux
    port map (
            O => \N__23911\,
            I => \N__23802\
        );

    \I__5581\ : InMux
    port map (
            O => \N__23910\,
            I => \N__23793\
        );

    \I__5580\ : InMux
    port map (
            O => \N__23909\,
            I => \N__23793\
        );

    \I__5579\ : InMux
    port map (
            O => \N__23906\,
            I => \N__23793\
        );

    \I__5578\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23793\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23790\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__23893\,
            I => \N__23783\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__23890\,
            I => \N__23783\
        );

    \I__5574\ : LocalMux
    port map (
            O => \N__23883\,
            I => \N__23783\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__23876\,
            I => \N__23776\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23776\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__23866\,
            I => \N__23776\
        );

    \I__5570\ : LocalMux
    port map (
            O => \N__23859\,
            I => \N__23769\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__23854\,
            I => \N__23769\
        );

    \I__5568\ : Span4Mux_s2_v
    port map (
            O => \N__23849\,
            I => \N__23769\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__23840\,
            I => \N__23762\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23762\
        );

    \I__5565\ : Span4Mux_s2_v
    port map (
            O => \N__23830\,
            I => \N__23762\
        );

    \I__5564\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23759\
        );

    \I__5563\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23754\
        );

    \I__5562\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23754\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23749\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__23821\,
            I => \N__23749\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__23818\,
            I => \N__23744\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__23805\,
            I => \N__23744\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__23802\,
            I => \N__23735\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__23793\,
            I => \N__23735\
        );

    \I__5555\ : Span12Mux_s4_h
    port map (
            O => \N__23790\,
            I => \N__23735\
        );

    \I__5554\ : Span12Mux_s5_v
    port map (
            O => \N__23783\,
            I => \N__23735\
        );

    \I__5553\ : Span4Mux_h
    port map (
            O => \N__23776\,
            I => \N__23728\
        );

    \I__5552\ : Span4Mux_h
    port map (
            O => \N__23769\,
            I => \N__23728\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__23762\,
            I => \N__23728\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23759\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__23754\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__23749\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5547\ : Odrv4
    port map (
            O => \N__23744\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5546\ : Odrv12
    port map (
            O => \N__23735\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5545\ : Odrv4
    port map (
            O => \N__23728\,
            I => \Lab_UT.dictrl.un1_next_state66_0\
        );

    \I__5544\ : InMux
    port map (
            O => \N__23715\,
            I => \N__23712\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__23712\,
            I => \N__23709\
        );

    \I__5542\ : Odrv12
    port map (
            O => \N__23709\,
            I => \Lab_UT.dictrl.N_1460_1\
        );

    \I__5541\ : CascadeMux
    port map (
            O => \N__23706\,
            I => \N__23701\
        );

    \I__5540\ : CascadeMux
    port map (
            O => \N__23705\,
            I => \N__23698\
        );

    \I__5539\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23694\
        );

    \I__5538\ : InMux
    port map (
            O => \N__23701\,
            I => \N__23684\
        );

    \I__5537\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23684\
        );

    \I__5536\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23684\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__23694\,
            I => \N__23681\
        );

    \I__5534\ : CascadeMux
    port map (
            O => \N__23693\,
            I => \N__23677\
        );

    \I__5533\ : CascadeMux
    port map (
            O => \N__23692\,
            I => \N__23673\
        );

    \I__5532\ : CascadeMux
    port map (
            O => \N__23691\,
            I => \N__23670\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__23684\,
            I => \N__23663\
        );

    \I__5530\ : Span4Mux_s2_h
    port map (
            O => \N__23681\,
            I => \N__23663\
        );

    \I__5529\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23655\
        );

    \I__5528\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23655\
        );

    \I__5527\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23655\
        );

    \I__5526\ : InMux
    port map (
            O => \N__23673\,
            I => \N__23646\
        );

    \I__5525\ : InMux
    port map (
            O => \N__23670\,
            I => \N__23646\
        );

    \I__5524\ : InMux
    port map (
            O => \N__23669\,
            I => \N__23646\
        );

    \I__5523\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23646\
        );

    \I__5522\ : Span4Mux_h
    port map (
            O => \N__23663\,
            I => \N__23643\
        );

    \I__5521\ : InMux
    port map (
            O => \N__23662\,
            I => \N__23638\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__23655\,
            I => \N__23635\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23646\,
            I => \N__23630\
        );

    \I__5518\ : IoSpan4Mux
    port map (
            O => \N__23643\,
            I => \N__23630\
        );

    \I__5517\ : InMux
    port map (
            O => \N__23642\,
            I => \N__23625\
        );

    \I__5516\ : InMux
    port map (
            O => \N__23641\,
            I => \N__23625\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__23638\,
            I => \L3_tx_data_rdy\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__23635\,
            I => \L3_tx_data_rdy\
        );

    \I__5513\ : Odrv4
    port map (
            O => \N__23630\,
            I => \L3_tx_data_rdy\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__23625\,
            I => \L3_tx_data_rdy\
        );

    \I__5511\ : InMux
    port map (
            O => \N__23616\,
            I => \N__23613\
        );

    \I__5510\ : LocalMux
    port map (
            O => \N__23613\,
            I => \N__23610\
        );

    \I__5509\ : Span4Mux_s1_h
    port map (
            O => \N__23610\,
            I => \N__23600\
        );

    \I__5508\ : InMux
    port map (
            O => \N__23609\,
            I => \N__23593\
        );

    \I__5507\ : InMux
    port map (
            O => \N__23608\,
            I => \N__23593\
        );

    \I__5506\ : InMux
    port map (
            O => \N__23607\,
            I => \N__23593\
        );

    \I__5505\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23581\
        );

    \I__5504\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23581\
        );

    \I__5503\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23581\
        );

    \I__5502\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23581\
        );

    \I__5501\ : Span4Mux_h
    port map (
            O => \N__23600\,
            I => \N__23575\
        );

    \I__5500\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23572\
        );

    \I__5499\ : InMux
    port map (
            O => \N__23592\,
            I => \N__23565\
        );

    \I__5498\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23565\
        );

    \I__5497\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23565\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__23581\,
            I => \N__23562\
        );

    \I__5495\ : InMux
    port map (
            O => \N__23580\,
            I => \N__23555\
        );

    \I__5494\ : InMux
    port map (
            O => \N__23579\,
            I => \N__23555\
        );

    \I__5493\ : InMux
    port map (
            O => \N__23578\,
            I => \N__23555\
        );

    \I__5492\ : Odrv4
    port map (
            O => \N__23575\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__5491\ : Odrv4
    port map (
            O => \N__23572\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__23565\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__5489\ : Odrv4
    port map (
            O => \N__23562\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__23555\,
            I => \uu2.un1_w_user_cr_0\
        );

    \I__5487\ : CascadeMux
    port map (
            O => \N__23544\,
            I => \N__23540\
        );

    \I__5486\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23537\
        );

    \I__5485\ : InMux
    port map (
            O => \N__23540\,
            I => \N__23534\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__23537\,
            I => \N__23530\
        );

    \I__5483\ : LocalMux
    port map (
            O => \N__23534\,
            I => \N__23527\
        );

    \I__5482\ : InMux
    port map (
            O => \N__23533\,
            I => \N__23524\
        );

    \I__5481\ : Span4Mux_s1_v
    port map (
            O => \N__23530\,
            I => \N__23521\
        );

    \I__5480\ : Span12Mux_s1_h
    port map (
            O => \N__23527\,
            I => \N__23518\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__23524\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__5478\ : Odrv4
    port map (
            O => \N__23521\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__5477\ : Odrv12
    port map (
            O => \N__23518\,
            I => \uu2.w_addr_userZ0Z_8\
        );

    \I__5476\ : CascadeMux
    port map (
            O => \N__23511\,
            I => \N__23508\
        );

    \I__5475\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23505\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__23505\,
            I => \N__23502\
        );

    \I__5473\ : Span4Mux_s1_v
    port map (
            O => \N__23502\,
            I => \N__23499\
        );

    \I__5472\ : Span4Mux_h
    port map (
            O => \N__23499\,
            I => \N__23496\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__23496\,
            I => \N__23493\
        );

    \I__5470\ : Odrv4
    port map (
            O => \N__23493\,
            I => \uu2.mem0.w_addr_8\
        );

    \I__5469\ : InMux
    port map (
            O => \N__23490\,
            I => \N__23482\
        );

    \I__5468\ : InMux
    port map (
            O => \N__23489\,
            I => \N__23475\
        );

    \I__5467\ : InMux
    port map (
            O => \N__23488\,
            I => \N__23475\
        );

    \I__5466\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23475\
        );

    \I__5465\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23468\
        );

    \I__5464\ : CascadeMux
    port map (
            O => \N__23485\,
            I => \N__23465\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__23482\,
            I => \N__23457\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23457\
        );

    \I__5461\ : InMux
    port map (
            O => \N__23474\,
            I => \N__23450\
        );

    \I__5460\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23450\
        );

    \I__5459\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23450\
        );

    \I__5458\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23447\
        );

    \I__5457\ : LocalMux
    port map (
            O => \N__23468\,
            I => \N__23444\
        );

    \I__5456\ : InMux
    port map (
            O => \N__23465\,
            I => \N__23435\
        );

    \I__5455\ : InMux
    port map (
            O => \N__23464\,
            I => \N__23435\
        );

    \I__5454\ : InMux
    port map (
            O => \N__23463\,
            I => \N__23435\
        );

    \I__5453\ : InMux
    port map (
            O => \N__23462\,
            I => \N__23435\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__23457\,
            I => \N__23432\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__23450\,
            I => \N__23429\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__23447\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__5449\ : Odrv12
    port map (
            O => \N__23444\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__23435\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__5447\ : Odrv4
    port map (
            O => \N__23432\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__23429\,
            I => \uu2.w_addr_displayingZ0Z_1\
        );

    \I__5445\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23414\
        );

    \I__5444\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23411\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23408\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__23411\,
            I => \N__23405\
        );

    \I__5441\ : Span4Mux_s1_v
    port map (
            O => \N__23408\,
            I => \N__23397\
        );

    \I__5440\ : Span4Mux_s2_h
    port map (
            O => \N__23405\,
            I => \N__23397\
        );

    \I__5439\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23390\
        );

    \I__5438\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23390\
        );

    \I__5437\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23390\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__23397\,
            I => \uu2.N_75_mux\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__23390\,
            I => \uu2.N_75_mux\
        );

    \I__5434\ : CascadeMux
    port map (
            O => \N__23385\,
            I => \N__23382\
        );

    \I__5433\ : InMux
    port map (
            O => \N__23382\,
            I => \N__23377\
        );

    \I__5432\ : InMux
    port map (
            O => \N__23381\,
            I => \N__23374\
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__23380\,
            I => \N__23369\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23366\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__23374\,
            I => \N__23363\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__23373\,
            I => \N__23359\
        );

    \I__5427\ : InMux
    port map (
            O => \N__23372\,
            I => \N__23354\
        );

    \I__5426\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23354\
        );

    \I__5425\ : Span4Mux_h
    port map (
            O => \N__23366\,
            I => \N__23349\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__23363\,
            I => \N__23349\
        );

    \I__5423\ : InMux
    port map (
            O => \N__23362\,
            I => \N__23344\
        );

    \I__5422\ : InMux
    port map (
            O => \N__23359\,
            I => \N__23344\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23335\
        );

    \I__5420\ : IoSpan4Mux
    port map (
            O => \N__23349\,
            I => \N__23335\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__23344\,
            I => \N__23335\
        );

    \I__5418\ : CascadeMux
    port map (
            O => \N__23343\,
            I => \N__23331\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__23342\,
            I => \N__23324\
        );

    \I__5416\ : Sp12to4
    port map (
            O => \N__23335\,
            I => \N__23321\
        );

    \I__5415\ : InMux
    port map (
            O => \N__23334\,
            I => \N__23310\
        );

    \I__5414\ : InMux
    port map (
            O => \N__23331\,
            I => \N__23310\
        );

    \I__5413\ : InMux
    port map (
            O => \N__23330\,
            I => \N__23310\
        );

    \I__5412\ : InMux
    port map (
            O => \N__23329\,
            I => \N__23310\
        );

    \I__5411\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23310\
        );

    \I__5410\ : InMux
    port map (
            O => \N__23327\,
            I => \N__23305\
        );

    \I__5409\ : InMux
    port map (
            O => \N__23324\,
            I => \N__23305\
        );

    \I__5408\ : Span12Mux_s1_v
    port map (
            O => \N__23321\,
            I => \N__23300\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__23310\,
            I => \N__23300\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__23305\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__5405\ : Odrv12
    port map (
            O => \N__23300\,
            I => \uu2.w_addr_displayingZ0Z_0\
        );

    \I__5404\ : InMux
    port map (
            O => \N__23295\,
            I => \N__23292\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__23292\,
            I => \N__23286\
        );

    \I__5402\ : InMux
    port map (
            O => \N__23291\,
            I => \N__23279\
        );

    \I__5401\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23279\
        );

    \I__5400\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23279\
        );

    \I__5399\ : Span4Mux_s2_h
    port map (
            O => \N__23286\,
            I => \N__23274\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23271\
        );

    \I__5397\ : InMux
    port map (
            O => \N__23278\,
            I => \N__23266\
        );

    \I__5396\ : InMux
    port map (
            O => \N__23277\,
            I => \N__23266\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__23274\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__5394\ : Odrv4
    port map (
            O => \N__23271\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__23266\,
            I => \uu2.w_addr_displayingZ0Z_5\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__23259\,
            I => \uu2.N_14_i_cascade_\
        );

    \I__5391\ : CascadeMux
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__5390\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23238\
        );

    \I__5389\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23238\
        );

    \I__5388\ : InMux
    port map (
            O => \N__23251\,
            I => \N__23238\
        );

    \I__5387\ : InMux
    port map (
            O => \N__23250\,
            I => \N__23238\
        );

    \I__5386\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23238\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__23235\,
            I => \N__23232\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__23232\,
            I => \uu2.N_15_i\
        );

    \I__5382\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23226\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23223\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__23223\,
            I => \Lab_UT.dictrl.state_ret_12and_0_ns_sn\
        );

    \I__5379\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23217\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__23217\,
            I => \N__23214\
        );

    \I__5377\ : Odrv12
    port map (
            O => \N__23214\,
            I => \Lab_UT.dictrl.state_ret_12and_0_ns_rn_0\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__23211\,
            I => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\
        );

    \I__5375\ : InMux
    port map (
            O => \N__23208\,
            I => \N__23205\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__23205\,
            I => \N__23199\
        );

    \I__5373\ : InMux
    port map (
            O => \N__23204\,
            I => \N__23192\
        );

    \I__5372\ : InMux
    port map (
            O => \N__23203\,
            I => \N__23192\
        );

    \I__5371\ : InMux
    port map (
            O => \N__23202\,
            I => \N__23192\
        );

    \I__5370\ : Span4Mux_s3_h
    port map (
            O => \N__23199\,
            I => \N__23188\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__23192\,
            I => \N__23185\
        );

    \I__5368\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23182\
        );

    \I__5367\ : Odrv4
    port map (
            O => \N__23188\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__5366\ : Odrv12
    port map (
            O => \N__23185\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__23182\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0\
        );

    \I__5364\ : CascadeMux
    port map (
            O => \N__23175\,
            I => \Lab_UT.dictrl.g2_0_cascade_\
        );

    \I__5363\ : InMux
    port map (
            O => \N__23172\,
            I => \N__23169\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__23169\,
            I => \Lab_UT.dictrl.next_state_2_0_1\
        );

    \I__5361\ : CascadeMux
    port map (
            O => \N__23166\,
            I => \N__23156\
        );

    \I__5360\ : CascadeMux
    port map (
            O => \N__23165\,
            I => \N__23149\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__23164\,
            I => \N__23145\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__23163\,
            I => \N__23142\
        );

    \I__5357\ : CascadeMux
    port map (
            O => \N__23162\,
            I => \N__23139\
        );

    \I__5356\ : CascadeMux
    port map (
            O => \N__23161\,
            I => \N__23134\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__23160\,
            I => \N__23129\
        );

    \I__5354\ : InMux
    port map (
            O => \N__23159\,
            I => \N__23124\
        );

    \I__5353\ : InMux
    port map (
            O => \N__23156\,
            I => \N__23124\
        );

    \I__5352\ : CascadeMux
    port map (
            O => \N__23155\,
            I => \N__23120\
        );

    \I__5351\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23104\
        );

    \I__5350\ : InMux
    port map (
            O => \N__23153\,
            I => \N__23104\
        );

    \I__5349\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23104\
        );

    \I__5348\ : InMux
    port map (
            O => \N__23149\,
            I => \N__23104\
        );

    \I__5347\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23104\
        );

    \I__5346\ : InMux
    port map (
            O => \N__23145\,
            I => \N__23104\
        );

    \I__5345\ : InMux
    port map (
            O => \N__23142\,
            I => \N__23104\
        );

    \I__5344\ : InMux
    port map (
            O => \N__23139\,
            I => \N__23101\
        );

    \I__5343\ : InMux
    port map (
            O => \N__23138\,
            I => \N__23098\
        );

    \I__5342\ : InMux
    port map (
            O => \N__23137\,
            I => \N__23095\
        );

    \I__5341\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23090\
        );

    \I__5340\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23090\
        );

    \I__5339\ : InMux
    port map (
            O => \N__23132\,
            I => \N__23085\
        );

    \I__5338\ : InMux
    port map (
            O => \N__23129\,
            I => \N__23085\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__23124\,
            I => \N__23079\
        );

    \I__5336\ : InMux
    port map (
            O => \N__23123\,
            I => \N__23074\
        );

    \I__5335\ : InMux
    port map (
            O => \N__23120\,
            I => \N__23074\
        );

    \I__5334\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23071\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__23104\,
            I => \N__23066\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__23101\,
            I => \N__23066\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__23098\,
            I => \N__23063\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__23095\,
            I => \N__23060\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__23090\,
            I => \N__23055\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__23085\,
            I => \N__23055\
        );

    \I__5327\ : InMux
    port map (
            O => \N__23084\,
            I => \N__23052\
        );

    \I__5326\ : InMux
    port map (
            O => \N__23083\,
            I => \N__23049\
        );

    \I__5325\ : InMux
    port map (
            O => \N__23082\,
            I => \N__23046\
        );

    \I__5324\ : Span4Mux_s2_v
    port map (
            O => \N__23079\,
            I => \N__23041\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__23074\,
            I => \N__23041\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23036\
        );

    \I__5321\ : Span4Mux_h
    port map (
            O => \N__23066\,
            I => \N__23036\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__23063\,
            I => \N__23029\
        );

    \I__5319\ : Span4Mux_v
    port map (
            O => \N__23060\,
            I => \N__23029\
        );

    \I__5318\ : Span4Mux_v
    port map (
            O => \N__23055\,
            I => \N__23029\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23026\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__23049\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__23046\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5314\ : Odrv4
    port map (
            O => \N__23041\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5313\ : Odrv4
    port map (
            O => \N__23036\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5312\ : Odrv4
    port map (
            O => \N__23029\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5311\ : Odrv12
    port map (
            O => \N__23026\,
            I => \Lab_UT.dictrl.stateZ0Z_1\
        );

    \I__5310\ : InMux
    port map (
            O => \N__23013\,
            I => \N__23010\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__23010\,
            I => \N__23007\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__23007\,
            I => \Lab_UT.dictrl.N_1460_0\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__23004\,
            I => \Lab_UT.dictrl.g2_cascade_\
        );

    \I__5306\ : InMux
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__22998\,
            I => \N__22995\
        );

    \I__5304\ : Odrv4
    port map (
            O => \N__22995\,
            I => \Lab_UT.dictrl.next_state_0_1\
        );

    \I__5303\ : InMux
    port map (
            O => \N__22992\,
            I => \N__22989\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22989\,
            I => \N__22986\
        );

    \I__5301\ : Odrv12
    port map (
            O => \N__22986\,
            I => \Lab_UT.dictrl.N_40_3\
        );

    \I__5300\ : CascadeMux
    port map (
            O => \N__22983\,
            I => \Lab_UT.dictrl.N_1105_1_cascade_\
        );

    \I__5299\ : InMux
    port map (
            O => \N__22980\,
            I => \N__22974\
        );

    \I__5298\ : InMux
    port map (
            O => \N__22979\,
            I => \N__22969\
        );

    \I__5297\ : InMux
    port map (
            O => \N__22978\,
            I => \N__22963\
        );

    \I__5296\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22960\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__22974\,
            I => \N__22957\
        );

    \I__5294\ : InMux
    port map (
            O => \N__22973\,
            I => \N__22952\
        );

    \I__5293\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22952\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22949\
        );

    \I__5291\ : InMux
    port map (
            O => \N__22968\,
            I => \N__22940\
        );

    \I__5290\ : InMux
    port map (
            O => \N__22967\,
            I => \N__22937\
        );

    \I__5289\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22934\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22963\,
            I => \N__22931\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__22960\,
            I => \N__22928\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__22957\,
            I => \N__22921\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__22952\,
            I => \N__22921\
        );

    \I__5284\ : Span4Mux_v
    port map (
            O => \N__22949\,
            I => \N__22921\
        );

    \I__5283\ : InMux
    port map (
            O => \N__22948\,
            I => \N__22914\
        );

    \I__5282\ : InMux
    port map (
            O => \N__22947\,
            I => \N__22914\
        );

    \I__5281\ : InMux
    port map (
            O => \N__22946\,
            I => \N__22914\
        );

    \I__5280\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22907\
        );

    \I__5279\ : InMux
    port map (
            O => \N__22944\,
            I => \N__22907\
        );

    \I__5278\ : InMux
    port map (
            O => \N__22943\,
            I => \N__22907\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__22940\,
            I => \N__22904\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__22937\,
            I => \N__22899\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__22934\,
            I => \N__22899\
        );

    \I__5274\ : Span4Mux_s3_v
    port map (
            O => \N__22931\,
            I => \N__22894\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__22928\,
            I => \N__22894\
        );

    \I__5272\ : Span4Mux_h
    port map (
            O => \N__22921\,
            I => \N__22889\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22889\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__22907\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__5269\ : Odrv4
    port map (
            O => \N__22904\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__5268\ : Odrv12
    port map (
            O => \N__22899\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__5267\ : Odrv4
    port map (
            O => \N__22894\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__5266\ : Odrv4
    port map (
            O => \N__22889\,
            I => \Lab_UT.dictrl.state_i_3_2\
        );

    \I__5265\ : InMux
    port map (
            O => \N__22878\,
            I => \N__22875\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22872\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__22872\,
            I => \N__22869\
        );

    \I__5262\ : Odrv4
    port map (
            O => \N__22869\,
            I => \Lab_UT.dictrl.N_79_0\
        );

    \I__5261\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__5260\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__22860\,
            I => \N__22857\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__22857\,
            I => \Lab_UT.dictrl.N_40_5\
        );

    \I__5257\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22851\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__22851\,
            I => \N__22848\
        );

    \I__5255\ : Odrv4
    port map (
            O => \N__22848\,
            I => \Lab_UT.dictrl.g1_2\
        );

    \I__5254\ : InMux
    port map (
            O => \N__22845\,
            I => \N__22842\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__22842\,
            I => \N__22839\
        );

    \I__5252\ : Span4Mux_s2_h
    port map (
            O => \N__22839\,
            I => \N__22836\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__22836\,
            I => \Lab_UT.dictrl.N_40_2\
        );

    \I__5250\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__22830\,
            I => \N__22827\
        );

    \I__5248\ : Odrv4
    port map (
            O => \N__22827\,
            I => \Lab_UT.dictrl.g1_0\
        );

    \I__5247\ : InMux
    port map (
            O => \N__22824\,
            I => \N__22809\
        );

    \I__5246\ : InMux
    port map (
            O => \N__22823\,
            I => \N__22802\
        );

    \I__5245\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22802\
        );

    \I__5244\ : InMux
    port map (
            O => \N__22821\,
            I => \N__22802\
        );

    \I__5243\ : CascadeMux
    port map (
            O => \N__22820\,
            I => \N__22798\
        );

    \I__5242\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22795\
        );

    \I__5241\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22792\
        );

    \I__5240\ : InMux
    port map (
            O => \N__22817\,
            I => \N__22781\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22781\
        );

    \I__5238\ : InMux
    port map (
            O => \N__22815\,
            I => \N__22781\
        );

    \I__5237\ : InMux
    port map (
            O => \N__22814\,
            I => \N__22781\
        );

    \I__5236\ : InMux
    port map (
            O => \N__22813\,
            I => \N__22781\
        );

    \I__5235\ : InMux
    port map (
            O => \N__22812\,
            I => \N__22778\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__22809\,
            I => \N__22770\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__22802\,
            I => \N__22770\
        );

    \I__5232\ : InMux
    port map (
            O => \N__22801\,
            I => \N__22767\
        );

    \I__5231\ : InMux
    port map (
            O => \N__22798\,
            I => \N__22762\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22795\,
            I => \N__22759\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__22792\,
            I => \N__22756\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__22781\,
            I => \N__22751\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__22778\,
            I => \N__22751\
        );

    \I__5226\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22745\
        );

    \I__5225\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22745\
        );

    \I__5224\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22742\
        );

    \I__5223\ : Sp12to4
    port map (
            O => \N__22770\,
            I => \N__22737\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__22767\,
            I => \N__22737\
        );

    \I__5221\ : InMux
    port map (
            O => \N__22766\,
            I => \N__22734\
        );

    \I__5220\ : InMux
    port map (
            O => \N__22765\,
            I => \N__22731\
        );

    \I__5219\ : LocalMux
    port map (
            O => \N__22762\,
            I => \N__22726\
        );

    \I__5218\ : Span4Mux_s3_v
    port map (
            O => \N__22759\,
            I => \N__22726\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__22756\,
            I => \N__22721\
        );

    \I__5216\ : Span4Mux_s2_h
    port map (
            O => \N__22751\,
            I => \N__22721\
        );

    \I__5215\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22718\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__22745\,
            I => \N__22713\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__22742\,
            I => \N__22713\
        );

    \I__5212\ : Span12Mux_s7_v
    port map (
            O => \N__22737\,
            I => \N__22706\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__22734\,
            I => \N__22706\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__22731\,
            I => \N__22706\
        );

    \I__5209\ : Span4Mux_v
    port map (
            O => \N__22726\,
            I => \N__22703\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__22721\,
            I => \N__22700\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__22718\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5206\ : Odrv12
    port map (
            O => \N__22713\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5205\ : Odrv12
    port map (
            O => \N__22706\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5204\ : Odrv4
    port map (
            O => \N__22703\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5203\ : Odrv4
    port map (
            O => \N__22700\,
            I => \Lab_UT.dictrl.stateZ0Z_2\
        );

    \I__5202\ : InMux
    port map (
            O => \N__22689\,
            I => \N__22686\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__22686\,
            I => \N__22683\
        );

    \I__5200\ : Span4Mux_s2_h
    port map (
            O => \N__22683\,
            I => \N__22680\
        );

    \I__5199\ : Span4Mux_v
    port map (
            O => \N__22680\,
            I => \N__22677\
        );

    \I__5198\ : Odrv4
    port map (
            O => \N__22677\,
            I => \Lab_UT.dictrl.N_1460_4\
        );

    \I__5197\ : CascadeMux
    port map (
            O => \N__22674\,
            I => \N__22671\
        );

    \I__5196\ : InMux
    port map (
            O => \N__22671\,
            I => \N__22668\
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__22668\,
            I => \N__22665\
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__22665\,
            I => \Lab_UT.dictrl.g2_4\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__22662\,
            I => \Lab_UT.dictrl.next_state_4_1_cascade_\
        );

    \I__5192\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22656\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22653\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__22653\,
            I => \Lab_UT.didp.ceZ0Z_0\
        );

    \I__5189\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22647\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__22647\,
            I => \Lab_UT.LdSones_i_4\
        );

    \I__5187\ : InMux
    port map (
            O => \N__22644\,
            I => \N__22638\
        );

    \I__5186\ : InMux
    port map (
            O => \N__22643\,
            I => \N__22635\
        );

    \I__5185\ : InMux
    port map (
            O => \N__22642\,
            I => \N__22630\
        );

    \I__5184\ : InMux
    port map (
            O => \N__22641\,
            I => \N__22630\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__22638\,
            I => \N__22627\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__22635\,
            I => \N__22624\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__22630\,
            I => \N__22621\
        );

    \I__5180\ : Span4Mux_v
    port map (
            O => \N__22627\,
            I => \N__22618\
        );

    \I__5179\ : Span4Mux_h
    port map (
            O => \N__22624\,
            I => \N__22615\
        );

    \I__5178\ : Span4Mux_h
    port map (
            O => \N__22621\,
            I => \N__22612\
        );

    \I__5177\ : Odrv4
    port map (
            O => \N__22618\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__5176\ : Odrv4
    port map (
            O => \N__22615\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__5175\ : Odrv4
    port map (
            O => \N__22612\,
            I => \Lab_UT.didp.un1_dicLdSones_0\
        );

    \I__5174\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22600\
        );

    \I__5173\ : InMux
    port map (
            O => \N__22604\,
            I => \N__22595\
        );

    \I__5172\ : InMux
    port map (
            O => \N__22603\,
            I => \N__22595\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22600\,
            I => \N__22590\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__22595\,
            I => \N__22590\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__22590\,
            I => \N__22584\
        );

    \I__5168\ : InMux
    port map (
            O => \N__22589\,
            I => \N__22579\
        );

    \I__5167\ : InMux
    port map (
            O => \N__22588\,
            I => \N__22579\
        );

    \I__5166\ : InMux
    port map (
            O => \N__22587\,
            I => \N__22576\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__22584\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__22579\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__22576\,
            I => \Lab_UT.dictrl.next_stateZ0Z_2\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__22569\,
            I => \N__22564\
        );

    \I__5161\ : CascadeMux
    port map (
            O => \N__22568\,
            I => \N__22561\
        );

    \I__5160\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22553\
        );

    \I__5159\ : InMux
    port map (
            O => \N__22564\,
            I => \N__22553\
        );

    \I__5158\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22553\
        );

    \I__5157\ : CascadeMux
    port map (
            O => \N__22560\,
            I => \N__22547\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22544\
        );

    \I__5155\ : InMux
    port map (
            O => \N__22552\,
            I => \N__22541\
        );

    \I__5154\ : InMux
    port map (
            O => \N__22551\,
            I => \N__22538\
        );

    \I__5153\ : InMux
    port map (
            O => \N__22550\,
            I => \N__22533\
        );

    \I__5152\ : InMux
    port map (
            O => \N__22547\,
            I => \N__22533\
        );

    \I__5151\ : Odrv12
    port map (
            O => \N__22544\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22541\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__22538\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__22533\,
            I => \Lab_UT.dictrl.next_stateZ0Z_3\
        );

    \I__5147\ : CascadeMux
    port map (
            O => \N__22524\,
            I => \N__22518\
        );

    \I__5146\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22513\
        );

    \I__5145\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22513\
        );

    \I__5144\ : InMux
    port map (
            O => \N__22521\,
            I => \N__22508\
        );

    \I__5143\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22508\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__22513\,
            I => \N__22505\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__22508\,
            I => \N__22502\
        );

    \I__5140\ : Span4Mux_h
    port map (
            O => \N__22505\,
            I => \N__22499\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__22502\,
            I => \N__22496\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__22499\,
            I => \Lab_UT.LdSones\
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__22496\,
            I => \Lab_UT.LdSones\
        );

    \I__5136\ : CEMux
    port map (
            O => \N__22491\,
            I => \N__22473\
        );

    \I__5135\ : CEMux
    port map (
            O => \N__22490\,
            I => \N__22473\
        );

    \I__5134\ : CEMux
    port map (
            O => \N__22489\,
            I => \N__22473\
        );

    \I__5133\ : CEMux
    port map (
            O => \N__22488\,
            I => \N__22473\
        );

    \I__5132\ : CEMux
    port map (
            O => \N__22487\,
            I => \N__22473\
        );

    \I__5131\ : CEMux
    port map (
            O => \N__22486\,
            I => \N__22473\
        );

    \I__5130\ : GlobalMux
    port map (
            O => \N__22473\,
            I => \N__22470\
        );

    \I__5129\ : gio2CtrlBuf
    port map (
            O => \N__22470\,
            I => bu_rx_data_rdy_0_g
        );

    \I__5128\ : CascadeMux
    port map (
            O => \N__22467\,
            I => \N__22464\
        );

    \I__5127\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22459\
        );

    \I__5126\ : CascadeMux
    port map (
            O => \N__22463\,
            I => \N__22455\
        );

    \I__5125\ : CascadeMux
    port map (
            O => \N__22462\,
            I => \N__22452\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22449\
        );

    \I__5123\ : InMux
    port map (
            O => \N__22458\,
            I => \N__22442\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22442\
        );

    \I__5121\ : InMux
    port map (
            O => \N__22452\,
            I => \N__22442\
        );

    \I__5120\ : Span4Mux_v
    port map (
            O => \N__22449\,
            I => \N__22439\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22442\,
            I => \N__22436\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__22439\,
            I => \N__22433\
        );

    \I__5117\ : Span4Mux_h
    port map (
            O => \N__22436\,
            I => \N__22430\
        );

    \I__5116\ : Odrv4
    port map (
            O => \N__22433\,
            I => \Lab_UT.dictrl.g2_5\
        );

    \I__5115\ : Odrv4
    port map (
            O => \N__22430\,
            I => \Lab_UT.dictrl.g2_5\
        );

    \I__5114\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22422\
        );

    \I__5113\ : LocalMux
    port map (
            O => \N__22422\,
            I => \N__22415\
        );

    \I__5112\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22408\
        );

    \I__5111\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22408\
        );

    \I__5110\ : InMux
    port map (
            O => \N__22419\,
            I => \N__22408\
        );

    \I__5109\ : InMux
    port map (
            O => \N__22418\,
            I => \N__22405\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__22415\,
            I => \N__22402\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__22408\,
            I => \N__22399\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__22405\,
            I => \N__22396\
        );

    \I__5105\ : Span4Mux_v
    port map (
            O => \N__22402\,
            I => \N__22393\
        );

    \I__5104\ : Span4Mux_h
    port map (
            O => \N__22399\,
            I => \N__22388\
        );

    \I__5103\ : Span4Mux_s2_h
    port map (
            O => \N__22396\,
            I => \N__22388\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__22393\,
            I => \Lab_UT.dictrl.g1_3\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__22388\,
            I => \Lab_UT.dictrl.g1_3\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__22383\,
            I => \Lab_UT.dictrl.g2_5_cascade_\
        );

    \I__5099\ : InMux
    port map (
            O => \N__22380\,
            I => \N__22376\
        );

    \I__5098\ : CascadeMux
    port map (
            O => \N__22379\,
            I => \N__22373\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__22376\,
            I => \N__22367\
        );

    \I__5096\ : InMux
    port map (
            O => \N__22373\,
            I => \N__22360\
        );

    \I__5095\ : InMux
    port map (
            O => \N__22372\,
            I => \N__22360\
        );

    \I__5094\ : InMux
    port map (
            O => \N__22371\,
            I => \N__22360\
        );

    \I__5093\ : InMux
    port map (
            O => \N__22370\,
            I => \N__22357\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__22367\,
            I => \N__22354\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__22360\,
            I => \N__22351\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22348\
        );

    \I__5089\ : Span4Mux_v
    port map (
            O => \N__22354\,
            I => \N__22345\
        );

    \I__5088\ : Span4Mux_h
    port map (
            O => \N__22351\,
            I => \N__22340\
        );

    \I__5087\ : Span4Mux_s2_h
    port map (
            O => \N__22348\,
            I => \N__22340\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__22345\,
            I => \Lab_UT.dictrl.N_1460_5\
        );

    \I__5085\ : Odrv4
    port map (
            O => \N__22340\,
            I => \Lab_UT.dictrl.N_1460_5\
        );

    \I__5084\ : InMux
    port map (
            O => \N__22335\,
            I => \N__22329\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22334\,
            I => \N__22329\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__22326\,
            I => \N__22323\
        );

    \I__5080\ : Odrv4
    port map (
            O => \N__22323\,
            I => \Lab_UT.didp.ceZ0Z_3\
        );

    \I__5079\ : InMux
    port map (
            O => \N__22320\,
            I => \N__22316\
        );

    \I__5078\ : InMux
    port map (
            O => \N__22319\,
            I => \N__22313\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22308\
        );

    \I__5076\ : LocalMux
    port map (
            O => \N__22313\,
            I => \N__22308\
        );

    \I__5075\ : Odrv4
    port map (
            O => \N__22308\,
            I => \Lab_UT.didp.ceZ0Z_2\
        );

    \I__5074\ : CascadeMux
    port map (
            O => \N__22305\,
            I => \N__22299\
        );

    \I__5073\ : InMux
    port map (
            O => \N__22304\,
            I => \N__22287\
        );

    \I__5072\ : InMux
    port map (
            O => \N__22303\,
            I => \N__22287\
        );

    \I__5071\ : InMux
    port map (
            O => \N__22302\,
            I => \N__22287\
        );

    \I__5070\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22287\
        );

    \I__5069\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22287\
        );

    \I__5068\ : LocalMux
    port map (
            O => \N__22287\,
            I => \N__22284\
        );

    \I__5067\ : Odrv12
    port map (
            O => \N__22284\,
            I => \Lab_UT.didp.un24_ce_2\
        );

    \I__5066\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22276\
        );

    \I__5065\ : InMux
    port map (
            O => \N__22280\,
            I => \N__22273\
        );

    \I__5064\ : InMux
    port map (
            O => \N__22279\,
            I => \N__22270\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22263\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22260\
        );

    \I__5061\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22257\
        );

    \I__5060\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22254\
        );

    \I__5059\ : InMux
    port map (
            O => \N__22268\,
            I => \N__22251\
        );

    \I__5058\ : InMux
    port map (
            O => \N__22267\,
            I => \N__22248\
        );

    \I__5057\ : InMux
    port map (
            O => \N__22266\,
            I => \N__22245\
        );

    \I__5056\ : Span4Mux_h
    port map (
            O => \N__22263\,
            I => \N__22242\
        );

    \I__5055\ : Span4Mux_s3_h
    port map (
            O => \N__22260\,
            I => \N__22237\
        );

    \I__5054\ : Span4Mux_h
    port map (
            O => \N__22257\,
            I => \N__22237\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22234\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__22251\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__22248\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5050\ : LocalMux
    port map (
            O => \N__22245\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5049\ : Odrv4
    port map (
            O => \N__22242\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5048\ : Odrv4
    port map (
            O => \N__22237\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__22234\,
            I => \Lab_UT.di_Mtens_1\
        );

    \I__5046\ : CascadeMux
    port map (
            O => \N__22221\,
            I => \Lab_UT.didp.ce_12_3_cascade_\
        );

    \I__5045\ : InMux
    port map (
            O => \N__22218\,
            I => \N__22215\
        );

    \I__5044\ : LocalMux
    port map (
            O => \N__22215\,
            I => \N__22210\
        );

    \I__5043\ : CascadeMux
    port map (
            O => \N__22214\,
            I => \N__22205\
        );

    \I__5042\ : InMux
    port map (
            O => \N__22213\,
            I => \N__22202\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__22210\,
            I => \N__22199\
        );

    \I__5040\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22192\
        );

    \I__5039\ : InMux
    port map (
            O => \N__22208\,
            I => \N__22192\
        );

    \I__5038\ : InMux
    port map (
            O => \N__22205\,
            I => \N__22192\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__22202\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__5036\ : Odrv4
    port map (
            O => \N__22199\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__22192\,
            I => \Lab_UT.di_Mtens_3\
        );

    \I__5034\ : InMux
    port map (
            O => \N__22185\,
            I => \N__22179\
        );

    \I__5033\ : InMux
    port map (
            O => \N__22184\,
            I => \N__22179\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__22179\,
            I => \N__22174\
        );

    \I__5031\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22171\
        );

    \I__5030\ : InMux
    port map (
            O => \N__22177\,
            I => \N__22168\
        );

    \I__5029\ : Span4Mux_v
    port map (
            O => \N__22174\,
            I => \N__22165\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__22160\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__22160\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__22165\,
            I => \N__22157\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__22160\,
            I => \N__22154\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__22157\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__5023\ : Odrv4
    port map (
            O => \N__22154\,
            I => \Lab_UT.didp.resetZ0Z_3\
        );

    \I__5022\ : InMux
    port map (
            O => \N__22149\,
            I => \N__22130\
        );

    \I__5021\ : InMux
    port map (
            O => \N__22148\,
            I => \N__22130\
        );

    \I__5020\ : InMux
    port map (
            O => \N__22147\,
            I => \N__22130\
        );

    \I__5019\ : InMux
    port map (
            O => \N__22146\,
            I => \N__22130\
        );

    \I__5018\ : InMux
    port map (
            O => \N__22145\,
            I => \N__22130\
        );

    \I__5017\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22130\
        );

    \I__5016\ : InMux
    port map (
            O => \N__22143\,
            I => \N__22127\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__22130\,
            I => \N__22124\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__22127\,
            I => \N__22121\
        );

    \I__5013\ : Span4Mux_s2_h
    port map (
            O => \N__22124\,
            I => \N__22118\
        );

    \I__5012\ : Odrv12
    port map (
            O => \N__22121\,
            I => \Lab_UT.didp.un18_ce\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__22118\,
            I => \Lab_UT.didp.un18_ce\
        );

    \I__5010\ : CascadeMux
    port map (
            O => \N__22113\,
            I => \N__22105\
        );

    \I__5009\ : CascadeMux
    port map (
            O => \N__22112\,
            I => \N__22102\
        );

    \I__5008\ : CascadeMux
    port map (
            O => \N__22111\,
            I => \N__22099\
        );

    \I__5007\ : CascadeMux
    port map (
            O => \N__22110\,
            I => \N__22096\
        );

    \I__5006\ : CascadeMux
    port map (
            O => \N__22109\,
            I => \N__22091\
        );

    \I__5005\ : InMux
    port map (
            O => \N__22108\,
            I => \N__22084\
        );

    \I__5004\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22084\
        );

    \I__5003\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22071\
        );

    \I__5002\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22071\
        );

    \I__5001\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22071\
        );

    \I__5000\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22071\
        );

    \I__4999\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22071\
        );

    \I__4998\ : InMux
    port map (
            O => \N__22091\,
            I => \N__22071\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__22090\,
            I => \N__22066\
        );

    \I__4996\ : InMux
    port map (
            O => \N__22089\,
            I => \N__22062\
        );

    \I__4995\ : LocalMux
    port map (
            O => \N__22084\,
            I => \N__22059\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__22071\,
            I => \N__22056\
        );

    \I__4993\ : CascadeMux
    port map (
            O => \N__22070\,
            I => \N__22053\
        );

    \I__4992\ : InMux
    port map (
            O => \N__22069\,
            I => \N__22047\
        );

    \I__4991\ : InMux
    port map (
            O => \N__22066\,
            I => \N__22047\
        );

    \I__4990\ : CascadeMux
    port map (
            O => \N__22065\,
            I => \N__22044\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__22062\,
            I => \N__22041\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__22059\,
            I => \N__22036\
        );

    \I__4987\ : Span4Mux_s2_h
    port map (
            O => \N__22056\,
            I => \N__22036\
        );

    \I__4986\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22031\
        );

    \I__4985\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22028\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__22025\
        );

    \I__4983\ : InMux
    port map (
            O => \N__22044\,
            I => \N__22022\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__22041\,
            I => \N__22017\
        );

    \I__4981\ : Span4Mux_h
    port map (
            O => \N__22036\,
            I => \N__22017\
        );

    \I__4980\ : InMux
    port map (
            O => \N__22035\,
            I => \N__22012\
        );

    \I__4979\ : InMux
    port map (
            O => \N__22034\,
            I => \N__22012\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__22031\,
            I => \oneSecStrb\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__22028\,
            I => \oneSecStrb\
        );

    \I__4976\ : Odrv4
    port map (
            O => \N__22025\,
            I => \oneSecStrb\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__22022\,
            I => \oneSecStrb\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__22017\,
            I => \oneSecStrb\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__22012\,
            I => \oneSecStrb\
        );

    \I__4972\ : CascadeMux
    port map (
            O => \N__21999\,
            I => \N__21994\
        );

    \I__4971\ : InMux
    port map (
            O => \N__21998\,
            I => \N__21987\
        );

    \I__4970\ : InMux
    port map (
            O => \N__21997\,
            I => \N__21987\
        );

    \I__4969\ : InMux
    port map (
            O => \N__21994\,
            I => \N__21987\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21983\
        );

    \I__4967\ : InMux
    port map (
            O => \N__21986\,
            I => \N__21980\
        );

    \I__4966\ : Span12Mux_s7_v
    port map (
            O => \N__21983\,
            I => \N__21975\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21975\
        );

    \I__4964\ : Odrv12
    port map (
            O => \N__21975\,
            I => \Lab_UT.didp.resetZ0Z_0\
        );

    \I__4963\ : InMux
    port map (
            O => \N__21972\,
            I => \N__21967\
        );

    \I__4962\ : InMux
    port map (
            O => \N__21971\,
            I => \N__21964\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21970\,
            I => \N__21961\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21967\,
            I => \N__21956\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__21964\,
            I => \N__21953\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__21961\,
            I => \N__21949\
        );

    \I__4957\ : InMux
    port map (
            O => \N__21960\,
            I => \N__21943\
        );

    \I__4956\ : InMux
    port map (
            O => \N__21959\,
            I => \N__21943\
        );

    \I__4955\ : Span4Mux_v
    port map (
            O => \N__21956\,
            I => \N__21938\
        );

    \I__4954\ : Span4Mux_v
    port map (
            O => \N__21953\,
            I => \N__21938\
        );

    \I__4953\ : InMux
    port map (
            O => \N__21952\,
            I => \N__21935\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__21949\,
            I => \N__21932\
        );

    \I__4951\ : InMux
    port map (
            O => \N__21948\,
            I => \N__21929\
        );

    \I__4950\ : LocalMux
    port map (
            O => \N__21943\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4949\ : Odrv4
    port map (
            O => \N__21938\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__21935\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4947\ : Odrv4
    port map (
            O => \N__21932\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__21929\,
            I => \Lab_UT.di_Mtens_0\
        );

    \I__4945\ : InMux
    port map (
            O => \N__21918\,
            I => \N__21915\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__21915\,
            I => \N__21911\
        );

    \I__4943\ : InMux
    port map (
            O => \N__21914\,
            I => \N__21908\
        );

    \I__4942\ : Span4Mux_v
    port map (
            O => \N__21911\,
            I => \N__21899\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21908\,
            I => \N__21899\
        );

    \I__4940\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21896\
        );

    \I__4939\ : InMux
    port map (
            O => \N__21906\,
            I => \N__21889\
        );

    \I__4938\ : InMux
    port map (
            O => \N__21905\,
            I => \N__21889\
        );

    \I__4937\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21889\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__21899\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__21896\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4934\ : LocalMux
    port map (
            O => \N__21889\,
            I => \Lab_UT.di_Mtens_2\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21882\,
            I => \N__21879\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__21879\,
            I => \Lab_UT.didp.reset_12_1_3\
        );

    \I__4931\ : InMux
    port map (
            O => \N__21876\,
            I => \N__21873\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__21873\,
            I => \N__21870\
        );

    \I__4929\ : Span4Mux_s2_h
    port map (
            O => \N__21870\,
            I => \N__21867\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__21867\,
            I => \Lab_UT.didp.ceZ0Z_1\
        );

    \I__4927\ : InMux
    port map (
            O => \N__21864\,
            I => \N__21861\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__21861\,
            I => \N__21858\
        );

    \I__4925\ : Span4Mux_s3_h
    port map (
            O => \N__21858\,
            I => \N__21855\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__21855\,
            I => \Lab_UT.LdStens_i_4\
        );

    \I__4923\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21849\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__21849\,
            I => \N__21844\
        );

    \I__4921\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21839\
        );

    \I__4920\ : InMux
    port map (
            O => \N__21847\,
            I => \N__21839\
        );

    \I__4919\ : Span4Mux_v
    port map (
            O => \N__21844\,
            I => \N__21834\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__21839\,
            I => \N__21834\
        );

    \I__4917\ : Span4Mux_h
    port map (
            O => \N__21834\,
            I => \N__21831\
        );

    \I__4916\ : Odrv4
    port map (
            O => \N__21831\,
            I => \Lab_UT.di_AMones_3\
        );

    \I__4915\ : CEMux
    port map (
            O => \N__21828\,
            I => \N__21825\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__21825\,
            I => \N__21822\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__21822\,
            I => \N__21818\
        );

    \I__4912\ : CEMux
    port map (
            O => \N__21821\,
            I => \N__21815\
        );

    \I__4911\ : Span4Mux_s1_h
    port map (
            O => \N__21818\,
            I => \N__21810\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21810\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__21810\,
            I => \Lab_UT.didp.regrce3.LdAMones_0\
        );

    \I__4908\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21799\
        );

    \I__4907\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21796\
        );

    \I__4906\ : InMux
    port map (
            O => \N__21805\,
            I => \N__21793\
        );

    \I__4905\ : InMux
    port map (
            O => \N__21804\,
            I => \N__21790\
        );

    \I__4904\ : InMux
    port map (
            O => \N__21803\,
            I => \N__21787\
        );

    \I__4903\ : InMux
    port map (
            O => \N__21802\,
            I => \N__21783\
        );

    \I__4902\ : LocalMux
    port map (
            O => \N__21799\,
            I => \N__21780\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__21796\,
            I => \N__21776\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__21793\,
            I => \N__21771\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__21790\,
            I => \N__21767\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21764\
        );

    \I__4897\ : InMux
    port map (
            O => \N__21786\,
            I => \N__21761\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__21783\,
            I => \N__21756\
        );

    \I__4895\ : Span4Mux_s2_h
    port map (
            O => \N__21780\,
            I => \N__21756\
        );

    \I__4894\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21753\
        );

    \I__4893\ : Span4Mux_s2_h
    port map (
            O => \N__21776\,
            I => \N__21750\
        );

    \I__4892\ : InMux
    port map (
            O => \N__21775\,
            I => \N__21746\
        );

    \I__4891\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21743\
        );

    \I__4890\ : Span4Mux_h
    port map (
            O => \N__21771\,
            I => \N__21740\
        );

    \I__4889\ : InMux
    port map (
            O => \N__21770\,
            I => \N__21737\
        );

    \I__4888\ : Span4Mux_v
    port map (
            O => \N__21767\,
            I => \N__21730\
        );

    \I__4887\ : Span4Mux_v
    port map (
            O => \N__21764\,
            I => \N__21730\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21730\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__21756\,
            I => \N__21725\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__21753\,
            I => \N__21725\
        );

    \I__4883\ : Span4Mux_h
    port map (
            O => \N__21750\,
            I => \N__21722\
        );

    \I__4882\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21719\
        );

    \I__4881\ : LocalMux
    port map (
            O => \N__21746\,
            I => \N__21714\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__21743\,
            I => \N__21714\
        );

    \I__4879\ : Span4Mux_v
    port map (
            O => \N__21740\,
            I => \N__21711\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__21737\,
            I => \N__21704\
        );

    \I__4877\ : Span4Mux_h
    port map (
            O => \N__21730\,
            I => \N__21704\
        );

    \I__4876\ : Span4Mux_h
    port map (
            O => \N__21725\,
            I => \N__21701\
        );

    \I__4875\ : Span4Mux_v
    port map (
            O => \N__21722\,
            I => \N__21696\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__21719\,
            I => \N__21696\
        );

    \I__4873\ : Span12Mux_s10_h
    port map (
            O => \N__21714\,
            I => \N__21693\
        );

    \I__4872\ : Span4Mux_h
    port map (
            O => \N__21711\,
            I => \N__21690\
        );

    \I__4871\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21685\
        );

    \I__4870\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21685\
        );

    \I__4869\ : Span4Mux_h
    port map (
            O => \N__21704\,
            I => \N__21680\
        );

    \I__4868\ : Span4Mux_v
    port map (
            O => \N__21701\,
            I => \N__21680\
        );

    \I__4867\ : Span4Mux_h
    port map (
            O => \N__21696\,
            I => \N__21677\
        );

    \I__4866\ : Odrv12
    port map (
            O => \N__21693\,
            I => bu_rx_data_0
        );

    \I__4865\ : Odrv4
    port map (
            O => \N__21690\,
            I => bu_rx_data_0
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__21685\,
            I => bu_rx_data_0
        );

    \I__4863\ : Odrv4
    port map (
            O => \N__21680\,
            I => bu_rx_data_0
        );

    \I__4862\ : Odrv4
    port map (
            O => \N__21677\,
            I => bu_rx_data_0
        );

    \I__4861\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21663\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__21663\,
            I => \Lab_UT.didp.countrce3.q_5_0\
        );

    \I__4859\ : CascadeMux
    port map (
            O => \N__21660\,
            I => \Lab_UT.didp.un1_dicLdMones_0_cascade_\
        );

    \I__4858\ : InMux
    port map (
            O => \N__21657\,
            I => \N__21654\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__21654\,
            I => \Lab_UT.didp.countrce3.q_5_1\
        );

    \I__4856\ : InMux
    port map (
            O => \N__21651\,
            I => \N__21647\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21650\,
            I => \N__21644\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__21647\,
            I => \N__21641\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__21644\,
            I => \N__21637\
        );

    \I__4852\ : Span4Mux_v
    port map (
            O => \N__21641\,
            I => \N__21634\
        );

    \I__4851\ : InMux
    port map (
            O => \N__21640\,
            I => \N__21631\
        );

    \I__4850\ : Odrv12
    port map (
            O => \N__21637\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4849\ : Odrv4
    port map (
            O => \N__21634\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4848\ : LocalMux
    port map (
            O => \N__21631\,
            I => \Lab_UT.di_AMones_2\
        );

    \I__4847\ : InMux
    port map (
            O => \N__21624\,
            I => \N__21621\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__21621\,
            I => \N__21617\
        );

    \I__4845\ : InMux
    port map (
            O => \N__21620\,
            I => \N__21614\
        );

    \I__4844\ : Span4Mux_v
    port map (
            O => \N__21617\,
            I => \N__21610\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21607\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__21613\,
            I => \N__21604\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__21610\,
            I => \N__21601\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__21607\,
            I => \N__21598\
        );

    \I__4839\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21595\
        );

    \I__4838\ : Odrv4
    port map (
            O => \N__21601\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__4837\ : Odrv4
    port map (
            O => \N__21598\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__21595\,
            I => \Lab_UT.di_AMones_1\
        );

    \I__4835\ : InMux
    port map (
            O => \N__21588\,
            I => \N__21585\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__21585\,
            I => \N__21582\
        );

    \I__4833\ : Odrv4
    port map (
            O => \N__21582\,
            I => \Lab_UT.dispString.m49Z0Z_2\
        );

    \I__4832\ : CascadeMux
    port map (
            O => \N__21579\,
            I => \N__21575\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__21578\,
            I => \N__21572\
        );

    \I__4830\ : InMux
    port map (
            O => \N__21575\,
            I => \N__21562\
        );

    \I__4829\ : InMux
    port map (
            O => \N__21572\,
            I => \N__21562\
        );

    \I__4828\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21562\
        );

    \I__4827\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21557\
        );

    \I__4826\ : InMux
    port map (
            O => \N__21569\,
            I => \N__21557\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__21562\,
            I => \N__21554\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__21557\,
            I => \N__21551\
        );

    \I__4823\ : Span4Mux_s3_h
    port map (
            O => \N__21554\,
            I => \N__21546\
        );

    \I__4822\ : Span4Mux_s3_h
    port map (
            O => \N__21551\,
            I => \N__21543\
        );

    \I__4821\ : InMux
    port map (
            O => \N__21550\,
            I => \N__21538\
        );

    \I__4820\ : InMux
    port map (
            O => \N__21549\,
            I => \N__21538\
        );

    \I__4819\ : Odrv4
    port map (
            O => \N__21546\,
            I => \Lab_UT.sec2_1\
        );

    \I__4818\ : Odrv4
    port map (
            O => \N__21543\,
            I => \Lab_UT.sec2_1\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__21538\,
            I => \Lab_UT.sec2_1\
        );

    \I__4816\ : CascadeMux
    port map (
            O => \N__21531\,
            I => \N__21526\
        );

    \I__4815\ : InMux
    port map (
            O => \N__21530\,
            I => \N__21518\
        );

    \I__4814\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21518\
        );

    \I__4813\ : InMux
    port map (
            O => \N__21526\,
            I => \N__21518\
        );

    \I__4812\ : CascadeMux
    port map (
            O => \N__21525\,
            I => \N__21514\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21510\
        );

    \I__4810\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21505\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21505\
        );

    \I__4808\ : CascadeMux
    port map (
            O => \N__21513\,
            I => \N__21501\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__21510\,
            I => \N__21498\
        );

    \I__4806\ : LocalMux
    port map (
            O => \N__21505\,
            I => \N__21495\
        );

    \I__4805\ : InMux
    port map (
            O => \N__21504\,
            I => \N__21490\
        );

    \I__4804\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21490\
        );

    \I__4803\ : Span4Mux_s1_h
    port map (
            O => \N__21498\,
            I => \N__21485\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__21495\,
            I => \N__21485\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21482\
        );

    \I__4800\ : Odrv4
    port map (
            O => \N__21485\,
            I => \Lab_UT.sec2_3\
        );

    \I__4799\ : Odrv4
    port map (
            O => \N__21482\,
            I => \Lab_UT.sec2_3\
        );

    \I__4798\ : CascadeMux
    port map (
            O => \N__21477\,
            I => \N__21471\
        );

    \I__4797\ : InMux
    port map (
            O => \N__21476\,
            I => \N__21463\
        );

    \I__4796\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21463\
        );

    \I__4795\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21463\
        );

    \I__4794\ : InMux
    port map (
            O => \N__21471\,
            I => \N__21458\
        );

    \I__4793\ : InMux
    port map (
            O => \N__21470\,
            I => \N__21458\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__21463\,
            I => \N__21454\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__21458\,
            I => \N__21451\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__21457\,
            I => \N__21448\
        );

    \I__4789\ : Span4Mux_s2_h
    port map (
            O => \N__21454\,
            I => \N__21444\
        );

    \I__4788\ : Span4Mux_s2_h
    port map (
            O => \N__21451\,
            I => \N__21441\
        );

    \I__4787\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21436\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21436\
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__21444\,
            I => \Lab_UT.sec2_2\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__21441\,
            I => \Lab_UT.sec2_2\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__21436\,
            I => \Lab_UT.sec2_2\
        );

    \I__4782\ : InMux
    port map (
            O => \N__21429\,
            I => \N__21423\
        );

    \I__4781\ : InMux
    port map (
            O => \N__21428\,
            I => \N__21423\
        );

    \I__4780\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21417\
        );

    \I__4779\ : InMux
    port map (
            O => \N__21422\,
            I => \N__21410\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21421\,
            I => \N__21410\
        );

    \I__4777\ : InMux
    port map (
            O => \N__21420\,
            I => \N__21410\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__21417\,
            I => \N__21405\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__21410\,
            I => \N__21402\
        );

    \I__4774\ : InMux
    port map (
            O => \N__21409\,
            I => \N__21397\
        );

    \I__4773\ : InMux
    port map (
            O => \N__21408\,
            I => \N__21397\
        );

    \I__4772\ : Sp12to4
    port map (
            O => \N__21405\,
            I => \N__21394\
        );

    \I__4771\ : Span4Mux_s3_h
    port map (
            O => \N__21402\,
            I => \N__21389\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21389\
        );

    \I__4769\ : Odrv12
    port map (
            O => \N__21394\,
            I => \Lab_UT.sec2_0\
        );

    \I__4768\ : Odrv4
    port map (
            O => \N__21389\,
            I => \Lab_UT.sec2_0\
        );

    \I__4767\ : InMux
    port map (
            O => \N__21384\,
            I => \N__21381\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__21381\,
            I => \uu2.bitmapZ0Z_58\
        );

    \I__4765\ : CascadeMux
    port map (
            O => \N__21378\,
            I => \Lab_UT.didp.countrce2.q_5_0_cascade_\
        );

    \I__4764\ : InMux
    port map (
            O => \N__21375\,
            I => \N__21371\
        );

    \I__4763\ : InMux
    port map (
            O => \N__21374\,
            I => \N__21368\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__21371\,
            I => \N__21365\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__21368\,
            I => \N__21362\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__21365\,
            I => \N__21356\
        );

    \I__4759\ : Span4Mux_v
    port map (
            O => \N__21362\,
            I => \N__21356\
        );

    \I__4758\ : InMux
    port map (
            O => \N__21361\,
            I => \N__21353\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__21356\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__21353\,
            I => \Lab_UT.di_AStens_0\
        );

    \I__4755\ : CascadeMux
    port map (
            O => \N__21348\,
            I => \N__21337\
        );

    \I__4754\ : InMux
    port map (
            O => \N__21347\,
            I => \N__21333\
        );

    \I__4753\ : InMux
    port map (
            O => \N__21346\,
            I => \N__21328\
        );

    \I__4752\ : InMux
    port map (
            O => \N__21345\,
            I => \N__21328\
        );

    \I__4751\ : InMux
    port map (
            O => \N__21344\,
            I => \N__21321\
        );

    \I__4750\ : InMux
    port map (
            O => \N__21343\,
            I => \N__21321\
        );

    \I__4749\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21318\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21341\,
            I => \N__21309\
        );

    \I__4747\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21309\
        );

    \I__4746\ : InMux
    port map (
            O => \N__21337\,
            I => \N__21309\
        );

    \I__4745\ : InMux
    port map (
            O => \N__21336\,
            I => \N__21309\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__21333\,
            I => \N__21304\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21304\
        );

    \I__4742\ : InMux
    port map (
            O => \N__21327\,
            I => \N__21298\
        );

    \I__4741\ : InMux
    port map (
            O => \N__21326\,
            I => \N__21295\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__21321\,
            I => \N__21288\
        );

    \I__4739\ : LocalMux
    port map (
            O => \N__21318\,
            I => \N__21288\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21288\
        );

    \I__4737\ : Span4Mux_s3_h
    port map (
            O => \N__21304\,
            I => \N__21285\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21303\,
            I => \N__21282\
        );

    \I__4735\ : InMux
    port map (
            O => \N__21302\,
            I => \N__21277\
        );

    \I__4734\ : InMux
    port map (
            O => \N__21301\,
            I => \N__21277\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__21298\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4732\ : LocalMux
    port map (
            O => \N__21295\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__21288\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__21285\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4729\ : LocalMux
    port map (
            O => \N__21282\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__21277\,
            I => \Lab_UT.loadalarm_0\
        );

    \I__4727\ : InMux
    port map (
            O => \N__21264\,
            I => \N__21260\
        );

    \I__4726\ : InMux
    port map (
            O => \N__21263\,
            I => \N__21252\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__21260\,
            I => \N__21249\
        );

    \I__4724\ : InMux
    port map (
            O => \N__21259\,
            I => \N__21240\
        );

    \I__4723\ : InMux
    port map (
            O => \N__21258\,
            I => \N__21240\
        );

    \I__4722\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21240\
        );

    \I__4721\ : InMux
    port map (
            O => \N__21256\,
            I => \N__21240\
        );

    \I__4720\ : InMux
    port map (
            O => \N__21255\,
            I => \N__21237\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__21252\,
            I => \N__21232\
        );

    \I__4718\ : Span4Mux_s2_h
    port map (
            O => \N__21249\,
            I => \N__21232\
        );

    \I__4717\ : LocalMux
    port map (
            O => \N__21240\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__21237\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4715\ : Odrv4
    port map (
            O => \N__21232\,
            I => \Lab_UT.di_Sones_1\
        );

    \I__4714\ : InMux
    port map (
            O => \N__21225\,
            I => \N__21222\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__21222\,
            I => \N__21217\
        );

    \I__4712\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21212\
        );

    \I__4711\ : InMux
    port map (
            O => \N__21220\,
            I => \N__21212\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__21217\,
            I => \N__21209\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__21212\,
            I => \N__21206\
        );

    \I__4708\ : Span4Mux_h
    port map (
            O => \N__21209\,
            I => \N__21203\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__21206\,
            I => \N__21200\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__21203\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__21200\,
            I => \Lab_UT.di_AStens_1\
        );

    \I__4704\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21191\
        );

    \I__4703\ : InMux
    port map (
            O => \N__21194\,
            I => \N__21187\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21184\
        );

    \I__4701\ : InMux
    port map (
            O => \N__21190\,
            I => \N__21181\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__21187\,
            I => \N__21178\
        );

    \I__4699\ : Odrv4
    port map (
            O => \N__21184\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__21181\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4697\ : Odrv4
    port map (
            O => \N__21178\,
            I => \Lab_UT.di_ASones_1\
        );

    \I__4696\ : InMux
    port map (
            O => \N__21171\,
            I => \N__21168\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__21168\,
            I => \N__21165\
        );

    \I__4694\ : Span4Mux_h
    port map (
            O => \N__21165\,
            I => \N__21162\
        );

    \I__4693\ : Odrv4
    port map (
            O => \N__21162\,
            I => \Lab_UT.dispString.m49Z0Z_5\
        );

    \I__4692\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21156\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__21156\,
            I => \uu2.bitmapZ0Z_218\
        );

    \I__4690\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21150\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__21150\,
            I => \uu2.bitmapZ0Z_90\
        );

    \I__4688\ : InMux
    port map (
            O => \N__21147\,
            I => \N__21144\
        );

    \I__4687\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__21141\
        );

    \I__4686\ : Span4Mux_h
    port map (
            O => \N__21141\,
            I => \N__21138\
        );

    \I__4685\ : Odrv4
    port map (
            O => \N__21138\,
            I => \uu2.N_20\
        );

    \I__4684\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21128\
        );

    \I__4683\ : InMux
    port map (
            O => \N__21134\,
            I => \N__21121\
        );

    \I__4682\ : InMux
    port map (
            O => \N__21133\,
            I => \N__21121\
        );

    \I__4681\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21118\
        );

    \I__4680\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21115\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__21128\,
            I => \N__21112\
        );

    \I__4678\ : InMux
    port map (
            O => \N__21127\,
            I => \N__21109\
        );

    \I__4677\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21106\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__21103\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__21118\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__21115\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4673\ : Odrv4
    port map (
            O => \N__21112\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__21109\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__21106\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4670\ : Odrv4
    port map (
            O => \N__21103\,
            I => \uu2.w_addr_displaying_fastZ0Z_7\
        );

    \I__4669\ : CascadeMux
    port map (
            O => \N__21090\,
            I => \uu2.bitmap_RNIE7RKZ0Z_58_cascade_\
        );

    \I__4668\ : InMux
    port map (
            O => \N__21087\,
            I => \N__21084\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__21084\,
            I => \uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7\
        );

    \I__4666\ : InMux
    port map (
            O => \N__21081\,
            I => \N__21076\
        );

    \I__4665\ : InMux
    port map (
            O => \N__21080\,
            I => \N__21073\
        );

    \I__4664\ : InMux
    port map (
            O => \N__21079\,
            I => \N__21070\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__21076\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__4662\ : LocalMux
    port map (
            O => \N__21073\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__21070\,
            I => \uu2.bitmapZ0Z_314\
        );

    \I__4660\ : InMux
    port map (
            O => \N__21063\,
            I => \N__21060\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__21060\,
            I => \uu2.bitmap_RNI020QZ0Z_186\
        );

    \I__4658\ : InMux
    port map (
            O => \N__21057\,
            I => \N__21054\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__21054\,
            I => \uu2.bitmapZ0Z_186\
        );

    \I__4656\ : InMux
    port map (
            O => \N__21051\,
            I => \N__21044\
        );

    \I__4655\ : InMux
    port map (
            O => \N__21050\,
            I => \N__21044\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__21049\,
            I => \N__21041\
        );

    \I__4653\ : LocalMux
    port map (
            O => \N__21044\,
            I => \N__21038\
        );

    \I__4652\ : InMux
    port map (
            O => \N__21041\,
            I => \N__21034\
        );

    \I__4651\ : Span4Mux_h
    port map (
            O => \N__21038\,
            I => \N__21031\
        );

    \I__4650\ : InMux
    port map (
            O => \N__21037\,
            I => \N__21028\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__21034\,
            I => \N__21025\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__21031\,
            I => \N__21022\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__21028\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4646\ : Odrv12
    port map (
            O => \N__21025\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__21022\,
            I => \uu2.w_addr_userZ0Z_5\
        );

    \I__4644\ : InMux
    port map (
            O => \N__21015\,
            I => \N__21009\
        );

    \I__4643\ : InMux
    port map (
            O => \N__21014\,
            I => \N__21006\
        );

    \I__4642\ : InMux
    port map (
            O => \N__21013\,
            I => \N__21003\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__21012\,
            I => \N__21000\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__20996\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20991\
        );

    \I__4638\ : LocalMux
    port map (
            O => \N__21003\,
            I => \N__20991\
        );

    \I__4637\ : InMux
    port map (
            O => \N__21000\,
            I => \N__20986\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20999\,
            I => \N__20986\
        );

    \I__4635\ : Span4Mux_s0_v
    port map (
            O => \N__20996\,
            I => \N__20983\
        );

    \I__4634\ : Span12Mux_s10_h
    port map (
            O => \N__20991\,
            I => \N__20980\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20986\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__20983\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4631\ : Odrv12
    port map (
            O => \N__20980\,
            I => \uu2.w_addr_userZ0Z_4\
        );

    \I__4630\ : InMux
    port map (
            O => \N__20973\,
            I => \N__20964\
        );

    \I__4629\ : InMux
    port map (
            O => \N__20972\,
            I => \N__20964\
        );

    \I__4628\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20964\
        );

    \I__4627\ : LocalMux
    port map (
            O => \N__20964\,
            I => \N__20961\
        );

    \I__4626\ : Span4Mux_s1_h
    port map (
            O => \N__20961\,
            I => \N__20955\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20960\,
            I => \N__20948\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20959\,
            I => \N__20948\
        );

    \I__4623\ : InMux
    port map (
            O => \N__20958\,
            I => \N__20948\
        );

    \I__4622\ : Span4Mux_h
    port map (
            O => \N__20955\,
            I => \N__20944\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__20948\,
            I => \N__20941\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20947\,
            I => \N__20938\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__20944\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4618\ : Odrv4
    port map (
            O => \N__20941\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__20938\,
            I => \uu2.un28_w_addr_user_i\
        );

    \I__4616\ : InMux
    port map (
            O => \N__20931\,
            I => \N__20922\
        );

    \I__4615\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20922\
        );

    \I__4614\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20922\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20917\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20921\,
            I => \N__20912\
        );

    \I__4611\ : InMux
    port map (
            O => \N__20920\,
            I => \N__20912\
        );

    \I__4610\ : Odrv12
    port map (
            O => \N__20917\,
            I => \uu2.un404_ci\
        );

    \I__4609\ : LocalMux
    port map (
            O => \N__20912\,
            I => \uu2.un404_ci\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__20907\,
            I => \N__20904\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20904\,
            I => \N__20901\
        );

    \I__4606\ : LocalMux
    port map (
            O => \N__20901\,
            I => \N__20898\
        );

    \I__4605\ : Span4Mux_s1_v
    port map (
            O => \N__20898\,
            I => \N__20895\
        );

    \I__4604\ : Span4Mux_h
    port map (
            O => \N__20895\,
            I => \N__20891\
        );

    \I__4603\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20888\
        );

    \I__4602\ : Odrv4
    port map (
            O => \N__20891\,
            I => \uu2.un426_ci_3\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__20888\,
            I => \uu2.un426_ci_3\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20883\,
            I => \N__20876\
        );

    \I__4599\ : InMux
    port map (
            O => \N__20882\,
            I => \N__20876\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__20881\,
            I => \N__20873\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__20876\,
            I => \N__20868\
        );

    \I__4596\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20865\
        );

    \I__4595\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20862\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20871\,
            I => \N__20859\
        );

    \I__4593\ : Span12Mux_v
    port map (
            O => \N__20868\,
            I => \N__20854\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20865\,
            I => \N__20854\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20862\,
            I => \N__20851\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__20859\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__4589\ : Odrv12
    port map (
            O => \N__20854\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__4588\ : Odrv4
    port map (
            O => \N__20851\,
            I => \uu2.w_addr_userZ0Z_6\
        );

    \I__4587\ : SRMux
    port map (
            O => \N__20844\,
            I => \N__20839\
        );

    \I__4586\ : SRMux
    port map (
            O => \N__20843\,
            I => \N__20836\
        );

    \I__4585\ : SRMux
    port map (
            O => \N__20842\,
            I => \N__20833\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20830\
        );

    \I__4583\ : LocalMux
    port map (
            O => \N__20836\,
            I => \N__20827\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20833\,
            I => \N__20824\
        );

    \I__4581\ : Span12Mux_s2_v
    port map (
            O => \N__20830\,
            I => \N__20820\
        );

    \I__4580\ : Span4Mux_s2_v
    port map (
            O => \N__20827\,
            I => \N__20817\
        );

    \I__4579\ : Span4Mux_h
    port map (
            O => \N__20824\,
            I => \N__20814\
        );

    \I__4578\ : InMux
    port map (
            O => \N__20823\,
            I => \N__20811\
        );

    \I__4577\ : Odrv12
    port map (
            O => \N__20820\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__4576\ : Odrv4
    port map (
            O => \N__20817\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__4575\ : Odrv4
    port map (
            O => \N__20814\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20811\,
            I => \uu2.w_addr_user_RNI43E87Z0Z_2\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__20802\,
            I => \uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_\
        );

    \I__4572\ : InMux
    port map (
            O => \N__20799\,
            I => \N__20796\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__20796\,
            I => \N__20793\
        );

    \I__4570\ : Odrv12
    port map (
            O => \N__20793\,
            I => \uu2.N_397\
        );

    \I__4569\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20785\
        );

    \I__4568\ : InMux
    port map (
            O => \N__20789\,
            I => \N__20778\
        );

    \I__4567\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20778\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__20785\,
            I => \N__20775\
        );

    \I__4565\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20770\
        );

    \I__4564\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20770\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__20778\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__20775\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__20770\,
            I => \uu2.w_addr_displaying_fastZ0Z_1\
        );

    \I__4560\ : InMux
    port map (
            O => \N__20763\,
            I => \N__20745\
        );

    \I__4559\ : InMux
    port map (
            O => \N__20762\,
            I => \N__20745\
        );

    \I__4558\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20745\
        );

    \I__4557\ : InMux
    port map (
            O => \N__20760\,
            I => \N__20745\
        );

    \I__4556\ : InMux
    port map (
            O => \N__20759\,
            I => \N__20737\
        );

    \I__4555\ : InMux
    port map (
            O => \N__20758\,
            I => \N__20737\
        );

    \I__4554\ : InMux
    port map (
            O => \N__20757\,
            I => \N__20734\
        );

    \I__4553\ : InMux
    port map (
            O => \N__20756\,
            I => \N__20731\
        );

    \I__4552\ : InMux
    port map (
            O => \N__20755\,
            I => \N__20728\
        );

    \I__4551\ : InMux
    port map (
            O => \N__20754\,
            I => \N__20725\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__20745\,
            I => \N__20722\
        );

    \I__4549\ : InMux
    port map (
            O => \N__20744\,
            I => \N__20717\
        );

    \I__4548\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20717\
        );

    \I__4547\ : InMux
    port map (
            O => \N__20742\,
            I => \N__20714\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20711\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__20734\,
            I => \N__20706\
        );

    \I__4544\ : LocalMux
    port map (
            O => \N__20731\,
            I => \N__20706\
        );

    \I__4543\ : LocalMux
    port map (
            O => \N__20728\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__20725\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__20722\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__20717\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__20714\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4538\ : Odrv4
    port map (
            O => \N__20711\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4537\ : Odrv4
    port map (
            O => \N__20706\,
            I => \uu2.w_addr_displayingZ1Z_3\
        );

    \I__4536\ : InMux
    port map (
            O => \N__20691\,
            I => \N__20688\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__20688\,
            I => \uu2.bitmap_pmux_sn_N_11\
        );

    \I__4534\ : CascadeMux
    port map (
            O => \N__20685\,
            I => \N__20682\
        );

    \I__4533\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20679\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__20679\,
            I => \uu2.N_32\
        );

    \I__4531\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20669\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20675\,
            I => \N__20664\
        );

    \I__4529\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20664\
        );

    \I__4528\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20656\
        );

    \I__4527\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20656\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__20669\,
            I => \N__20653\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__20664\,
            I => \N__20650\
        );

    \I__4524\ : InMux
    port map (
            O => \N__20663\,
            I => \N__20643\
        );

    \I__4523\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20643\
        );

    \I__4522\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20643\
        );

    \I__4521\ : LocalMux
    port map (
            O => \N__20656\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__4520\ : Odrv4
    port map (
            O => \N__20653\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__4519\ : Odrv12
    port map (
            O => \N__20650\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20643\,
            I => \uu2.w_addr_displaying_fastZ0Z_3\
        );

    \I__4517\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20630\
        );

    \I__4516\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20625\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__20630\,
            I => \N__20622\
        );

    \I__4514\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20617\
        );

    \I__4513\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20617\
        );

    \I__4512\ : LocalMux
    port map (
            O => \N__20625\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__4511\ : Odrv4
    port map (
            O => \N__20622\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__20617\,
            I => \uu2.w_addr_displaying_fastZ0Z_2\
        );

    \I__4509\ : InMux
    port map (
            O => \N__20610\,
            I => \N__20607\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__20607\,
            I => \N__20604\
        );

    \I__4507\ : Odrv4
    port map (
            O => \N__20604\,
            I => \uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2\
        );

    \I__4506\ : CascadeMux
    port map (
            O => \N__20601\,
            I => \N__20598\
        );

    \I__4505\ : InMux
    port map (
            O => \N__20598\,
            I => \N__20586\
        );

    \I__4504\ : InMux
    port map (
            O => \N__20597\,
            I => \N__20586\
        );

    \I__4503\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20581\
        );

    \I__4502\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20581\
        );

    \I__4501\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20567\
        );

    \I__4500\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20567\
        );

    \I__4499\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20567\
        );

    \I__4498\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20567\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__20586\,
            I => \N__20562\
        );

    \I__4496\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20562\
        );

    \I__4495\ : InMux
    port map (
            O => \N__20580\,
            I => \N__20555\
        );

    \I__4494\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20555\
        );

    \I__4493\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20555\
        );

    \I__4492\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20552\
        );

    \I__4491\ : InMux
    port map (
            O => \N__20576\,
            I => \N__20549\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__20567\,
            I => \N__20546\
        );

    \I__4489\ : Span4Mux_v
    port map (
            O => \N__20562\,
            I => \N__20541\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__20555\,
            I => \N__20541\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__20552\,
            I => \Lab_UT.dictrl.m23_aZ0Z0\
        );

    \I__4486\ : LocalMux
    port map (
            O => \N__20549\,
            I => \Lab_UT.dictrl.m23_aZ0Z0\
        );

    \I__4485\ : Odrv12
    port map (
            O => \N__20546\,
            I => \Lab_UT.dictrl.m23_aZ0Z0\
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__20541\,
            I => \Lab_UT.dictrl.m23_aZ0Z0\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20532\,
            I => \N__20529\
        );

    \I__4482\ : LocalMux
    port map (
            O => \N__20529\,
            I => \Lab_UT.dictrl.N_40_7\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__20526\,
            I => \Lab_UT.dictrl.N_40_7_cascade_\
        );

    \I__4480\ : InMux
    port map (
            O => \N__20523\,
            I => \N__20520\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__20520\,
            I => \Lab_UT.dictrl.g2_1_5\
        );

    \I__4478\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \Lab_UT.dictrl.N_1462_5_cascade_\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20514\,
            I => \N__20511\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__20511\,
            I => \Lab_UT.dictrl.N_1102_5\
        );

    \I__4475\ : InMux
    port map (
            O => \N__20508\,
            I => \N__20505\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20499\
        );

    \I__4473\ : InMux
    port map (
            O => \N__20504\,
            I => \N__20494\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__20503\,
            I => \N__20490\
        );

    \I__4471\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20484\
        );

    \I__4470\ : Span4Mux_v
    port map (
            O => \N__20499\,
            I => \N__20481\
        );

    \I__4469\ : InMux
    port map (
            O => \N__20498\,
            I => \N__20476\
        );

    \I__4468\ : InMux
    port map (
            O => \N__20497\,
            I => \N__20476\
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__20494\,
            I => \N__20473\
        );

    \I__4466\ : InMux
    port map (
            O => \N__20493\,
            I => \N__20470\
        );

    \I__4465\ : InMux
    port map (
            O => \N__20490\,
            I => \N__20465\
        );

    \I__4464\ : InMux
    port map (
            O => \N__20489\,
            I => \N__20465\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__20488\,
            I => \N__20462\
        );

    \I__4462\ : InMux
    port map (
            O => \N__20487\,
            I => \N__20459\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__20484\,
            I => \N__20456\
        );

    \I__4460\ : Sp12to4
    port map (
            O => \N__20481\,
            I => \N__20453\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20450\
        );

    \I__4458\ : Span4Mux_h
    port map (
            O => \N__20473\,
            I => \N__20445\
        );

    \I__4457\ : LocalMux
    port map (
            O => \N__20470\,
            I => \N__20445\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__20465\,
            I => \N__20442\
        );

    \I__4455\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20439\
        );

    \I__4454\ : LocalMux
    port map (
            O => \N__20459\,
            I => \N__20436\
        );

    \I__4453\ : Span4Mux_v
    port map (
            O => \N__20456\,
            I => \N__20433\
        );

    \I__4452\ : Span12Mux_s8_h
    port map (
            O => \N__20453\,
            I => \N__20430\
        );

    \I__4451\ : Span4Mux_h
    port map (
            O => \N__20450\,
            I => \N__20423\
        );

    \I__4450\ : Span4Mux_h
    port map (
            O => \N__20445\,
            I => \N__20423\
        );

    \I__4449\ : Span4Mux_s3_h
    port map (
            O => \N__20442\,
            I => \N__20423\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20418\
        );

    \I__4447\ : Span4Mux_h
    port map (
            O => \N__20436\,
            I => \N__20418\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__20433\,
            I => bu_rx_data_0_rep1
        );

    \I__4445\ : Odrv12
    port map (
            O => \N__20430\,
            I => bu_rx_data_0_rep1
        );

    \I__4444\ : Odrv4
    port map (
            O => \N__20423\,
            I => bu_rx_data_0_rep1
        );

    \I__4443\ : Odrv4
    port map (
            O => \N__20418\,
            I => bu_rx_data_0_rep1
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__20409\,
            I => \N__20403\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20408\,
            I => \N__20399\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__20407\,
            I => \N__20396\
        );

    \I__4439\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20387\
        );

    \I__4438\ : InMux
    port map (
            O => \N__20403\,
            I => \N__20387\
        );

    \I__4437\ : InMux
    port map (
            O => \N__20402\,
            I => \N__20387\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20399\,
            I => \N__20384\
        );

    \I__4435\ : InMux
    port map (
            O => \N__20396\,
            I => \N__20379\
        );

    \I__4434\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20379\
        );

    \I__4433\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20376\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__20387\,
            I => \N__20372\
        );

    \I__4431\ : Span4Mux_s2_v
    port map (
            O => \N__20384\,
            I => \N__20367\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__20379\,
            I => \N__20367\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__20376\,
            I => \N__20364\
        );

    \I__4428\ : CascadeMux
    port map (
            O => \N__20375\,
            I => \N__20361\
        );

    \I__4427\ : Span4Mux_s2_v
    port map (
            O => \N__20372\,
            I => \N__20357\
        );

    \I__4426\ : Span4Mux_v
    port map (
            O => \N__20367\,
            I => \N__20354\
        );

    \I__4425\ : Span4Mux_s2_v
    port map (
            O => \N__20364\,
            I => \N__20351\
        );

    \I__4424\ : InMux
    port map (
            O => \N__20361\,
            I => \N__20348\
        );

    \I__4423\ : InMux
    port map (
            O => \N__20360\,
            I => \N__20345\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__20357\,
            I => \N__20342\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__20354\,
            I => \N__20337\
        );

    \I__4420\ : Span4Mux_v
    port map (
            O => \N__20351\,
            I => \N__20337\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__20348\,
            I => \N__20332\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__20345\,
            I => \N__20332\
        );

    \I__4417\ : Odrv4
    port map (
            O => \N__20342\,
            I => bu_rx_data_5_rep1
        );

    \I__4416\ : Odrv4
    port map (
            O => \N__20337\,
            I => bu_rx_data_5_rep1
        );

    \I__4415\ : Odrv12
    port map (
            O => \N__20332\,
            I => bu_rx_data_5_rep1
        );

    \I__4414\ : InMux
    port map (
            O => \N__20325\,
            I => \N__20311\
        );

    \I__4413\ : InMux
    port map (
            O => \N__20324\,
            I => \N__20311\
        );

    \I__4412\ : InMux
    port map (
            O => \N__20323\,
            I => \N__20311\
        );

    \I__4411\ : InMux
    port map (
            O => \N__20322\,
            I => \N__20301\
        );

    \I__4410\ : InMux
    port map (
            O => \N__20321\,
            I => \N__20301\
        );

    \I__4409\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20301\
        );

    \I__4408\ : InMux
    port map (
            O => \N__20319\,
            I => \N__20301\
        );

    \I__4407\ : InMux
    port map (
            O => \N__20318\,
            I => \N__20298\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20311\,
            I => \N__20292\
        );

    \I__4405\ : InMux
    port map (
            O => \N__20310\,
            I => \N__20289\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__20301\,
            I => \N__20284\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__20298\,
            I => \N__20284\
        );

    \I__4402\ : InMux
    port map (
            O => \N__20297\,
            I => \N__20279\
        );

    \I__4401\ : InMux
    port map (
            O => \N__20296\,
            I => \N__20274\
        );

    \I__4400\ : InMux
    port map (
            O => \N__20295\,
            I => \N__20274\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__20292\,
            I => \N__20269\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__20289\,
            I => \N__20269\
        );

    \I__4397\ : Span4Mux_s3_v
    port map (
            O => \N__20284\,
            I => \N__20264\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20283\,
            I => \N__20259\
        );

    \I__4395\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20259\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20256\
        );

    \I__4393\ : LocalMux
    port map (
            O => \N__20274\,
            I => \N__20251\
        );

    \I__4392\ : Span4Mux_h
    port map (
            O => \N__20269\,
            I => \N__20251\
        );

    \I__4391\ : InMux
    port map (
            O => \N__20268\,
            I => \N__20246\
        );

    \I__4390\ : InMux
    port map (
            O => \N__20267\,
            I => \N__20246\
        );

    \I__4389\ : Span4Mux_h
    port map (
            O => \N__20264\,
            I => \N__20241\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__20259\,
            I => \N__20241\
        );

    \I__4387\ : Odrv4
    port map (
            O => \N__20256\,
            I => bu_rx_data_4_rep2
        );

    \I__4386\ : Odrv4
    port map (
            O => \N__20251\,
            I => bu_rx_data_4_rep2
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__20246\,
            I => bu_rx_data_4_rep2
        );

    \I__4384\ : Odrv4
    port map (
            O => \N__20241\,
            I => bu_rx_data_4_rep2
        );

    \I__4383\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20229\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__20229\,
            I => \N__20226\
        );

    \I__4381\ : Odrv4
    port map (
            O => \N__20226\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_4_8\
        );

    \I__4380\ : CascadeMux
    port map (
            O => \N__20223\,
            I => \N__20211\
        );

    \I__4379\ : CascadeMux
    port map (
            O => \N__20222\,
            I => \N__20208\
        );

    \I__4378\ : CascadeMux
    port map (
            O => \N__20221\,
            I => \N__20202\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__20220\,
            I => \N__20199\
        );

    \I__4376\ : InMux
    port map (
            O => \N__20219\,
            I => \N__20193\
        );

    \I__4375\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20186\
        );

    \I__4374\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20186\
        );

    \I__4373\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20183\
        );

    \I__4372\ : InMux
    port map (
            O => \N__20215\,
            I => \N__20178\
        );

    \I__4371\ : InMux
    port map (
            O => \N__20214\,
            I => \N__20178\
        );

    \I__4370\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20169\
        );

    \I__4369\ : InMux
    port map (
            O => \N__20208\,
            I => \N__20169\
        );

    \I__4368\ : InMux
    port map (
            O => \N__20207\,
            I => \N__20169\
        );

    \I__4367\ : InMux
    port map (
            O => \N__20206\,
            I => \N__20169\
        );

    \I__4366\ : InMux
    port map (
            O => \N__20205\,
            I => \N__20160\
        );

    \I__4365\ : InMux
    port map (
            O => \N__20202\,
            I => \N__20160\
        );

    \I__4364\ : InMux
    port map (
            O => \N__20199\,
            I => \N__20160\
        );

    \I__4363\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20160\
        );

    \I__4362\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20152\
        );

    \I__4361\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20152\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__20193\,
            I => \N__20149\
        );

    \I__4359\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20144\
        );

    \I__4358\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20144\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__20186\,
            I => \N__20140\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__20183\,
            I => \N__20135\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__20178\,
            I => \N__20135\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__20169\,
            I => \N__20130\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__20160\,
            I => \N__20130\
        );

    \I__4352\ : InMux
    port map (
            O => \N__20159\,
            I => \N__20123\
        );

    \I__4351\ : InMux
    port map (
            O => \N__20158\,
            I => \N__20123\
        );

    \I__4350\ : InMux
    port map (
            O => \N__20157\,
            I => \N__20123\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__20152\,
            I => \N__20116\
        );

    \I__4348\ : Span4Mux_v
    port map (
            O => \N__20149\,
            I => \N__20116\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__20144\,
            I => \N__20116\
        );

    \I__4346\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20113\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__20140\,
            I => \N__20104\
        );

    \I__4344\ : Span4Mux_s2_v
    port map (
            O => \N__20135\,
            I => \N__20104\
        );

    \I__4343\ : Span4Mux_h
    port map (
            O => \N__20130\,
            I => \N__20104\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__20123\,
            I => \N__20104\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__20116\,
            I => \N__20099\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__20113\,
            I => \N__20099\
        );

    \I__4339\ : Odrv4
    port map (
            O => \N__20104\,
            I => \Lab_UT.dictrl.N_19_0\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__20099\,
            I => \Lab_UT.dictrl.N_19_0\
        );

    \I__4337\ : CascadeMux
    port map (
            O => \N__20094\,
            I => \N__20087\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__20093\,
            I => \N__20083\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__20092\,
            I => \N__20079\
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__20091\,
            I => \N__20072\
        );

    \I__4333\ : InMux
    port map (
            O => \N__20090\,
            I => \N__20067\
        );

    \I__4332\ : InMux
    port map (
            O => \N__20087\,
            I => \N__20064\
        );

    \I__4331\ : InMux
    port map (
            O => \N__20086\,
            I => \N__20055\
        );

    \I__4330\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20055\
        );

    \I__4329\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20055\
        );

    \I__4328\ : InMux
    port map (
            O => \N__20079\,
            I => \N__20055\
        );

    \I__4327\ : InMux
    port map (
            O => \N__20078\,
            I => \N__20050\
        );

    \I__4326\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20050\
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__20076\,
            I => \N__20046\
        );

    \I__4324\ : InMux
    port map (
            O => \N__20075\,
            I => \N__20040\
        );

    \I__4323\ : InMux
    port map (
            O => \N__20072\,
            I => \N__20040\
        );

    \I__4322\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20035\
        );

    \I__4321\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20035\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__20067\,
            I => \N__20032\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20028\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__20055\,
            I => \N__20023\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__20050\,
            I => \N__20023\
        );

    \I__4316\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20018\
        );

    \I__4315\ : InMux
    port map (
            O => \N__20046\,
            I => \N__20018\
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__20045\,
            I => \N__20015\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__20040\,
            I => \N__20012\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__20035\,
            I => \N__20009\
        );

    \I__4311\ : Span4Mux_s1_v
    port map (
            O => \N__20032\,
            I => \N__20006\
        );

    \I__4310\ : InMux
    port map (
            O => \N__20031\,
            I => \N__20003\
        );

    \I__4309\ : Span4Mux_h
    port map (
            O => \N__20028\,
            I => \N__19998\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__20023\,
            I => \N__19998\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__20018\,
            I => \N__19995\
        );

    \I__4306\ : InMux
    port map (
            O => \N__20015\,
            I => \N__19992\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__20012\,
            I => \N__19987\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__20009\,
            I => \N__19987\
        );

    \I__4303\ : Sp12to4
    port map (
            O => \N__20006\,
            I => \N__19982\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__19982\
        );

    \I__4301\ : Span4Mux_h
    port map (
            O => \N__19998\,
            I => \N__19979\
        );

    \I__4300\ : Span4Mux_h
    port map (
            O => \N__19995\,
            I => \N__19974\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19992\,
            I => \N__19974\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__19987\,
            I => \N__19971\
        );

    \I__4297\ : Odrv12
    port map (
            O => \N__19982\,
            I => bu_rx_data_6_rep2
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__19979\,
            I => bu_rx_data_6_rep2
        );

    \I__4295\ : Odrv4
    port map (
            O => \N__19974\,
            I => bu_rx_data_6_rep2
        );

    \I__4294\ : Odrv4
    port map (
            O => \N__19971\,
            I => bu_rx_data_6_rep2
        );

    \I__4293\ : InMux
    port map (
            O => \N__19962\,
            I => \N__19948\
        );

    \I__4292\ : InMux
    port map (
            O => \N__19961\,
            I => \N__19945\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19942\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19959\,
            I => \N__19939\
        );

    \I__4289\ : InMux
    port map (
            O => \N__19958\,
            I => \N__19936\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19957\,
            I => \N__19933\
        );

    \I__4287\ : InMux
    port map (
            O => \N__19956\,
            I => \N__19926\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19955\,
            I => \N__19926\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19926\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19921\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19952\,
            I => \N__19921\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19951\,
            I => \N__19918\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19914\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__19945\,
            I => \N__19909\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19942\,
            I => \N__19909\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19904\
        );

    \I__4277\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19904\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__19933\,
            I => \N__19901\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19898\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19921\,
            I => \N__19893\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__19918\,
            I => \N__19893\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19917\,
            I => \N__19890\
        );

    \I__4271\ : Span12Mux_s2_v
    port map (
            O => \N__19914\,
            I => \N__19885\
        );

    \I__4270\ : Span12Mux_v
    port map (
            O => \N__19909\,
            I => \N__19885\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__19904\,
            I => \N__19880\
        );

    \I__4268\ : Span4Mux_s2_v
    port map (
            O => \N__19901\,
            I => \N__19880\
        );

    \I__4267\ : Span4Mux_h
    port map (
            O => \N__19898\,
            I => \N__19875\
        );

    \I__4266\ : Span4Mux_s2_v
    port map (
            O => \N__19893\,
            I => \N__19875\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__19890\,
            I => \N__19872\
        );

    \I__4264\ : Odrv12
    port map (
            O => \N__19885\,
            I => \Lab_UT.dictrl.m40Z0Z_1\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__19880\,
            I => \Lab_UT.dictrl.m40Z0Z_1\
        );

    \I__4262\ : Odrv4
    port map (
            O => \N__19875\,
            I => \Lab_UT.dictrl.m40Z0Z_1\
        );

    \I__4261\ : Odrv12
    port map (
            O => \N__19872\,
            I => \Lab_UT.dictrl.m40Z0Z_1\
        );

    \I__4260\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19860\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__19860\,
            I => \N__19857\
        );

    \I__4258\ : Span4Mux_h
    port map (
            O => \N__19857\,
            I => \N__19854\
        );

    \I__4257\ : Odrv4
    port map (
            O => \N__19854\,
            I => \Lab_UT.dictrl.m53_d_1_4\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19851\,
            I => \N__19845\
        );

    \I__4255\ : InMux
    port map (
            O => \N__19850\,
            I => \N__19845\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19845\,
            I => \N__19840\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19844\,
            I => \N__19837\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19834\
        );

    \I__4251\ : Span4Mux_v
    port map (
            O => \N__19840\,
            I => \N__19825\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__19837\,
            I => \N__19825\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__19834\,
            I => \N__19816\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19833\,
            I => \N__19813\
        );

    \I__4247\ : InMux
    port map (
            O => \N__19832\,
            I => \N__19810\
        );

    \I__4246\ : InMux
    port map (
            O => \N__19831\,
            I => \N__19805\
        );

    \I__4245\ : InMux
    port map (
            O => \N__19830\,
            I => \N__19805\
        );

    \I__4244\ : Span4Mux_v
    port map (
            O => \N__19825\,
            I => \N__19802\
        );

    \I__4243\ : InMux
    port map (
            O => \N__19824\,
            I => \N__19799\
        );

    \I__4242\ : InMux
    port map (
            O => \N__19823\,
            I => \N__19788\
        );

    \I__4241\ : InMux
    port map (
            O => \N__19822\,
            I => \N__19788\
        );

    \I__4240\ : InMux
    port map (
            O => \N__19821\,
            I => \N__19788\
        );

    \I__4239\ : InMux
    port map (
            O => \N__19820\,
            I => \N__19788\
        );

    \I__4238\ : InMux
    port map (
            O => \N__19819\,
            I => \N__19788\
        );

    \I__4237\ : Span4Mux_s3_v
    port map (
            O => \N__19816\,
            I => \N__19783\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__19813\,
            I => \N__19783\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19780\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__19805\,
            I => \N__19775\
        );

    \I__4233\ : Span4Mux_s0_v
    port map (
            O => \N__19802\,
            I => \N__19768\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__19799\,
            I => \N__19768\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__19788\,
            I => \N__19768\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__19783\,
            I => \N__19762\
        );

    \I__4229\ : Span4Mux_v
    port map (
            O => \N__19780\,
            I => \N__19762\
        );

    \I__4228\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19757\
        );

    \I__4227\ : InMux
    port map (
            O => \N__19778\,
            I => \N__19757\
        );

    \I__4226\ : Span4Mux_v
    port map (
            O => \N__19775\,
            I => \N__19752\
        );

    \I__4225\ : Span4Mux_v
    port map (
            O => \N__19768\,
            I => \N__19752\
        );

    \I__4224\ : InMux
    port map (
            O => \N__19767\,
            I => \N__19749\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__19762\,
            I => \Lab_UT.dictrl.state_2_rep2\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__19757\,
            I => \Lab_UT.dictrl.state_2_rep2\
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__19752\,
            I => \Lab_UT.dictrl.state_2_rep2\
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__19749\,
            I => \Lab_UT.dictrl.state_2_rep2\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__19740\,
            I => \Lab_UT.dictrl.N_97_mux_6_cascade_\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__19737\,
            I => \N__19731\
        );

    \I__4217\ : CascadeMux
    port map (
            O => \N__19736\,
            I => \N__19726\
        );

    \I__4216\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19721\
        );

    \I__4215\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19717\
        );

    \I__4214\ : InMux
    port map (
            O => \N__19731\,
            I => \N__19707\
        );

    \I__4213\ : InMux
    port map (
            O => \N__19730\,
            I => \N__19704\
        );

    \I__4212\ : InMux
    port map (
            O => \N__19729\,
            I => \N__19701\
        );

    \I__4211\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19697\
        );

    \I__4210\ : InMux
    port map (
            O => \N__19725\,
            I => \N__19694\
        );

    \I__4209\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19691\
        );

    \I__4208\ : LocalMux
    port map (
            O => \N__19721\,
            I => \N__19688\
        );

    \I__4207\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19685\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19682\
        );

    \I__4205\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19679\
        );

    \I__4204\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19672\
        );

    \I__4203\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19672\
        );

    \I__4202\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19672\
        );

    \I__4201\ : InMux
    port map (
            O => \N__19712\,
            I => \N__19667\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19711\,
            I => \N__19667\
        );

    \I__4199\ : InMux
    port map (
            O => \N__19710\,
            I => \N__19662\
        );

    \I__4198\ : LocalMux
    port map (
            O => \N__19707\,
            I => \N__19655\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__19704\,
            I => \N__19655\
        );

    \I__4196\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19655\
        );

    \I__4195\ : InMux
    port map (
            O => \N__19700\,
            I => \N__19652\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__19697\,
            I => \N__19645\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__19694\,
            I => \N__19645\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__19691\,
            I => \N__19645\
        );

    \I__4191\ : Span4Mux_s2_v
    port map (
            O => \N__19688\,
            I => \N__19642\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__19685\,
            I => \N__19639\
        );

    \I__4189\ : Span4Mux_s2_v
    port map (
            O => \N__19682\,
            I => \N__19632\
        );

    \I__4188\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19632\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__19672\,
            I => \N__19632\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19629\
        );

    \I__4185\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19624\
        );

    \I__4184\ : InMux
    port map (
            O => \N__19665\,
            I => \N__19624\
        );

    \I__4183\ : LocalMux
    port map (
            O => \N__19662\,
            I => \N__19619\
        );

    \I__4182\ : Span4Mux_v
    port map (
            O => \N__19655\,
            I => \N__19619\
        );

    \I__4181\ : LocalMux
    port map (
            O => \N__19652\,
            I => \N__19610\
        );

    \I__4180\ : Span4Mux_s3_v
    port map (
            O => \N__19645\,
            I => \N__19610\
        );

    \I__4179\ : Span4Mux_v
    port map (
            O => \N__19642\,
            I => \N__19607\
        );

    \I__4178\ : Span4Mux_v
    port map (
            O => \N__19639\,
            I => \N__19596\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__19632\,
            I => \N__19596\
        );

    \I__4176\ : Span4Mux_v
    port map (
            O => \N__19629\,
            I => \N__19596\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__19624\,
            I => \N__19596\
        );

    \I__4174\ : Span4Mux_h
    port map (
            O => \N__19619\,
            I => \N__19596\
        );

    \I__4173\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19593\
        );

    \I__4172\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19590\
        );

    \I__4171\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19585\
        );

    \I__4170\ : InMux
    port map (
            O => \N__19615\,
            I => \N__19585\
        );

    \I__4169\ : Odrv4
    port map (
            O => \N__19610\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__19607\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4167\ : Odrv4
    port map (
            O => \N__19596\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__19593\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__19590\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__19585\,
            I => \Lab_UT.dictrl.state_3_rep2\
        );

    \I__4163\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19569\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19566\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__19566\,
            I => \N__19563\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__19563\,
            I => \N__19560\
        );

    \I__4159\ : Odrv4
    port map (
            O => \N__19560\,
            I => \Lab_UT.dictrl.g2_1_4\
        );

    \I__4158\ : InMux
    port map (
            O => \N__19557\,
            I => \N__19554\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__19554\,
            I => \Lab_UT.dictrl.N_1462_4\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__19551\,
            I => \Lab_UT.dictrl.N_1102_4_cascade_\
        );

    \I__4155\ : InMux
    port map (
            O => \N__19548\,
            I => \N__19545\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__19545\,
            I => \Lab_UT.dictrl.N_6_0\
        );

    \I__4153\ : CascadeMux
    port map (
            O => \N__19542\,
            I => \N__19539\
        );

    \I__4152\ : InMux
    port map (
            O => \N__19539\,
            I => \N__19535\
        );

    \I__4151\ : InMux
    port map (
            O => \N__19538\,
            I => \N__19529\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__19535\,
            I => \N__19524\
        );

    \I__4149\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19519\
        );

    \I__4148\ : InMux
    port map (
            O => \N__19533\,
            I => \N__19519\
        );

    \I__4147\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19516\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19513\
        );

    \I__4145\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19510\
        );

    \I__4144\ : CascadeMux
    port map (
            O => \N__19527\,
            I => \N__19507\
        );

    \I__4143\ : Span4Mux_s2_v
    port map (
            O => \N__19524\,
            I => \N__19502\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__19519\,
            I => \N__19502\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19497\
        );

    \I__4140\ : Span4Mux_s2_v
    port map (
            O => \N__19513\,
            I => \N__19497\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__19510\,
            I => \N__19494\
        );

    \I__4138\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19491\
        );

    \I__4137\ : Span4Mux_v
    port map (
            O => \N__19502\,
            I => \N__19488\
        );

    \I__4136\ : Span4Mux_v
    port map (
            O => \N__19497\,
            I => \N__19485\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__19494\,
            I => \N__19478\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__19491\,
            I => \N__19478\
        );

    \I__4133\ : Span4Mux_s2_h
    port map (
            O => \N__19488\,
            I => \N__19478\
        );

    \I__4132\ : Odrv4
    port map (
            O => \N__19485\,
            I => \Lab_UT.dictrl.next_state_2_1\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__19478\,
            I => \Lab_UT.dictrl.next_state_2_1\
        );

    \I__4130\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19470\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__19470\,
            I => \N__19467\
        );

    \I__4128\ : Span4Mux_h
    port map (
            O => \N__19467\,
            I => \N__19464\
        );

    \I__4127\ : Span4Mux_h
    port map (
            O => \N__19464\,
            I => \N__19461\
        );

    \I__4126\ : Odrv4
    port map (
            O => \N__19461\,
            I => \Lab_UT.dictrl.g0_i_0\
        );

    \I__4125\ : CascadeMux
    port map (
            O => \N__19458\,
            I => \N__19455\
        );

    \I__4124\ : InMux
    port map (
            O => \N__19455\,
            I => \N__19452\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__19452\,
            I => \Lab_UT.dictrl.g1_1_1_0\
        );

    \I__4122\ : InMux
    port map (
            O => \N__19449\,
            I => \N__19440\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19448\,
            I => \N__19440\
        );

    \I__4120\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19434\
        );

    \I__4119\ : InMux
    port map (
            O => \N__19446\,
            I => \N__19434\
        );

    \I__4118\ : InMux
    port map (
            O => \N__19445\,
            I => \N__19431\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__19440\,
            I => \N__19428\
        );

    \I__4116\ : InMux
    port map (
            O => \N__19439\,
            I => \N__19425\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19418\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__19431\,
            I => \N__19415\
        );

    \I__4113\ : Span4Mux_v
    port map (
            O => \N__19428\,
            I => \N__19412\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__19425\,
            I => \N__19409\
        );

    \I__4111\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19404\
        );

    \I__4110\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19404\
        );

    \I__4109\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19399\
        );

    \I__4108\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19399\
        );

    \I__4107\ : Span12Mux_s10_h
    port map (
            O => \N__19418\,
            I => \N__19396\
        );

    \I__4106\ : Span4Mux_v
    port map (
            O => \N__19415\,
            I => \N__19385\
        );

    \I__4105\ : Span4Mux_h
    port map (
            O => \N__19412\,
            I => \N__19385\
        );

    \I__4104\ : Span4Mux_v
    port map (
            O => \N__19409\,
            I => \N__19385\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19385\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__19399\,
            I => \N__19385\
        );

    \I__4101\ : Odrv12
    port map (
            O => \N__19396\,
            I => bu_rx_data_7_rep1
        );

    \I__4100\ : Odrv4
    port map (
            O => \N__19385\,
            I => bu_rx_data_7_rep1
        );

    \I__4099\ : InMux
    port map (
            O => \N__19380\,
            I => \N__19377\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__19377\,
            I => \N__19374\
        );

    \I__4097\ : Span4Mux_h
    port map (
            O => \N__19374\,
            I => \N__19371\
        );

    \I__4096\ : Odrv4
    port map (
            O => \N__19371\,
            I => \Lab_UT.dictrl.N_59\
        );

    \I__4095\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19363\
        );

    \I__4094\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19358\
        );

    \I__4093\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19358\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__19363\,
            I => \N__19352\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__19358\,
            I => \N__19352\
        );

    \I__4090\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19348\
        );

    \I__4089\ : Span4Mux_v
    port map (
            O => \N__19352\,
            I => \N__19345\
        );

    \I__4088\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19342\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__19348\,
            I => \Lab_UT.dictrl.N_97_mux\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__19345\,
            I => \Lab_UT.dictrl.N_97_mux\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__19342\,
            I => \Lab_UT.dictrl.N_97_mux\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__19335\,
            I => \Lab_UT.dictrl.N_59_cascade_\
        );

    \I__4083\ : InMux
    port map (
            O => \N__19332\,
            I => \N__19321\
        );

    \I__4082\ : InMux
    port map (
            O => \N__19331\,
            I => \N__19321\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__19330\,
            I => \N__19318\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__19329\,
            I => \N__19307\
        );

    \I__4079\ : InMux
    port map (
            O => \N__19328\,
            I => \N__19298\
        );

    \I__4078\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19298\
        );

    \I__4077\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19298\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__19321\,
            I => \N__19295\
        );

    \I__4075\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19290\
        );

    \I__4074\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19290\
        );

    \I__4073\ : InMux
    port map (
            O => \N__19316\,
            I => \N__19285\
        );

    \I__4072\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19285\
        );

    \I__4071\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19280\
        );

    \I__4070\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19280\
        );

    \I__4069\ : InMux
    port map (
            O => \N__19312\,
            I => \N__19275\
        );

    \I__4068\ : InMux
    port map (
            O => \N__19311\,
            I => \N__19275\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__19310\,
            I => \N__19272\
        );

    \I__4066\ : InMux
    port map (
            O => \N__19307\,
            I => \N__19264\
        );

    \I__4065\ : InMux
    port map (
            O => \N__19306\,
            I => \N__19264\
        );

    \I__4064\ : InMux
    port map (
            O => \N__19305\,
            I => \N__19264\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__19298\,
            I => \N__19261\
        );

    \I__4062\ : Span4Mux_h
    port map (
            O => \N__19295\,
            I => \N__19256\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__19290\,
            I => \N__19256\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__19285\,
            I => \N__19249\
        );

    \I__4059\ : LocalMux
    port map (
            O => \N__19280\,
            I => \N__19249\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__19275\,
            I => \N__19249\
        );

    \I__4057\ : InMux
    port map (
            O => \N__19272\,
            I => \N__19246\
        );

    \I__4056\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19243\
        );

    \I__4055\ : LocalMux
    port map (
            O => \N__19264\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__19261\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4053\ : Odrv4
    port map (
            O => \N__19256\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4052\ : Odrv12
    port map (
            O => \N__19249\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__19246\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__19243\,
            I => \Lab_UT.dictrl.state_0_rep2\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__19230\,
            I => \Lab_UT.dictrl.N_40_5_cascade_\
        );

    \I__4048\ : InMux
    port map (
            O => \N__19227\,
            I => \N__19223\
        );

    \I__4047\ : InMux
    port map (
            O => \N__19226\,
            I => \N__19220\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__19223\,
            I => \Lab_UT.dictrl.N_40_4\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__19220\,
            I => \Lab_UT.dictrl.N_40_4\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__19215\,
            I => \Lab_UT.dictrl.N_40_2_cascade_\
        );

    \I__4043\ : InMux
    port map (
            O => \N__19212\,
            I => \N__19205\
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__19211\,
            I => \N__19200\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__19210\,
            I => \N__19194\
        );

    \I__4040\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19185\
        );

    \I__4039\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19185\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__19205\,
            I => \N__19182\
        );

    \I__4037\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19177\
        );

    \I__4036\ : InMux
    port map (
            O => \N__19203\,
            I => \N__19177\
        );

    \I__4035\ : InMux
    port map (
            O => \N__19200\,
            I => \N__19172\
        );

    \I__4034\ : InMux
    port map (
            O => \N__19199\,
            I => \N__19172\
        );

    \I__4033\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19165\
        );

    \I__4032\ : InMux
    port map (
            O => \N__19197\,
            I => \N__19165\
        );

    \I__4031\ : InMux
    port map (
            O => \N__19194\,
            I => \N__19165\
        );

    \I__4030\ : CascadeMux
    port map (
            O => \N__19193\,
            I => \N__19161\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__19192\,
            I => \N__19158\
        );

    \I__4028\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19154\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__19190\,
            I => \N__19151\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__19185\,
            I => \N__19146\
        );

    \I__4025\ : Span4Mux_s3_h
    port map (
            O => \N__19182\,
            I => \N__19143\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__19177\,
            I => \N__19140\
        );

    \I__4023\ : LocalMux
    port map (
            O => \N__19172\,
            I => \N__19137\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__19165\,
            I => \N__19134\
        );

    \I__4021\ : InMux
    port map (
            O => \N__19164\,
            I => \N__19129\
        );

    \I__4020\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19129\
        );

    \I__4019\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19124\
        );

    \I__4018\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19124\
        );

    \I__4017\ : LocalMux
    port map (
            O => \N__19154\,
            I => \N__19121\
        );

    \I__4016\ : InMux
    port map (
            O => \N__19151\,
            I => \N__19118\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__19150\,
            I => \N__19112\
        );

    \I__4014\ : InMux
    port map (
            O => \N__19149\,
            I => \N__19109\
        );

    \I__4013\ : Span4Mux_s3_h
    port map (
            O => \N__19146\,
            I => \N__19106\
        );

    \I__4012\ : Sp12to4
    port map (
            O => \N__19143\,
            I => \N__19101\
        );

    \I__4011\ : Span12Mux_s8_h
    port map (
            O => \N__19140\,
            I => \N__19101\
        );

    \I__4010\ : Span4Mux_v
    port map (
            O => \N__19137\,
            I => \N__19094\
        );

    \I__4009\ : Span4Mux_v
    port map (
            O => \N__19134\,
            I => \N__19094\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__19129\,
            I => \N__19094\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19091\
        );

    \I__4006\ : Span4Mux_s3_h
    port map (
            O => \N__19121\,
            I => \N__19088\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__19118\,
            I => \N__19085\
        );

    \I__4004\ : InMux
    port map (
            O => \N__19117\,
            I => \N__19076\
        );

    \I__4003\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19076\
        );

    \I__4002\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19076\
        );

    \I__4001\ : InMux
    port map (
            O => \N__19112\,
            I => \N__19076\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__19109\,
            I => bu_rx_data_6
        );

    \I__3999\ : Odrv4
    port map (
            O => \N__19106\,
            I => bu_rx_data_6
        );

    \I__3998\ : Odrv12
    port map (
            O => \N__19101\,
            I => bu_rx_data_6
        );

    \I__3997\ : Odrv4
    port map (
            O => \N__19094\,
            I => bu_rx_data_6
        );

    \I__3996\ : Odrv4
    port map (
            O => \N__19091\,
            I => bu_rx_data_6
        );

    \I__3995\ : Odrv4
    port map (
            O => \N__19088\,
            I => bu_rx_data_6
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__19085\,
            I => bu_rx_data_6
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__19076\,
            I => bu_rx_data_6
        );

    \I__3992\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19056\
        );

    \I__3991\ : LocalMux
    port map (
            O => \N__19056\,
            I => \Lab_UT.dictrl.g0_i_a4_1_5\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__19053\,
            I => \Lab_UT.dictrl.g0_i_a4_1_4_cascade_\
        );

    \I__3989\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19042\
        );

    \I__3988\ : InMux
    port map (
            O => \N__19049\,
            I => \N__19042\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__19048\,
            I => \N__19037\
        );

    \I__3986\ : InMux
    port map (
            O => \N__19047\,
            I => \N__19033\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19030\
        );

    \I__3984\ : InMux
    port map (
            O => \N__19041\,
            I => \N__19023\
        );

    \I__3983\ : InMux
    port map (
            O => \N__19040\,
            I => \N__19023\
        );

    \I__3982\ : InMux
    port map (
            O => \N__19037\,
            I => \N__19023\
        );

    \I__3981\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19020\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__19033\,
            I => \N__19014\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__19030\,
            I => \N__19009\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__19023\,
            I => \N__19009\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__19020\,
            I => \N__19006\
        );

    \I__3976\ : InMux
    port map (
            O => \N__19019\,
            I => \N__18999\
        );

    \I__3975\ : InMux
    port map (
            O => \N__19018\,
            I => \N__18999\
        );

    \I__3974\ : InMux
    port map (
            O => \N__19017\,
            I => \N__18999\
        );

    \I__3973\ : Span12Mux_s3_h
    port map (
            O => \N__19014\,
            I => \N__18991\
        );

    \I__3972\ : Span4Mux_h
    port map (
            O => \N__19009\,
            I => \N__18988\
        );

    \I__3971\ : Span4Mux_s3_h
    port map (
            O => \N__19006\,
            I => \N__18985\
        );

    \I__3970\ : LocalMux
    port map (
            O => \N__18999\,
            I => \N__18982\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18998\,
            I => \N__18971\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18997\,
            I => \N__18971\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18996\,
            I => \N__18971\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18995\,
            I => \N__18971\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18994\,
            I => \N__18971\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__18991\,
            I => bu_rx_data_5
        );

    \I__3963\ : Odrv4
    port map (
            O => \N__18988\,
            I => bu_rx_data_5
        );

    \I__3962\ : Odrv4
    port map (
            O => \N__18985\,
            I => bu_rx_data_5
        );

    \I__3961\ : Odrv12
    port map (
            O => \N__18982\,
            I => bu_rx_data_5
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18971\,
            I => bu_rx_data_5
        );

    \I__3959\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18957\
        );

    \I__3958\ : LocalMux
    port map (
            O => \N__18957\,
            I => \N__18954\
        );

    \I__3957\ : Span4Mux_h
    port map (
            O => \N__18954\,
            I => \N__18951\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__18951\,
            I => \Lab_UT.dictrl.N_12\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18948\,
            I => \N__18945\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18945\,
            I => \N__18942\
        );

    \I__3953\ : Odrv12
    port map (
            O => \N__18942\,
            I => \Lab_UT.dictrl.N_4\
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__18939\,
            I => \N__18928\
        );

    \I__3951\ : CascadeMux
    port map (
            O => \N__18938\,
            I => \N__18924\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18921\
        );

    \I__3949\ : InMux
    port map (
            O => \N__18936\,
            I => \N__18914\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18935\,
            I => \N__18914\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__18934\,
            I => \N__18911\
        );

    \I__3946\ : InMux
    port map (
            O => \N__18933\,
            I => \N__18906\
        );

    \I__3945\ : InMux
    port map (
            O => \N__18932\,
            I => \N__18901\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18931\,
            I => \N__18901\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18928\,
            I => \N__18898\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18927\,
            I => \N__18893\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18924\,
            I => \N__18893\
        );

    \I__3940\ : InMux
    port map (
            O => \N__18921\,
            I => \N__18886\
        );

    \I__3939\ : InMux
    port map (
            O => \N__18920\,
            I => \N__18886\
        );

    \I__3938\ : CascadeMux
    port map (
            O => \N__18919\,
            I => \N__18883\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18914\,
            I => \N__18880\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18911\,
            I => \N__18877\
        );

    \I__3935\ : InMux
    port map (
            O => \N__18910\,
            I => \N__18872\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18909\,
            I => \N__18869\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__18906\,
            I => \N__18864\
        );

    \I__3932\ : LocalMux
    port map (
            O => \N__18901\,
            I => \N__18864\
        );

    \I__3931\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18861\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__18893\,
            I => \N__18858\
        );

    \I__3929\ : CascadeMux
    port map (
            O => \N__18892\,
            I => \N__18855\
        );

    \I__3928\ : InMux
    port map (
            O => \N__18891\,
            I => \N__18850\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__18886\,
            I => \N__18847\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18883\,
            I => \N__18844\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__18880\,
            I => \N__18839\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18877\,
            I => \N__18839\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18876\,
            I => \N__18834\
        );

    \I__3922\ : InMux
    port map (
            O => \N__18875\,
            I => \N__18834\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__18872\,
            I => \N__18831\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__18869\,
            I => \N__18822\
        );

    \I__3919\ : Span4Mux_v
    port map (
            O => \N__18864\,
            I => \N__18822\
        );

    \I__3918\ : Span4Mux_v
    port map (
            O => \N__18861\,
            I => \N__18822\
        );

    \I__3917\ : Span4Mux_v
    port map (
            O => \N__18858\,
            I => \N__18822\
        );

    \I__3916\ : InMux
    port map (
            O => \N__18855\,
            I => \N__18817\
        );

    \I__3915\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18817\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18853\,
            I => \N__18814\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__18850\,
            I => \N__18811\
        );

    \I__3912\ : Span4Mux_v
    port map (
            O => \N__18847\,
            I => \N__18804\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__18844\,
            I => \N__18804\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__18839\,
            I => \N__18804\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__18834\,
            I => \N__18797\
        );

    \I__3908\ : Span4Mux_v
    port map (
            O => \N__18831\,
            I => \N__18797\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__18822\,
            I => \N__18797\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__18817\,
            I => \N__18792\
        );

    \I__3905\ : LocalMux
    port map (
            O => \N__18814\,
            I => \N__18792\
        );

    \I__3904\ : Span4Mux_h
    port map (
            O => \N__18811\,
            I => \N__18787\
        );

    \I__3903\ : Span4Mux_h
    port map (
            O => \N__18804\,
            I => \N__18787\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__18797\,
            I => bu_rx_data_4
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__18792\,
            I => bu_rx_data_4
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__18787\,
            I => bu_rx_data_4
        );

    \I__3899\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18777\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18777\,
            I => \N__18774\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__18774\,
            I => \Lab_UT.dictrl.N_7\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__18771\,
            I => \N__18768\
        );

    \I__3895\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18765\
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__18765\,
            I => \N__18760\
        );

    \I__3893\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18756\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__18763\,
            I => \N__18753\
        );

    \I__3891\ : Span4Mux_v
    port map (
            O => \N__18760\,
            I => \N__18747\
        );

    \I__3890\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18744\
        );

    \I__3889\ : LocalMux
    port map (
            O => \N__18756\,
            I => \N__18741\
        );

    \I__3888\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18737\
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__18752\,
            I => \N__18734\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__18751\,
            I => \N__18731\
        );

    \I__3885\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18726\
        );

    \I__3884\ : Span4Mux_h
    port map (
            O => \N__18747\,
            I => \N__18719\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__18744\,
            I => \N__18719\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__18741\,
            I => \N__18716\
        );

    \I__3881\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18713\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__18737\,
            I => \N__18710\
        );

    \I__3879\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18701\
        );

    \I__3878\ : InMux
    port map (
            O => \N__18731\,
            I => \N__18701\
        );

    \I__3877\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18701\
        );

    \I__3876\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18701\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__18726\,
            I => \N__18698\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__18725\,
            I => \N__18695\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__18724\,
            I => \N__18692\
        );

    \I__3872\ : Span4Mux_h
    port map (
            O => \N__18719\,
            I => \N__18689\
        );

    \I__3871\ : Span4Mux_v
    port map (
            O => \N__18716\,
            I => \N__18686\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18713\,
            I => \N__18679\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__18710\,
            I => \N__18679\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18679\
        );

    \I__3867\ : Span4Mux_v
    port map (
            O => \N__18698\,
            I => \N__18676\
        );

    \I__3866\ : InMux
    port map (
            O => \N__18695\,
            I => \N__18673\
        );

    \I__3865\ : InMux
    port map (
            O => \N__18692\,
            I => \N__18670\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__18689\,
            I => \N__18665\
        );

    \I__3863\ : Span4Mux_h
    port map (
            O => \N__18686\,
            I => \N__18665\
        );

    \I__3862\ : Span4Mux_h
    port map (
            O => \N__18679\,
            I => \N__18662\
        );

    \I__3861\ : Odrv4
    port map (
            O => \N__18676\,
            I => bu_rx_data_3_rep2
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__18673\,
            I => bu_rx_data_3_rep2
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__18670\,
            I => bu_rx_data_3_rep2
        );

    \I__3858\ : Odrv4
    port map (
            O => \N__18665\,
            I => bu_rx_data_3_rep2
        );

    \I__3857\ : Odrv4
    port map (
            O => \N__18662\,
            I => bu_rx_data_3_rep2
        );

    \I__3856\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18646\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18650\,
            I => \N__18641\
        );

    \I__3854\ : InMux
    port map (
            O => \N__18649\,
            I => \N__18641\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18638\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__18641\,
            I => \N__18635\
        );

    \I__3851\ : Odrv12
    port map (
            O => \N__18638\,
            I => \Lab_UT.N_115\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__18635\,
            I => \Lab_UT.N_115\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18630\,
            I => \N__18627\
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__18627\,
            I => \N__18622\
        );

    \I__3847\ : InMux
    port map (
            O => \N__18626\,
            I => \N__18617\
        );

    \I__3846\ : InMux
    port map (
            O => \N__18625\,
            I => \N__18617\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__18622\,
            I => \N__18614\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__18617\,
            I => \N__18611\
        );

    \I__3843\ : Odrv4
    port map (
            O => \N__18614\,
            I => \Lab_UT.dictrl.N_39\
        );

    \I__3842\ : Odrv12
    port map (
            O => \N__18611\,
            I => \Lab_UT.dictrl.N_39\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__18606\,
            I => \N__18599\
        );

    \I__3840\ : CascadeMux
    port map (
            O => \N__18605\,
            I => \N__18596\
        );

    \I__3839\ : CascadeMux
    port map (
            O => \N__18604\,
            I => \N__18591\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__18603\,
            I => \N__18588\
        );

    \I__3837\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18580\
        );

    \I__3836\ : InMux
    port map (
            O => \N__18599\,
            I => \N__18580\
        );

    \I__3835\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18577\
        );

    \I__3834\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18574\
        );

    \I__3833\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18571\
        );

    \I__3832\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18566\
        );

    \I__3831\ : InMux
    port map (
            O => \N__18588\,
            I => \N__18563\
        );

    \I__3830\ : InMux
    port map (
            O => \N__18587\,
            I => \N__18560\
        );

    \I__3829\ : InMux
    port map (
            O => \N__18586\,
            I => \N__18556\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__18585\,
            I => \N__18553\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__18580\,
            I => \N__18548\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__18577\,
            I => \N__18548\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__18574\,
            I => \N__18545\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__18571\,
            I => \N__18542\
        );

    \I__3823\ : InMux
    port map (
            O => \N__18570\,
            I => \N__18537\
        );

    \I__3822\ : InMux
    port map (
            O => \N__18569\,
            I => \N__18537\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18532\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18532\
        );

    \I__3819\ : LocalMux
    port map (
            O => \N__18560\,
            I => \N__18529\
        );

    \I__3818\ : InMux
    port map (
            O => \N__18559\,
            I => \N__18526\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__18556\,
            I => \N__18523\
        );

    \I__3816\ : InMux
    port map (
            O => \N__18553\,
            I => \N__18520\
        );

    \I__3815\ : Span4Mux_v
    port map (
            O => \N__18548\,
            I => \N__18517\
        );

    \I__3814\ : Span4Mux_v
    port map (
            O => \N__18545\,
            I => \N__18512\
        );

    \I__3813\ : Span4Mux_v
    port map (
            O => \N__18542\,
            I => \N__18512\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__18537\,
            I => \N__18509\
        );

    \I__3811\ : Span4Mux_s3_v
    port map (
            O => \N__18532\,
            I => \N__18506\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__18529\,
            I => \N__18503\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__18526\,
            I => \N__18496\
        );

    \I__3808\ : Span4Mux_v
    port map (
            O => \N__18523\,
            I => \N__18496\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__18520\,
            I => \N__18496\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__18517\,
            I => \N__18491\
        );

    \I__3805\ : Span4Mux_v
    port map (
            O => \N__18512\,
            I => \N__18491\
        );

    \I__3804\ : Span4Mux_v
    port map (
            O => \N__18509\,
            I => \N__18488\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__18506\,
            I => \N__18485\
        );

    \I__3802\ : Span4Mux_v
    port map (
            O => \N__18503\,
            I => \N__18480\
        );

    \I__3801\ : Span4Mux_h
    port map (
            O => \N__18496\,
            I => \N__18480\
        );

    \I__3800\ : Odrv4
    port map (
            O => \N__18491\,
            I => bu_rx_data_6_rep1
        );

    \I__3799\ : Odrv4
    port map (
            O => \N__18488\,
            I => bu_rx_data_6_rep1
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__18485\,
            I => bu_rx_data_6_rep1
        );

    \I__3797\ : Odrv4
    port map (
            O => \N__18480\,
            I => bu_rx_data_6_rep1
        );

    \I__3796\ : InMux
    port map (
            O => \N__18471\,
            I => \N__18468\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__18468\,
            I => \N__18465\
        );

    \I__3794\ : Span4Mux_h
    port map (
            O => \N__18465\,
            I => \N__18462\
        );

    \I__3793\ : Odrv4
    port map (
            O => \N__18462\,
            I => \Lab_UT.dictrl.m53_d_1_0\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \Lab_UT.dictrl.N_97_mux_2_cascade_\
        );

    \I__3791\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18453\
        );

    \I__3790\ : LocalMux
    port map (
            O => \N__18453\,
            I => \N__18450\
        );

    \I__3789\ : Span4Mux_v
    port map (
            O => \N__18450\,
            I => \N__18447\
        );

    \I__3788\ : Odrv4
    port map (
            O => \N__18447\,
            I => \Lab_UT.dictrl.g2_1\
        );

    \I__3787\ : InMux
    port map (
            O => \N__18444\,
            I => \N__18441\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__18441\,
            I => \N__18438\
        );

    \I__3785\ : Odrv4
    port map (
            O => \N__18438\,
            I => \Lab_UT.dictrl.N_1462_0\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__18435\,
            I => \Lab_UT.dictrl.N_1102_0_cascade_\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__18432\,
            I => \N__18428\
        );

    \I__3782\ : InMux
    port map (
            O => \N__18431\,
            I => \N__18425\
        );

    \I__3781\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18422\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__18425\,
            I => \Lab_UT.dictrl.N_97_mux_7\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__18422\,
            I => \Lab_UT.dictrl.N_97_mux_7\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__18417\,
            I => \Lab_UT.dictrl.N_1106_1_cascade_\
        );

    \I__3777\ : CascadeMux
    port map (
            O => \N__18414\,
            I => \Lab_UT.didp.countrce4.q_5_0_cascade_\
        );

    \I__3776\ : InMux
    port map (
            O => \N__18411\,
            I => \N__18408\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__18408\,
            I => \N__18403\
        );

    \I__3774\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18400\
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__18406\,
            I => \N__18396\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__18403\,
            I => \N__18392\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__18400\,
            I => \N__18389\
        );

    \I__3770\ : InMux
    port map (
            O => \N__18399\,
            I => \N__18382\
        );

    \I__3769\ : InMux
    port map (
            O => \N__18396\,
            I => \N__18382\
        );

    \I__3768\ : InMux
    port map (
            O => \N__18395\,
            I => \N__18382\
        );

    \I__3767\ : Odrv4
    port map (
            O => \N__18392\,
            I => \Lab_UT.LdMtens\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__18389\,
            I => \Lab_UT.LdMtens\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__18382\,
            I => \Lab_UT.LdMtens\
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__18375\,
            I => \Lab_UT.didp.countrce4.q_5_1_cascade_\
        );

    \I__3763\ : InMux
    port map (
            O => \N__18372\,
            I => \N__18368\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18365\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__18368\,
            I => \N__18360\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__18365\,
            I => \N__18360\
        );

    \I__3759\ : Span4Mux_h
    port map (
            O => \N__18360\,
            I => \N__18356\
        );

    \I__3758\ : InMux
    port map (
            O => \N__18359\,
            I => \N__18353\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__18356\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__18353\,
            I => \Lab_UT.didp.un1_dicLdMtens_0\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__18348\,
            I => \N__18342\
        );

    \I__3754\ : InMux
    port map (
            O => \N__18347\,
            I => \N__18328\
        );

    \I__3753\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18328\
        );

    \I__3752\ : InMux
    port map (
            O => \N__18345\,
            I => \N__18328\
        );

    \I__3751\ : InMux
    port map (
            O => \N__18342\,
            I => \N__18328\
        );

    \I__3750\ : InMux
    port map (
            O => \N__18341\,
            I => \N__18325\
        );

    \I__3749\ : InMux
    port map (
            O => \N__18340\,
            I => \N__18316\
        );

    \I__3748\ : InMux
    port map (
            O => \N__18339\,
            I => \N__18316\
        );

    \I__3747\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18313\
        );

    \I__3746\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18310\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__18328\,
            I => \N__18307\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__18325\,
            I => \N__18304\
        );

    \I__3743\ : InMux
    port map (
            O => \N__18324\,
            I => \N__18297\
        );

    \I__3742\ : InMux
    port map (
            O => \N__18323\,
            I => \N__18297\
        );

    \I__3741\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18297\
        );

    \I__3740\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18294\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__18316\,
            I => \N__18291\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__18313\,
            I => \N__18288\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18284\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__18307\,
            I => \N__18275\
        );

    \I__3735\ : Span4Mux_s3_v
    port map (
            O => \N__18304\,
            I => \N__18275\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__18297\,
            I => \N__18275\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__18294\,
            I => \N__18275\
        );

    \I__3732\ : Span4Mux_s3_h
    port map (
            O => \N__18291\,
            I => \N__18272\
        );

    \I__3731\ : Span4Mux_v
    port map (
            O => \N__18288\,
            I => \N__18268\
        );

    \I__3730\ : InMux
    port map (
            O => \N__18287\,
            I => \N__18265\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__18284\,
            I => \N__18260\
        );

    \I__3728\ : Span4Mux_h
    port map (
            O => \N__18275\,
            I => \N__18260\
        );

    \I__3727\ : Span4Mux_h
    port map (
            O => \N__18272\,
            I => \N__18257\
        );

    \I__3726\ : InMux
    port map (
            O => \N__18271\,
            I => \N__18254\
        );

    \I__3725\ : Odrv4
    port map (
            O => \N__18268\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__18265\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__3723\ : Odrv4
    port map (
            O => \N__18260\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__3722\ : Odrv4
    port map (
            O => \N__18257\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__18254\,
            I => \Lab_UT.dictrl.state_0_rep1\
        );

    \I__3720\ : InMux
    port map (
            O => \N__18243\,
            I => \N__18240\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__18240\,
            I => \N__18237\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__18237\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0\
        );

    \I__3717\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18229\
        );

    \I__3716\ : InMux
    port map (
            O => \N__18233\,
            I => \N__18226\
        );

    \I__3715\ : InMux
    port map (
            O => \N__18232\,
            I => \N__18221\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__18229\,
            I => \N__18218\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__18226\,
            I => \N__18214\
        );

    \I__3712\ : InMux
    port map (
            O => \N__18225\,
            I => \N__18211\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__18224\,
            I => \N__18208\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__18221\,
            I => \N__18203\
        );

    \I__3709\ : Span4Mux_v
    port map (
            O => \N__18218\,
            I => \N__18203\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__18217\,
            I => \N__18200\
        );

    \I__3707\ : Span4Mux_v
    port map (
            O => \N__18214\,
            I => \N__18194\
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__18211\,
            I => \N__18194\
        );

    \I__3705\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18191\
        );

    \I__3704\ : Span4Mux_h
    port map (
            O => \N__18203\,
            I => \N__18188\
        );

    \I__3703\ : InMux
    port map (
            O => \N__18200\,
            I => \N__18185\
        );

    \I__3702\ : InMux
    port map (
            O => \N__18199\,
            I => \N__18182\
        );

    \I__3701\ : Odrv4
    port map (
            O => \N__18194\,
            I => \Lab_UT.state_i_4_0\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__18191\,
            I => \Lab_UT.state_i_4_0\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__18188\,
            I => \Lab_UT.state_i_4_0\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__18185\,
            I => \Lab_UT.state_i_4_0\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__18182\,
            I => \Lab_UT.state_i_4_0\
        );

    \I__3696\ : InMux
    port map (
            O => \N__18171\,
            I => \N__18167\
        );

    \I__3695\ : InMux
    port map (
            O => \N__18170\,
            I => \N__18164\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__18167\,
            I => \Lab_UT.dicRun_2\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__18164\,
            I => \Lab_UT.dicRun_2\
        );

    \I__3692\ : InMux
    port map (
            O => \N__18159\,
            I => \N__18145\
        );

    \I__3691\ : InMux
    port map (
            O => \N__18158\,
            I => \N__18145\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__18157\,
            I => \N__18142\
        );

    \I__3689\ : InMux
    port map (
            O => \N__18156\,
            I => \N__18138\
        );

    \I__3688\ : InMux
    port map (
            O => \N__18155\,
            I => \N__18130\
        );

    \I__3687\ : InMux
    port map (
            O => \N__18154\,
            I => \N__18130\
        );

    \I__3686\ : InMux
    port map (
            O => \N__18153\,
            I => \N__18130\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__18152\,
            I => \N__18126\
        );

    \I__3684\ : InMux
    port map (
            O => \N__18151\,
            I => \N__18123\
        );

    \I__3683\ : InMux
    port map (
            O => \N__18150\,
            I => \N__18120\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__18145\,
            I => \N__18117\
        );

    \I__3681\ : InMux
    port map (
            O => \N__18142\,
            I => \N__18114\
        );

    \I__3680\ : CascadeMux
    port map (
            O => \N__18141\,
            I => \N__18111\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__18138\,
            I => \N__18108\
        );

    \I__3678\ : InMux
    port map (
            O => \N__18137\,
            I => \N__18105\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__18130\,
            I => \N__18102\
        );

    \I__3676\ : InMux
    port map (
            O => \N__18129\,
            I => \N__18099\
        );

    \I__3675\ : InMux
    port map (
            O => \N__18126\,
            I => \N__18096\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__18123\,
            I => \N__18087\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__18120\,
            I => \N__18087\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__18117\,
            I => \N__18087\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18087\
        );

    \I__3670\ : InMux
    port map (
            O => \N__18111\,
            I => \N__18084\
        );

    \I__3669\ : Span4Mux_v
    port map (
            O => \N__18108\,
            I => \N__18079\
        );

    \I__3668\ : LocalMux
    port map (
            O => \N__18105\,
            I => \N__18079\
        );

    \I__3667\ : Span4Mux_h
    port map (
            O => \N__18102\,
            I => \N__18076\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__18099\,
            I => \N__18071\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__18096\,
            I => \N__18071\
        );

    \I__3664\ : Span4Mux_v
    port map (
            O => \N__18087\,
            I => \N__18066\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__18084\,
            I => \N__18066\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__18079\,
            I => \N__18063\
        );

    \I__3661\ : Span4Mux_h
    port map (
            O => \N__18076\,
            I => \N__18060\
        );

    \I__3660\ : Span4Mux_v
    port map (
            O => \N__18071\,
            I => \N__18055\
        );

    \I__3659\ : Span4Mux_h
    port map (
            O => \N__18066\,
            I => \N__18055\
        );

    \I__3658\ : Odrv4
    port map (
            O => \N__18063\,
            I => bu_rx_data_7
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__18060\,
            I => bu_rx_data_7
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__18055\,
            I => bu_rx_data_7
        );

    \I__3655\ : InMux
    port map (
            O => \N__18048\,
            I => \N__18045\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__18045\,
            I => \N__18042\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__18042\,
            I => \Lab_UT.didp.countrce1.q_5_1\
        );

    \I__3652\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__18036\,
            I => \N__18033\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__18033\,
            I => \N__18029\
        );

    \I__3649\ : InMux
    port map (
            O => \N__18032\,
            I => \N__18026\
        );

    \I__3648\ : Odrv4
    port map (
            O => \N__18029\,
            I => \Lab_UT.LdASones\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__18026\,
            I => \Lab_UT.LdASones\
        );

    \I__3646\ : CEMux
    port map (
            O => \N__18021\,
            I => \N__18018\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__18018\,
            I => \N__18015\
        );

    \I__3644\ : Span4Mux_h
    port map (
            O => \N__18015\,
            I => \N__18011\
        );

    \I__3643\ : CEMux
    port map (
            O => \N__18014\,
            I => \N__18008\
        );

    \I__3642\ : Odrv4
    port map (
            O => \N__18011\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__18008\,
            I => \Lab_UT.didp.regrce1.LdASones_0\
        );

    \I__3640\ : InMux
    port map (
            O => \N__18003\,
            I => \N__18000\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__18000\,
            I => \N__17995\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17999\,
            I => \N__17992\
        );

    \I__3637\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17989\
        );

    \I__3636\ : Odrv4
    port map (
            O => \N__17995\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17992\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17989\,
            I => \Lab_UT.di_ASones_0\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__17982\,
            I => \N__17979\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17976\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17976\,
            I => \N__17973\
        );

    \I__3630\ : Odrv12
    port map (
            O => \N__17973\,
            I => \Lab_UT.dispString.N_180\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17970\,
            I => \N__17967\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17967\,
            I => \Lab_UT.dispString.m49Z0Z_7\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17964\,
            I => \N__17961\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__17961\,
            I => \Lab_UT.dispString.m49Z0Z_11\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__17958\,
            I => \Lab_UT.didp.countrce1.q_5_0_cascade_\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \N__17950\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__17954\,
            I => \N__17947\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17953\,
            I => \N__17940\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17940\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17947\,
            I => \N__17940\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17932\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17939\,
            I => \N__17929\
        );

    \I__3617\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17920\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17920\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17936\,
            I => \N__17920\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17935\,
            I => \N__17920\
        );

    \I__3613\ : Odrv4
    port map (
            O => \N__17932\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__17929\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__17920\,
            I => \Lab_UT.di_Sones_0\
        );

    \I__3610\ : CascadeMux
    port map (
            O => \N__17913\,
            I => \Lab_UT.LdMtens_cascade_\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__17910\,
            I => \Lab_UT.didp.countrce1.un13_qPone_cascade_\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__17907\,
            I => \Lab_UT.didp.countrce1.q_5_2_cascade_\
        );

    \I__3607\ : InMux
    port map (
            O => \N__17904\,
            I => \N__17896\
        );

    \I__3606\ : InMux
    port map (
            O => \N__17903\,
            I => \N__17889\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17902\,
            I => \N__17889\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17901\,
            I => \N__17889\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17900\,
            I => \N__17886\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17899\,
            I => \N__17883\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__17896\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__17889\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__17886\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__17883\,
            I => \Lab_UT.di_Sones_2\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17874\,
            I => \N__17871\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__17871\,
            I => \Lab_UT.dispString.m49Z0Z_12\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__17868\,
            I => \Lab_UT.dispString.m49Z0Z_4_cascade_\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17865\,
            I => \N__17861\
        );

    \I__3593\ : InMux
    port map (
            O => \N__17864\,
            I => \N__17858\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__17861\,
            I => \N__17853\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__17858\,
            I => \N__17853\
        );

    \I__3590\ : Odrv12
    port map (
            O => \N__17853\,
            I => \Lab_UT.dispString.N_128_mux\
        );

    \I__3589\ : InMux
    port map (
            O => \N__17850\,
            I => \N__17847\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17842\
        );

    \I__3587\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17837\
        );

    \I__3586\ : InMux
    port map (
            O => \N__17845\,
            I => \N__17837\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__17842\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__17837\,
            I => \Lab_UT.di_AStens_2\
        );

    \I__3583\ : InMux
    port map (
            O => \N__17832\,
            I => \N__17829\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__17829\,
            I => \N__17825\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17828\,
            I => \N__17822\
        );

    \I__3580\ : Span4Mux_v
    port map (
            O => \N__17825\,
            I => \N__17818\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__17822\,
            I => \N__17815\
        );

    \I__3578\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17812\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__17818\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__17815\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__17812\,
            I => \Lab_UT.di_ASones_2\
        );

    \I__3574\ : InMux
    port map (
            O => \N__17805\,
            I => \N__17802\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__17802\,
            I => \N__17794\
        );

    \I__3572\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17791\
        );

    \I__3571\ : InMux
    port map (
            O => \N__17800\,
            I => \N__17782\
        );

    \I__3570\ : InMux
    port map (
            O => \N__17799\,
            I => \N__17782\
        );

    \I__3569\ : InMux
    port map (
            O => \N__17798\,
            I => \N__17782\
        );

    \I__3568\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17782\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__17794\,
            I => \N__17777\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__17791\,
            I => \N__17777\
        );

    \I__3565\ : LocalMux
    port map (
            O => \N__17782\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__17777\,
            I => \uu2.w_addr_displaying_0_repZ0Z1\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__17772\,
            I => \N__17769\
        );

    \I__3562\ : InMux
    port map (
            O => \N__17769\,
            I => \N__17766\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__17766\,
            I => \N__17763\
        );

    \I__3560\ : Odrv4
    port map (
            O => \N__17763\,
            I => \uu2.N_15\
        );

    \I__3559\ : InMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__17757\,
            I => \uu2.N_17\
        );

    \I__3557\ : CascadeMux
    port map (
            O => \N__17754\,
            I => \uu2.bitmap_pmux_25_i_m2_ns_1_cascade_\
        );

    \I__3556\ : CascadeMux
    port map (
            O => \N__17751\,
            I => \N__17748\
        );

    \I__3555\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17745\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__17745\,
            I => \N__17742\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__17742\,
            I => \uu2.N_49\
        );

    \I__3552\ : InMux
    port map (
            O => \N__17739\,
            I => \N__17736\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__17736\,
            I => \uu2.bitmapZ0Z_221\
        );

    \I__3550\ : InMux
    port map (
            O => \N__17733\,
            I => \N__17730\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__17730\,
            I => \uu2.bitmapZ0Z_93\
        );

    \I__3548\ : InMux
    port map (
            O => \N__17727\,
            I => \N__17724\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17724\,
            I => \uu2.N_13\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__17721\,
            I => \Lab_UT.didp.countrce1.un20_qPone_cascade_\
        );

    \I__3545\ : CascadeMux
    port map (
            O => \N__17718\,
            I => \Lab_UT.didp.countrce1.q_5_3_cascade_\
        );

    \I__3544\ : CascadeMux
    port map (
            O => \N__17715\,
            I => \N__17708\
        );

    \I__3543\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17705\
        );

    \I__3542\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17700\
        );

    \I__3541\ : InMux
    port map (
            O => \N__17712\,
            I => \N__17700\
        );

    \I__3540\ : InMux
    port map (
            O => \N__17711\,
            I => \N__17695\
        );

    \I__3539\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17695\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__17705\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__17700\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__17695\,
            I => \Lab_UT.di_Sones_3\
        );

    \I__3535\ : InMux
    port map (
            O => \N__17688\,
            I => \N__17682\
        );

    \I__3534\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17682\
        );

    \I__3533\ : LocalMux
    port map (
            O => \N__17682\,
            I => \uu2.w_addr_displaying_0_rep1_RNIDASJZ0\
        );

    \I__3532\ : CascadeMux
    port map (
            O => \N__17679\,
            I => \N__17676\
        );

    \I__3531\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17673\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__17673\,
            I => \uu2.w_addr_displaying_RNIR2PLZ0Z_8\
        );

    \I__3529\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17667\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__17667\,
            I => \uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1\
        );

    \I__3527\ : InMux
    port map (
            O => \N__17664\,
            I => \N__17661\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__17661\,
            I => \N__17658\
        );

    \I__3525\ : Odrv4
    port map (
            O => \N__17658\,
            I => \uu2.bitmap_pmux_29_0\
        );

    \I__3524\ : InMux
    port map (
            O => \N__17655\,
            I => \N__17650\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17654\,
            I => \N__17647\
        );

    \I__3522\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17644\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__17650\,
            I => \uu2.N_24_0\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__17647\,
            I => \uu2.N_24_0\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__17644\,
            I => \uu2.N_24_0\
        );

    \I__3518\ : InMux
    port map (
            O => \N__17637\,
            I => \N__17634\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__17634\,
            I => \uu2.w_addr_displaying_RNIU1AF7Z0Z_0\
        );

    \I__3516\ : InMux
    port map (
            O => \N__17631\,
            I => \N__17625\
        );

    \I__3515\ : InMux
    port map (
            O => \N__17630\,
            I => \N__17625\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17622\
        );

    \I__3513\ : Span4Mux_h
    port map (
            O => \N__17622\,
            I => \N__17619\
        );

    \I__3512\ : Span4Mux_v
    port map (
            O => \N__17619\,
            I => \N__17616\
        );

    \I__3511\ : Odrv4
    port map (
            O => \N__17616\,
            I => \Lab_UT.dictrl.m12Z0Z_2\
        );

    \I__3510\ : InMux
    port map (
            O => \N__17613\,
            I => \N__17610\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__17610\,
            I => \uu2.bitmapZ0Z_215\
        );

    \I__3508\ : CascadeMux
    port map (
            O => \N__17607\,
            I => \uu2.N_198_cascade_\
        );

    \I__3507\ : InMux
    port map (
            O => \N__17604\,
            I => \N__17601\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__17601\,
            I => \N__17598\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__17598\,
            I => \uu2.N_199\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__17595\,
            I => \uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_\
        );

    \I__3503\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17589\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__17589\,
            I => \uu2.N_196\
        );

    \I__3501\ : InMux
    port map (
            O => \N__17586\,
            I => \N__17583\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__17583\,
            I => \uu2.bitmap_pmux_27_i_m2_ns_1\
        );

    \I__3499\ : InMux
    port map (
            O => \N__17580\,
            I => \N__17577\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__17577\,
            I => \N__17574\
        );

    \I__3497\ : Span4Mux_s3_v
    port map (
            O => \N__17574\,
            I => \N__17571\
        );

    \I__3496\ : Odrv4
    port map (
            O => \N__17571\,
            I => \Lab_UT.dictrl.m53_d_1_1\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__17568\,
            I => \Lab_UT.dictrl.N_97_mux_3_cascade_\
        );

    \I__3494\ : InMux
    port map (
            O => \N__17565\,
            I => \N__17562\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__17562\,
            I => \uu2.bitmap_pmux_sn_N_42\
        );

    \I__3492\ : CascadeMux
    port map (
            O => \N__17559\,
            I => \N__17552\
        );

    \I__3491\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17548\
        );

    \I__3490\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17545\
        );

    \I__3489\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17540\
        );

    \I__3488\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17540\
        );

    \I__3487\ : InMux
    port map (
            O => \N__17552\,
            I => \N__17535\
        );

    \I__3486\ : InMux
    port map (
            O => \N__17551\,
            I => \N__17535\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__17548\,
            I => \N__17532\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__17545\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__17540\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__17535\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3481\ : Odrv12
    port map (
            O => \N__17532\,
            I => \uu2.w_addr_userZ0Z_1\
        );

    \I__3480\ : InMux
    port map (
            O => \N__17523\,
            I => \N__17519\
        );

    \I__3479\ : CascadeMux
    port map (
            O => \N__17522\,
            I => \N__17515\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__17519\,
            I => \N__17510\
        );

    \I__3477\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17507\
        );

    \I__3476\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17502\
        );

    \I__3475\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17502\
        );

    \I__3474\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17499\
        );

    \I__3473\ : Span4Mux_s0_v
    port map (
            O => \N__17510\,
            I => \N__17496\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__17507\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__17502\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__17499\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3469\ : Odrv4
    port map (
            O => \N__17496\,
            I => \uu2.w_addr_userZ0Z_2\
        );

    \I__3468\ : CascadeMux
    port map (
            O => \N__17487\,
            I => \uu2.un3_w_addr_user_4_cascade_\
        );

    \I__3467\ : InMux
    port map (
            O => \N__17484\,
            I => \N__17481\
        );

    \I__3466\ : LocalMux
    port map (
            O => \N__17481\,
            I => \N__17478\
        );

    \I__3465\ : Span4Mux_s1_v
    port map (
            O => \N__17478\,
            I => \N__17475\
        );

    \I__3464\ : Odrv4
    port map (
            O => \N__17475\,
            I => \uu2.un3_w_addr_user_5\
        );

    \I__3463\ : CascadeMux
    port map (
            O => \N__17472\,
            I => \N__17469\
        );

    \I__3462\ : InMux
    port map (
            O => \N__17469\,
            I => \N__17465\
        );

    \I__3461\ : InMux
    port map (
            O => \N__17468\,
            I => \N__17462\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__17465\,
            I => \N__17457\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__17462\,
            I => \N__17457\
        );

    \I__3458\ : IoSpan4Mux
    port map (
            O => \N__17457\,
            I => \N__17454\
        );

    \I__3457\ : Span4Mux_s0_v
    port map (
            O => \N__17454\,
            I => \N__17451\
        );

    \I__3456\ : Odrv4
    port map (
            O => \N__17451\,
            I => \uu2.un3_w_addr_user\
        );

    \I__3455\ : CEMux
    port map (
            O => \N__17448\,
            I => \N__17445\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__17445\,
            I => \N__17442\
        );

    \I__3453\ : Span4Mux_s0_v
    port map (
            O => \N__17442\,
            I => \N__17439\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__17439\,
            I => \N__17436\
        );

    \I__3451\ : Odrv4
    port map (
            O => \N__17436\,
            I => \uu2.un21_w_addr_displaying_0_0\
        );

    \I__3450\ : InMux
    port map (
            O => \N__17433\,
            I => \N__17430\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__17430\,
            I => \N__17427\
        );

    \I__3448\ : Span4Mux_s1_v
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__3447\ : Odrv4
    port map (
            O => \N__17424\,
            I => \uu2.bitmap_pmux_sn_N_33\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__17421\,
            I => \N__17416\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__17420\,
            I => \N__17410\
        );

    \I__3444\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17402\
        );

    \I__3443\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17402\
        );

    \I__3442\ : InMux
    port map (
            O => \N__17415\,
            I => \N__17402\
        );

    \I__3441\ : InMux
    port map (
            O => \N__17414\,
            I => \N__17393\
        );

    \I__3440\ : InMux
    port map (
            O => \N__17413\,
            I => \N__17393\
        );

    \I__3439\ : InMux
    port map (
            O => \N__17410\,
            I => \N__17393\
        );

    \I__3438\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17393\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__17402\,
            I => \N__17390\
        );

    \I__3436\ : LocalMux
    port map (
            O => \N__17393\,
            I => \uu2.w_addr_displayingZ1Z_4\
        );

    \I__3435\ : Odrv4
    port map (
            O => \N__17390\,
            I => \uu2.w_addr_displayingZ1Z_4\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__17385\,
            I => \uu2.bitmap_pmux_sn_N_33_cascade_\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__17382\,
            I => \N__17378\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__17381\,
            I => \N__17371\
        );

    \I__3431\ : InMux
    port map (
            O => \N__17378\,
            I => \N__17368\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \N__17363\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__17376\,
            I => \N__17360\
        );

    \I__3428\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17353\
        );

    \I__3427\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17353\
        );

    \I__3426\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17353\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__17368\,
            I => \N__17350\
        );

    \I__3424\ : InMux
    port map (
            O => \N__17367\,
            I => \N__17345\
        );

    \I__3423\ : InMux
    port map (
            O => \N__17366\,
            I => \N__17345\
        );

    \I__3422\ : InMux
    port map (
            O => \N__17363\,
            I => \N__17342\
        );

    \I__3421\ : InMux
    port map (
            O => \N__17360\,
            I => \N__17339\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__17353\,
            I => \N__17334\
        );

    \I__3419\ : Span4Mux_s1_v
    port map (
            O => \N__17350\,
            I => \N__17334\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__17345\,
            I => \N__17331\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__17342\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__17339\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3415\ : Odrv4
    port map (
            O => \N__17334\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3414\ : Odrv12
    port map (
            O => \N__17331\,
            I => \uu2.w_addr_displayingZ0Z_2\
        );

    \I__3413\ : InMux
    port map (
            O => \N__17322\,
            I => \N__17319\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__17319\,
            I => \N__17316\
        );

    \I__3411\ : Span4Mux_s1_v
    port map (
            O => \N__17316\,
            I => \N__17313\
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__17313\,
            I => \uu2.bitmap_pmux_sn_m15_0_1\
        );

    \I__3409\ : InMux
    port map (
            O => \N__17310\,
            I => \N__17307\
        );

    \I__3408\ : LocalMux
    port map (
            O => \N__17307\,
            I => \Lab_UT.dictrl.g1_1\
        );

    \I__3407\ : InMux
    port map (
            O => \N__17304\,
            I => \N__17301\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__17301\,
            I => \N__17298\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__17298\,
            I => \Lab_UT.dictrl.N_5\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__17295\,
            I => \Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_\
        );

    \I__3403\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17289\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17286\
        );

    \I__3401\ : Odrv4
    port map (
            O => \N__17286\,
            I => \Lab_UT.dictrl.N_9\
        );

    \I__3400\ : InMux
    port map (
            O => \N__17283\,
            I => \N__17280\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__17280\,
            I => \Lab_UT.dictrl.g2_1_3\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__17277\,
            I => \Lab_UT.dictrl.N_1462_3_cascade_\
        );

    \I__3397\ : InMux
    port map (
            O => \N__17274\,
            I => \N__17271\
        );

    \I__3396\ : LocalMux
    port map (
            O => \N__17271\,
            I => \Lab_UT.dictrl.N_1102_3\
        );

    \I__3395\ : InMux
    port map (
            O => \N__17268\,
            I => \N__17265\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__17265\,
            I => \Lab_UT.dictrl.N_1460_3\
        );

    \I__3393\ : InMux
    port map (
            O => \N__17262\,
            I => \N__17259\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__17259\,
            I => \N__17256\
        );

    \I__3391\ : Odrv12
    port map (
            O => \N__17256\,
            I => \Lab_UT.dictrl.N_6\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__17253\,
            I => \Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_\
        );

    \I__3389\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17247\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__17247\,
            I => \Lab_UT.dictrl.g0_i_m2_i_1\
        );

    \I__3387\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17241\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__17241\,
            I => \Lab_UT.dictrl.N_97_mux_1\
        );

    \I__3385\ : InMux
    port map (
            O => \N__17238\,
            I => \N__17235\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__17235\,
            I => \N__17232\
        );

    \I__3383\ : Odrv12
    port map (
            O => \N__17232\,
            I => \Lab_UT.dictrl.g0_i_a5_0_2\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__17229\,
            I => \N__17226\
        );

    \I__3381\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17223\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__17223\,
            I => \N__17220\
        );

    \I__3379\ : Odrv12
    port map (
            O => \N__17220\,
            I => \Lab_UT.dictrl.g2_2\
        );

    \I__3378\ : CascadeMux
    port map (
            O => \N__17217\,
            I => \Lab_UT.dictrl.g2_3_cascade_\
        );

    \I__3377\ : InMux
    port map (
            O => \N__17214\,
            I => \N__17211\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__17211\,
            I => \N__17208\
        );

    \I__3375\ : Odrv12
    port map (
            O => \N__17208\,
            I => \Lab_UT.dictrl.next_state_3_1\
        );

    \I__3374\ : InMux
    port map (
            O => \N__17205\,
            I => \N__17202\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__17202\,
            I => \N__17199\
        );

    \I__3372\ : Span4Mux_h
    port map (
            O => \N__17199\,
            I => \N__17196\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__17196\,
            I => \Lab_UT.dictrl.g0_12_a6_2_2\
        );

    \I__3370\ : InMux
    port map (
            O => \N__17193\,
            I => \N__17190\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__17190\,
            I => \N__17187\
        );

    \I__3368\ : Span4Mux_h
    port map (
            O => \N__17187\,
            I => \N__17184\
        );

    \I__3367\ : Odrv4
    port map (
            O => \N__17184\,
            I => \Lab_UT.dictrl.N_19\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__17181\,
            I => \Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_\
        );

    \I__3365\ : InMux
    port map (
            O => \N__17178\,
            I => \N__17175\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__17175\,
            I => \N__17172\
        );

    \I__3363\ : Span4Mux_h
    port map (
            O => \N__17172\,
            I => \N__17169\
        );

    \I__3362\ : Odrv4
    port map (
            O => \N__17169\,
            I => \Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3\
        );

    \I__3361\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17160\
        );

    \I__3360\ : InMux
    port map (
            O => \N__17165\,
            I => \N__17160\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__17160\,
            I => \N__17157\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__17157\,
            I => \N__17154\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__17154\,
            I => \Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2\
        );

    \I__3356\ : CascadeMux
    port map (
            O => \N__17151\,
            I => \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_\
        );

    \I__3355\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17133\
        );

    \I__3354\ : InMux
    port map (
            O => \N__17147\,
            I => \N__17133\
        );

    \I__3353\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17133\
        );

    \I__3352\ : InMux
    port map (
            O => \N__17145\,
            I => \N__17133\
        );

    \I__3351\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17133\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__17133\,
            I => \N__17130\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__17130\,
            I => \Lab_UT.dictrl.N_1792_0_0_0\
        );

    \I__3348\ : InMux
    port map (
            O => \N__17127\,
            I => \N__17124\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__17124\,
            I => \N__17121\
        );

    \I__3346\ : Odrv4
    port map (
            O => \N__17121\,
            I => \Lab_UT.dictrl.m53_d_1_5\
        );

    \I__3345\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17114\
        );

    \I__3344\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17108\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__17114\,
            I => \N__17104\
        );

    \I__3342\ : InMux
    port map (
            O => \N__17113\,
            I => \N__17097\
        );

    \I__3341\ : InMux
    port map (
            O => \N__17112\,
            I => \N__17097\
        );

    \I__3340\ : InMux
    port map (
            O => \N__17111\,
            I => \N__17097\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__17108\,
            I => \N__17090\
        );

    \I__3338\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17087\
        );

    \I__3337\ : Span4Mux_v
    port map (
            O => \N__17104\,
            I => \N__17082\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__17097\,
            I => \N__17082\
        );

    \I__3335\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17075\
        );

    \I__3334\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17075\
        );

    \I__3333\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17075\
        );

    \I__3332\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17072\
        );

    \I__3331\ : Span4Mux_s3_h
    port map (
            O => \N__17090\,
            I => \N__17069\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__17087\,
            I => \N__17066\
        );

    \I__3329\ : Span4Mux_h
    port map (
            O => \N__17082\,
            I => \N__17061\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__17075\,
            I => \N__17061\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__17072\,
            I => bu_rx_data_4_rep1
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__17069\,
            I => bu_rx_data_4_rep1
        );

    \I__3325\ : Odrv12
    port map (
            O => \N__17066\,
            I => bu_rx_data_4_rep1
        );

    \I__3324\ : Odrv4
    port map (
            O => \N__17061\,
            I => bu_rx_data_4_rep1
        );

    \I__3323\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17049\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__17049\,
            I => \Lab_UT.dictrl.N_40_0\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__17046\,
            I => \N__17042\
        );

    \I__3320\ : CascadeMux
    port map (
            O => \N__17045\,
            I => \N__17038\
        );

    \I__3319\ : InMux
    port map (
            O => \N__17042\,
            I => \N__17025\
        );

    \I__3318\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17025\
        );

    \I__3317\ : InMux
    port map (
            O => \N__17038\,
            I => \N__17025\
        );

    \I__3316\ : InMux
    port map (
            O => \N__17037\,
            I => \N__17025\
        );

    \I__3315\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17025\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__17022\
        );

    \I__3313\ : Span4Mux_h
    port map (
            O => \N__17022\,
            I => \N__17019\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__17019\,
            I => \Lab_UT.dictrl.N_23_1\
        );

    \I__3311\ : InMux
    port map (
            O => \N__17016\,
            I => \N__17001\
        );

    \I__3310\ : InMux
    port map (
            O => \N__17015\,
            I => \N__17001\
        );

    \I__3309\ : InMux
    port map (
            O => \N__17014\,
            I => \N__17001\
        );

    \I__3308\ : InMux
    port map (
            O => \N__17013\,
            I => \N__17001\
        );

    \I__3307\ : InMux
    port map (
            O => \N__17012\,
            I => \N__17001\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__17001\,
            I => \N__16998\
        );

    \I__3305\ : Span4Mux_h
    port map (
            O => \N__16998\,
            I => \N__16995\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__16995\,
            I => \G_17_i_0\
        );

    \I__3303\ : CascadeMux
    port map (
            O => \N__16992\,
            I => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__16989\,
            I => \N__16984\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__16988\,
            I => \N__16980\
        );

    \I__3300\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16965\
        );

    \I__3299\ : InMux
    port map (
            O => \N__16984\,
            I => \N__16965\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16983\,
            I => \N__16965\
        );

    \I__3297\ : InMux
    port map (
            O => \N__16980\,
            I => \N__16965\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16979\,
            I => \N__16965\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16978\,
            I => \N__16965\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16965\,
            I => \N__16962\
        );

    \I__3293\ : Odrv4
    port map (
            O => \N__16962\,
            I => \Lab_UT.dictrl.next_state_latmux_2_1\
        );

    \I__3292\ : CascadeMux
    port map (
            O => \N__16959\,
            I => \N__16956\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16956\,
            I => \N__16952\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16955\,
            I => \N__16948\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__16952\,
            I => \N__16945\
        );

    \I__3288\ : IoInMux
    port map (
            O => \N__16951\,
            I => \N__16941\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16948\,
            I => \N__16938\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__16945\,
            I => \N__16935\
        );

    \I__3285\ : SRMux
    port map (
            O => \N__16944\,
            I => \N__16932\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__16941\,
            I => \N__16929\
        );

    \I__3283\ : Span4Mux_v
    port map (
            O => \N__16938\,
            I => \N__16926\
        );

    \I__3282\ : Span4Mux_v
    port map (
            O => \N__16935\,
            I => \N__16919\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__16932\,
            I => \N__16919\
        );

    \I__3280\ : Span4Mux_s1_v
    port map (
            O => \N__16929\,
            I => \N__16919\
        );

    \I__3279\ : Span4Mux_v
    port map (
            O => \N__16926\,
            I => \N__16916\
        );

    \I__3278\ : Span4Mux_h
    port map (
            O => \N__16919\,
            I => \N__16913\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__16916\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__16913\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__16908\,
            I => \N__16905\
        );

    \I__3274\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16902\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__16902\,
            I => \Lab_UT.dictrl.next_state_0_3\
        );

    \I__3272\ : CEMux
    port map (
            O => \N__16899\,
            I => \N__16896\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__16896\,
            I => \N__16891\
        );

    \I__3270\ : CEMux
    port map (
            O => \N__16895\,
            I => \N__16888\
        );

    \I__3269\ : CEMux
    port map (
            O => \N__16894\,
            I => \N__16885\
        );

    \I__3268\ : Span4Mux_s3_v
    port map (
            O => \N__16891\,
            I => \N__16881\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__16888\,
            I => \N__16878\
        );

    \I__3266\ : LocalMux
    port map (
            O => \N__16885\,
            I => \N__16875\
        );

    \I__3265\ : CEMux
    port map (
            O => \N__16884\,
            I => \N__16872\
        );

    \I__3264\ : Odrv4
    port map (
            O => \N__16881\,
            I => \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\
        );

    \I__3263\ : Odrv12
    port map (
            O => \N__16878\,
            I => \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__16875\,
            I => \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16872\,
            I => \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__16863\,
            I => \N__16857\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__16862\,
            I => \N__16853\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__16861\,
            I => \N__16850\
        );

    \I__3257\ : InMux
    port map (
            O => \N__16860\,
            I => \N__16839\
        );

    \I__3256\ : InMux
    port map (
            O => \N__16857\,
            I => \N__16839\
        );

    \I__3255\ : InMux
    port map (
            O => \N__16856\,
            I => \N__16839\
        );

    \I__3254\ : InMux
    port map (
            O => \N__16853\,
            I => \N__16839\
        );

    \I__3253\ : InMux
    port map (
            O => \N__16850\,
            I => \N__16839\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__16839\,
            I => \Lab_UT.dictrl.G_17_i_a5_1_1\
        );

    \I__3251\ : InMux
    port map (
            O => \N__16836\,
            I => \N__16822\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16835\,
            I => \N__16822\
        );

    \I__3249\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16822\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16833\,
            I => \N__16819\
        );

    \I__3247\ : InMux
    port map (
            O => \N__16832\,
            I => \N__16812\
        );

    \I__3246\ : InMux
    port map (
            O => \N__16831\,
            I => \N__16812\
        );

    \I__3245\ : InMux
    port map (
            O => \N__16830\,
            I => \N__16812\
        );

    \I__3244\ : InMux
    port map (
            O => \N__16829\,
            I => \N__16809\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__16822\,
            I => \N__16806\
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__16819\,
            I => \N__16801\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__16812\,
            I => \N__16801\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__16809\,
            I => \N__16798\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__16806\,
            I => \N__16792\
        );

    \I__3238\ : Span4Mux_v
    port map (
            O => \N__16801\,
            I => \N__16789\
        );

    \I__3237\ : Span4Mux_h
    port map (
            O => \N__16798\,
            I => \N__16786\
        );

    \I__3236\ : InMux
    port map (
            O => \N__16797\,
            I => \N__16779\
        );

    \I__3235\ : InMux
    port map (
            O => \N__16796\,
            I => \N__16779\
        );

    \I__3234\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16779\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__16792\,
            I => \Lab_UT.dictrl.state_1_rep2\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__16789\,
            I => \Lab_UT.dictrl.state_1_rep2\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__16786\,
            I => \Lab_UT.dictrl.state_1_rep2\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__16779\,
            I => \Lab_UT.dictrl.state_1_rep2\
        );

    \I__3229\ : InMux
    port map (
            O => \N__16770\,
            I => \N__16767\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__16767\,
            I => \N__16764\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__16764\,
            I => \Lab_UT.dictrl.N_15_0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16758\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__16758\,
            I => \N__16755\
        );

    \I__3224\ : Span4Mux_h
    port map (
            O => \N__16755\,
            I => \N__16752\
        );

    \I__3223\ : Odrv4
    port map (
            O => \N__16752\,
            I => \Lab_UT.dictrl.g0_i_m2_0_1\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__16749\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_\
        );

    \I__3221\ : InMux
    port map (
            O => \N__16746\,
            I => \N__16743\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__16743\,
            I => \N__16740\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__16740\,
            I => \Lab_UT.dictrl.g0_i_m2_0_2\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__16737\,
            I => \Lab_UT.dictrl.next_state_0_0_2_cascade_\
        );

    \I__3217\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16730\
        );

    \I__3216\ : InMux
    port map (
            O => \N__16733\,
            I => \N__16727\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__16730\,
            I => \N__16721\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__16727\,
            I => \N__16721\
        );

    \I__3213\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16716\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__16721\,
            I => \N__16713\
        );

    \I__3211\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16710\
        );

    \I__3210\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16707\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__16716\,
            I => \N__16704\
        );

    \I__3208\ : Span4Mux_v
    port map (
            O => \N__16713\,
            I => \N__16697\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__16710\,
            I => \N__16697\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__16707\,
            I => \N__16697\
        );

    \I__3205\ : Span4Mux_s3_v
    port map (
            O => \N__16704\,
            I => \N__16694\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__16697\,
            I => \N__16690\
        );

    \I__3203\ : Span4Mux_h
    port map (
            O => \N__16694\,
            I => \N__16687\
        );

    \I__3202\ : IoInMux
    port map (
            O => \N__16693\,
            I => \N__16684\
        );

    \I__3201\ : Odrv4
    port map (
            O => \N__16690\,
            I => rst
        );

    \I__3200\ : Odrv4
    port map (
            O => \N__16687\,
            I => rst
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16684\,
            I => rst
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__16677\,
            I => \N__16674\
        );

    \I__3197\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16671\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__16671\,
            I => \N__16668\
        );

    \I__3195\ : Odrv4
    port map (
            O => \N__16668\,
            I => \Lab_UT.didp.countrce4.un13_qPone\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16662\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__16662\,
            I => \N__16659\
        );

    \I__3192\ : Span4Mux_v
    port map (
            O => \N__16659\,
            I => \N__16656\
        );

    \I__3191\ : Span4Mux_h
    port map (
            O => \N__16656\,
            I => \N__16652\
        );

    \I__3190\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16649\
        );

    \I__3189\ : Odrv4
    port map (
            O => \N__16652\,
            I => \Lab_UT.LdAMtens\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__16649\,
            I => \Lab_UT.LdAMtens\
        );

    \I__3187\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16638\
        );

    \I__3186\ : InMux
    port map (
            O => \N__16643\,
            I => \N__16638\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__16638\,
            I => \Lab_UT.LdAMones\
        );

    \I__3184\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16632\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__16632\,
            I => \N__16629\
        );

    \I__3182\ : Span4Mux_s3_h
    port map (
            O => \N__16629\,
            I => \N__16625\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__16628\,
            I => \N__16622\
        );

    \I__3180\ : Span4Mux_h
    port map (
            O => \N__16625\,
            I => \N__16619\
        );

    \I__3179\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16616\
        );

    \I__3178\ : Odrv4
    port map (
            O => \N__16619\,
            I => \Lab_UT.LdAStens\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__16616\,
            I => \Lab_UT.LdAStens\
        );

    \I__3176\ : InMux
    port map (
            O => \N__16611\,
            I => \N__16608\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__16608\,
            I => \N__16605\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__16605\,
            I => \Lab_UT.dictrl.N_1460_2\
        );

    \I__3173\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16594\
        );

    \I__3172\ : InMux
    port map (
            O => \N__16601\,
            I => \N__16594\
        );

    \I__3171\ : InMux
    port map (
            O => \N__16600\,
            I => \N__16589\
        );

    \I__3170\ : InMux
    port map (
            O => \N__16599\,
            I => \N__16586\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16583\
        );

    \I__3168\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16578\
        );

    \I__3167\ : InMux
    port map (
            O => \N__16592\,
            I => \N__16578\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16575\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__16586\,
            I => \N__16570\
        );

    \I__3164\ : Span4Mux_s2_v
    port map (
            O => \N__16583\,
            I => \N__16570\
        );

    \I__3163\ : LocalMux
    port map (
            O => \N__16578\,
            I => \N__16567\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__16575\,
            I => \N__16562\
        );

    \I__3161\ : Span4Mux_v
    port map (
            O => \N__16570\,
            I => \N__16562\
        );

    \I__3160\ : Odrv12
    port map (
            O => \N__16567\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__3159\ : Odrv4
    port map (
            O => \N__16562\,
            I => \Lab_UT.dictrl.state_fast_0\
        );

    \I__3158\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16554\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__16554\,
            I => \N__16551\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__16551\,
            I => \Lab_UT.dispString.m49Z0Z_0\
        );

    \I__3155\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16545\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__16545\,
            I => \Lab_UT.dispString.m49Z0Z_1\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__16542\,
            I => \Lab_UT.dispString.m49Z0Z_3_cascade_\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__16539\,
            I => \Lab_UT.loadalarm_0_cascade_\
        );

    \I__3151\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16517\
        );

    \I__3150\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16517\
        );

    \I__3149\ : InMux
    port map (
            O => \N__16534\,
            I => \N__16517\
        );

    \I__3148\ : InMux
    port map (
            O => \N__16533\,
            I => \N__16517\
        );

    \I__3147\ : InMux
    port map (
            O => \N__16532\,
            I => \N__16517\
        );

    \I__3146\ : InMux
    port map (
            O => \N__16531\,
            I => \N__16517\
        );

    \I__3145\ : InMux
    port map (
            O => \N__16530\,
            I => \N__16514\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__16517\,
            I => \N__16511\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__16514\,
            I => \N__16508\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__16511\,
            I => \N__16505\
        );

    \I__3141\ : Odrv12
    port map (
            O => \N__16508\,
            I => \Lab_UT.min2_0\
        );

    \I__3140\ : Odrv4
    port map (
            O => \N__16505\,
            I => \Lab_UT.min2_0\
        );

    \I__3139\ : CascadeMux
    port map (
            O => \N__16500\,
            I => \N__16497\
        );

    \I__3138\ : InMux
    port map (
            O => \N__16497\,
            I => \N__16494\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__16494\,
            I => \N__16491\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__16491\,
            I => \N__16486\
        );

    \I__3135\ : InMux
    port map (
            O => \N__16490\,
            I => \N__16481\
        );

    \I__3134\ : InMux
    port map (
            O => \N__16489\,
            I => \N__16481\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__16486\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__16481\,
            I => \Lab_UT.di_AMones_0\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__16476\,
            I => \N__16472\
        );

    \I__3130\ : InMux
    port map (
            O => \N__16475\,
            I => \N__16468\
        );

    \I__3129\ : InMux
    port map (
            O => \N__16472\,
            I => \N__16465\
        );

    \I__3128\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16462\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__16468\,
            I => \N__16457\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__16465\,
            I => \N__16457\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__16462\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__3124\ : Odrv4
    port map (
            O => \N__16457\,
            I => \Lab_UT.di_AMtens_0\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__16452\,
            I => \Lab_UT.dictrl.g0_12_a6_1_3_cascade_\
        );

    \I__3122\ : InMux
    port map (
            O => \N__16449\,
            I => \N__16446\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16443\
        );

    \I__3120\ : Odrv4
    port map (
            O => \N__16443\,
            I => \Lab_UT.dictrl.N_18\
        );

    \I__3119\ : CascadeMux
    port map (
            O => \N__16440\,
            I => \N__16437\
        );

    \I__3118\ : InMux
    port map (
            O => \N__16437\,
            I => \N__16434\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__16434\,
            I => \N__16431\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__16431\,
            I => \N__16428\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__16428\,
            I => \Lab_UT.dictrl.m35_0\
        );

    \I__3114\ : InMux
    port map (
            O => \N__16425\,
            I => \N__16419\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__16424\,
            I => \N__16415\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__16423\,
            I => \N__16412\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__16422\,
            I => \N__16409\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__16419\,
            I => \N__16404\
        );

    \I__3109\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16391\
        );

    \I__3108\ : InMux
    port map (
            O => \N__16415\,
            I => \N__16391\
        );

    \I__3107\ : InMux
    port map (
            O => \N__16412\,
            I => \N__16391\
        );

    \I__3106\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16391\
        );

    \I__3105\ : InMux
    port map (
            O => \N__16408\,
            I => \N__16391\
        );

    \I__3104\ : InMux
    port map (
            O => \N__16407\,
            I => \N__16391\
        );

    \I__3103\ : Span4Mux_s1_v
    port map (
            O => \N__16404\,
            I => \N__16386\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__16391\,
            I => \N__16386\
        );

    \I__3101\ : Odrv4
    port map (
            O => \N__16386\,
            I => \Lab_UT.min2_1\
        );

    \I__3100\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16380\
        );

    \I__3099\ : LocalMux
    port map (
            O => \N__16380\,
            I => \N__16371\
        );

    \I__3098\ : InMux
    port map (
            O => \N__16379\,
            I => \N__16358\
        );

    \I__3097\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16358\
        );

    \I__3096\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16358\
        );

    \I__3095\ : InMux
    port map (
            O => \N__16376\,
            I => \N__16358\
        );

    \I__3094\ : InMux
    port map (
            O => \N__16375\,
            I => \N__16358\
        );

    \I__3093\ : InMux
    port map (
            O => \N__16374\,
            I => \N__16358\
        );

    \I__3092\ : Span4Mux_h
    port map (
            O => \N__16371\,
            I => \N__16353\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__16358\,
            I => \N__16353\
        );

    \I__3090\ : Span4Mux_v
    port map (
            O => \N__16353\,
            I => \N__16350\
        );

    \I__3089\ : Odrv4
    port map (
            O => \N__16350\,
            I => \Lab_UT.min2_2\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__16347\,
            I => \N__16344\
        );

    \I__3087\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16341\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__16341\,
            I => \N__16338\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__16338\,
            I => \N__16333\
        );

    \I__3084\ : InMux
    port map (
            O => \N__16337\,
            I => \N__16328\
        );

    \I__3083\ : InMux
    port map (
            O => \N__16336\,
            I => \N__16328\
        );

    \I__3082\ : Odrv4
    port map (
            O => \N__16333\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__16328\,
            I => \Lab_UT.di_AStens_3\
        );

    \I__3080\ : CEMux
    port map (
            O => \N__16323\,
            I => \N__16320\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__16320\,
            I => \N__16317\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__16317\,
            I => \N__16314\
        );

    \I__3077\ : Odrv4
    port map (
            O => \N__16314\,
            I => \Lab_UT.didp.regrce2.LdAStens_0\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__16311\,
            I => \Lab_UT.didp.countrce4.q_5_2_cascade_\
        );

    \I__3075\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16304\
        );

    \I__3074\ : InMux
    port map (
            O => \N__16307\,
            I => \N__16300\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__16304\,
            I => \N__16297\
        );

    \I__3072\ : InMux
    port map (
            O => \N__16303\,
            I => \N__16294\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__16300\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3070\ : Odrv4
    port map (
            O => \N__16297\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__16294\,
            I => \Lab_UT.di_AMtens_2\
        );

    \I__3068\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16283\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__16286\,
            I => \N__16279\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__16283\,
            I => \N__16276\
        );

    \I__3065\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16273\
        );

    \I__3064\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16270\
        );

    \I__3063\ : Span4Mux_v
    port map (
            O => \N__16276\,
            I => \N__16267\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__16273\,
            I => \N__16264\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16261\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__16267\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__16264\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__16261\,
            I => \Lab_UT.di_AMtens_1\
        );

    \I__3057\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16246\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__16253\,
            I => \N__16243\
        );

    \I__3055\ : InMux
    port map (
            O => \N__16252\,
            I => \N__16235\
        );

    \I__3054\ : InMux
    port map (
            O => \N__16251\,
            I => \N__16232\
        );

    \I__3053\ : InMux
    port map (
            O => \N__16250\,
            I => \N__16229\
        );

    \I__3052\ : InMux
    port map (
            O => \N__16249\,
            I => \N__16226\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__16246\,
            I => \N__16223\
        );

    \I__3050\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16214\
        );

    \I__3049\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16214\
        );

    \I__3048\ : InMux
    port map (
            O => \N__16241\,
            I => \N__16214\
        );

    \I__3047\ : InMux
    port map (
            O => \N__16240\,
            I => \N__16214\
        );

    \I__3046\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16209\
        );

    \I__3045\ : InMux
    port map (
            O => \N__16238\,
            I => \N__16209\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__16235\,
            I => \N__16198\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__16232\,
            I => \N__16198\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__16229\,
            I => \N__16198\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__16226\,
            I => \N__16198\
        );

    \I__3040\ : Span12Mux_s11_h
    port map (
            O => \N__16223\,
            I => \N__16198\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__16214\,
            I => \buart__rx_startbit\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__16209\,
            I => \buart__rx_startbit\
        );

    \I__3037\ : Odrv12
    port map (
            O => \N__16198\,
            I => \buart__rx_startbit\
        );

    \I__3036\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16188\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__16188\,
            I => \N__16185\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__16185\,
            I => \N__16182\
        );

    \I__3033\ : Span4Mux_v
    port map (
            O => \N__16182\,
            I => \N__16178\
        );

    \I__3032\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16175\
        );

    \I__3031\ : Span4Mux_h
    port map (
            O => \N__16178\,
            I => \N__16170\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__16175\,
            I => \N__16167\
        );

    \I__3029\ : InMux
    port map (
            O => \N__16174\,
            I => \N__16164\
        );

    \I__3028\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16161\
        );

    \I__3027\ : Odrv4
    port map (
            O => \N__16170\,
            I => \buart__rx_N_27_0_i\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__16167\,
            I => \buart__rx_N_27_0_i\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__16164\,
            I => \buart__rx_N_27_0_i\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__16161\,
            I => \buart__rx_N_27_0_i\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__16152\,
            I => \N__16149\
        );

    \I__3022\ : InMux
    port map (
            O => \N__16149\,
            I => \N__16146\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__16146\,
            I => \N__16143\
        );

    \I__3020\ : Span4Mux_h
    port map (
            O => \N__16143\,
            I => \N__16140\
        );

    \I__3019\ : Span4Mux_v
    port map (
            O => \N__16140\,
            I => \N__16137\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__16137\,
            I => \N__16134\
        );

    \I__3017\ : Odrv4
    port map (
            O => \N__16134\,
            I => \buart.Z_rx.bitcount_cry_1_THRU_CO\
        );

    \I__3016\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16125\
        );

    \I__3015\ : InMux
    port map (
            O => \N__16130\,
            I => \N__16122\
        );

    \I__3014\ : InMux
    port map (
            O => \N__16129\,
            I => \N__16117\
        );

    \I__3013\ : InMux
    port map (
            O => \N__16128\,
            I => \N__16117\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__16125\,
            I => \N__16114\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__16122\,
            I => \N__16109\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__16117\,
            I => \N__16109\
        );

    \I__3009\ : Span4Mux_v
    port map (
            O => \N__16114\,
            I => \N__16104\
        );

    \I__3008\ : Span4Mux_v
    port map (
            O => \N__16109\,
            I => \N__16104\
        );

    \I__3007\ : Span4Mux_h
    port map (
            O => \N__16104\,
            I => \N__16100\
        );

    \I__3006\ : InMux
    port map (
            O => \N__16103\,
            I => \N__16097\
        );

    \I__3005\ : Span4Mux_v
    port map (
            O => \N__16100\,
            I => \N__16094\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__16097\,
            I => \buart__rx_bitcount_2\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__16094\,
            I => \buart__rx_bitcount_2\
        );

    \I__3002\ : CEMux
    port map (
            O => \N__16089\,
            I => \N__16086\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__16086\,
            I => \N__16082\
        );

    \I__3000\ : CEMux
    port map (
            O => \N__16085\,
            I => \N__16078\
        );

    \I__2999\ : Sp12to4
    port map (
            O => \N__16082\,
            I => \N__16074\
        );

    \I__2998\ : CEMux
    port map (
            O => \N__16081\,
            I => \N__16071\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16068\
        );

    \I__2996\ : CEMux
    port map (
            O => \N__16077\,
            I => \N__16065\
        );

    \I__2995\ : Span12Mux_s9_v
    port map (
            O => \N__16074\,
            I => \N__16062\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__16071\,
            I => \N__16059\
        );

    \I__2993\ : Span4Mux_v
    port map (
            O => \N__16068\,
            I => \N__16056\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16053\
        );

    \I__2991\ : Odrv12
    port map (
            O => \N__16062\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2990\ : Odrv4
    port map (
            O => \N__16059\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2989\ : Odrv4
    port map (
            O => \N__16056\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__16053\,
            I => \buart.Z_rx.bitcounte_0_0\
        );

    \I__2987\ : InMux
    port map (
            O => \N__16044\,
            I => \N__16041\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__16041\,
            I => \uu2.bitmapZ0Z_75\
        );

    \I__2985\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16035\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__16035\,
            I => \uu2.bitmapZ0Z_72\
        );

    \I__2983\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16029\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__16029\,
            I => \N__16026\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__16026\,
            I => \uu2.vram_rd_clk_detZ0Z_1\
        );

    \I__2980\ : InMux
    port map (
            O => \N__16023\,
            I => \N__16019\
        );

    \I__2979\ : InMux
    port map (
            O => \N__16022\,
            I => \N__16016\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__16019\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__16016\,
            I => \uu2.vram_rd_clk_detZ0Z_0\
        );

    \I__2976\ : CEMux
    port map (
            O => \N__16011\,
            I => \N__16008\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__16008\,
            I => \N__16005\
        );

    \I__2974\ : Span4Mux_s3_h
    port map (
            O => \N__16005\,
            I => \N__16002\
        );

    \I__2973\ : Span4Mux_h
    port map (
            O => \N__16002\,
            I => \N__15999\
        );

    \I__2972\ : Odrv4
    port map (
            O => \N__15999\,
            I => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15993\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__15993\,
            I => \N__15990\
        );

    \I__2969\ : Span4Mux_h
    port map (
            O => \N__15990\,
            I => \N__15985\
        );

    \I__2968\ : InMux
    port map (
            O => \N__15989\,
            I => \N__15980\
        );

    \I__2967\ : InMux
    port map (
            O => \N__15988\,
            I => \N__15980\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__15985\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__15980\,
            I => \Lab_UT.di_ASones_3\
        );

    \I__2964\ : CascadeMux
    port map (
            O => \N__15975\,
            I => \uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15968\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__15971\,
            I => \N__15965\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15968\,
            I => \N__15957\
        );

    \I__2960\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15950\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15950\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15963\,
            I => \N__15950\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15962\,
            I => \N__15943\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15961\,
            I => \N__15943\
        );

    \I__2955\ : InMux
    port map (
            O => \N__15960\,
            I => \N__15943\
        );

    \I__2954\ : Span4Mux_s3_v
    port map (
            O => \N__15957\,
            I => \N__15940\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__15950\,
            I => \N__15935\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15943\,
            I => \N__15935\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__15940\,
            I => \Lab_UT.min1_2\
        );

    \I__2950\ : Odrv12
    port map (
            O => \N__15935\,
            I => \Lab_UT.min1_2\
        );

    \I__2949\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15926\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__15929\,
            I => \N__15919\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__15926\,
            I => \N__15915\
        );

    \I__2946\ : InMux
    port map (
            O => \N__15925\,
            I => \N__15908\
        );

    \I__2945\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15908\
        );

    \I__2944\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15908\
        );

    \I__2943\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15901\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15901\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15901\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__15915\,
            I => \N__15898\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__15908\,
            I => \N__15895\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__15901\,
            I => \N__15892\
        );

    \I__2937\ : Odrv4
    port map (
            O => \N__15898\,
            I => \Lab_UT.min1_1\
        );

    \I__2936\ : Odrv12
    port map (
            O => \N__15895\,
            I => \Lab_UT.min1_1\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__15892\,
            I => \Lab_UT.min1_1\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__15885\,
            I => \N__15882\
        );

    \I__2933\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15875\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__15881\,
            I => \N__15871\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \N__15868\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__15879\,
            I => \N__15865\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__15878\,
            I => \N__15861\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__15875\,
            I => \N__15858\
        );

    \I__2927\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15851\
        );

    \I__2926\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15851\
        );

    \I__2925\ : InMux
    port map (
            O => \N__15868\,
            I => \N__15851\
        );

    \I__2924\ : InMux
    port map (
            O => \N__15865\,
            I => \N__15844\
        );

    \I__2923\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15844\
        );

    \I__2922\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15844\
        );

    \I__2921\ : Span4Mux_h
    port map (
            O => \N__15858\,
            I => \N__15839\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__15851\,
            I => \N__15839\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__15844\,
            I => \N__15836\
        );

    \I__2918\ : Odrv4
    port map (
            O => \N__15839\,
            I => \Lab_UT.min1_3\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__15836\,
            I => \Lab_UT.min1_3\
        );

    \I__2916\ : InMux
    port map (
            O => \N__15831\,
            I => \N__15828\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__15828\,
            I => \N__15819\
        );

    \I__2914\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15812\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15812\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15812\
        );

    \I__2911\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15805\
        );

    \I__2910\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15805\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15805\
        );

    \I__2908\ : Span4Mux_s3_v
    port map (
            O => \N__15819\,
            I => \N__15802\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__15812\,
            I => \N__15799\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15805\,
            I => \N__15796\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__15802\,
            I => \Lab_UT.min1_0\
        );

    \I__2904\ : Odrv12
    port map (
            O => \N__15799\,
            I => \Lab_UT.min1_0\
        );

    \I__2903\ : Odrv4
    port map (
            O => \N__15796\,
            I => \Lab_UT.min1_0\
        );

    \I__2902\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15786\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__15786\,
            I => \uu2.bitmapZ0Z_69\
        );

    \I__2900\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15780\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__15780\,
            I => \uu2.bitmapZ0Z_197\
        );

    \I__2898\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15757\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15757\
        );

    \I__2896\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15757\
        );

    \I__2895\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15757\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15757\
        );

    \I__2893\ : InMux
    port map (
            O => \N__15772\,
            I => \N__15750\
        );

    \I__2892\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15750\
        );

    \I__2891\ : InMux
    port map (
            O => \N__15770\,
            I => \N__15750\
        );

    \I__2890\ : InMux
    port map (
            O => \N__15769\,
            I => \N__15745\
        );

    \I__2889\ : InMux
    port map (
            O => \N__15768\,
            I => \N__15745\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__15757\,
            I => \N__15742\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__15750\,
            I => \N__15737\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__15745\,
            I => \N__15737\
        );

    \I__2885\ : Odrv4
    port map (
            O => \N__15742\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__15737\,
            I => \uu2.un4_w_user_data_rdyZ0Z_0\
        );

    \I__2883\ : InMux
    port map (
            O => \N__15732\,
            I => \N__15729\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__15729\,
            I => \uu2.bitmap_pmux_sn_N_65\
        );

    \I__2881\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15723\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__15723\,
            I => \uu2.N_54\
        );

    \I__2879\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15717\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__15717\,
            I => \uu2.N_53\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15714\,
            I => \N__15711\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__15711\,
            I => \N__15708\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__15708\,
            I => \Lab_UT.dictrl.m53_d_1_3\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__15705\,
            I => \Lab_UT.dictrl.N_97_mux_5_cascade_\
        );

    \I__2873\ : InMux
    port map (
            O => \N__15702\,
            I => \N__15697\
        );

    \I__2872\ : InMux
    port map (
            O => \N__15701\,
            I => \N__15694\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__15700\,
            I => \N__15689\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__15697\,
            I => \N__15684\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__15694\,
            I => \N__15684\
        );

    \I__2868\ : InMux
    port map (
            O => \N__15693\,
            I => \N__15681\
        );

    \I__2867\ : InMux
    port map (
            O => \N__15692\,
            I => \N__15676\
        );

    \I__2866\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15676\
        );

    \I__2865\ : Span4Mux_s1_v
    port map (
            O => \N__15684\,
            I => \N__15673\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__15681\,
            I => \Lab_UT.dictrl.N_40\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__15676\,
            I => \Lab_UT.dictrl.N_40\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__15673\,
            I => \Lab_UT.dictrl.N_40\
        );

    \I__2861\ : InMux
    port map (
            O => \N__15666\,
            I => \N__15662\
        );

    \I__2860\ : InMux
    port map (
            O => \N__15665\,
            I => \N__15659\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__15662\,
            I => \N__15656\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__15659\,
            I => \Lab_UT.dictrl.N_62\
        );

    \I__2857\ : Odrv12
    port map (
            O => \N__15656\,
            I => \Lab_UT.dictrl.N_62\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__15651\,
            I => \Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_\
        );

    \I__2855\ : InMux
    port map (
            O => \N__15648\,
            I => \N__15645\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__15645\,
            I => \Lab_UT.dictrl.next_state_RNO_1Z0Z_2\
        );

    \I__2853\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15639\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__15639\,
            I => \Lab_UT.dictrl.next_state_RNO_0Z0Z_2\
        );

    \I__2851\ : InMux
    port map (
            O => \N__15636\,
            I => \N__15633\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__15633\,
            I => \N__15620\
        );

    \I__2849\ : InMux
    port map (
            O => \N__15632\,
            I => \N__15615\
        );

    \I__2848\ : InMux
    port map (
            O => \N__15631\,
            I => \N__15615\
        );

    \I__2847\ : InMux
    port map (
            O => \N__15630\,
            I => \N__15608\
        );

    \I__2846\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15608\
        );

    \I__2845\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15608\
        );

    \I__2844\ : InMux
    port map (
            O => \N__15627\,
            I => \N__15603\
        );

    \I__2843\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15598\
        );

    \I__2842\ : InMux
    port map (
            O => \N__15625\,
            I => \N__15598\
        );

    \I__2841\ : InMux
    port map (
            O => \N__15624\,
            I => \N__15595\
        );

    \I__2840\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15592\
        );

    \I__2839\ : Span4Mux_h
    port map (
            O => \N__15620\,
            I => \N__15587\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__15615\,
            I => \N__15587\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__15608\,
            I => \N__15584\
        );

    \I__2836\ : InMux
    port map (
            O => \N__15607\,
            I => \N__15581\
        );

    \I__2835\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15578\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__15603\,
            I => \N__15575\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__15598\,
            I => \N__15564\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__15595\,
            I => \N__15564\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__15592\,
            I => \N__15564\
        );

    \I__2830\ : Sp12to4
    port map (
            O => \N__15587\,
            I => \N__15564\
        );

    \I__2829\ : Sp12to4
    port map (
            O => \N__15584\,
            I => \N__15564\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__15581\,
            I => \N__15561\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__15578\,
            I => \N__15558\
        );

    \I__2826\ : Span12Mux_s5_h
    port map (
            O => \N__15575\,
            I => \N__15553\
        );

    \I__2825\ : Span12Mux_s6_v
    port map (
            O => \N__15564\,
            I => \N__15553\
        );

    \I__2824\ : Span4Mux_s3_v
    port map (
            O => \N__15561\,
            I => \N__15548\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__15558\,
            I => \N__15548\
        );

    \I__2822\ : Odrv12
    port map (
            O => \N__15553\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__15548\,
            I => \Lab_UT.dictrl.state_3_rep1\
        );

    \I__2820\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__15540\,
            I => \N__15536\
        );

    \I__2818\ : InMux
    port map (
            O => \N__15539\,
            I => \N__15533\
        );

    \I__2817\ : Odrv4
    port map (
            O => \N__15536\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__15533\,
            I => \Lab_UT.dictrl.next_state_0_2\
        );

    \I__2815\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15525\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__15525\,
            I => \N__15522\
        );

    \I__2813\ : Span4Mux_h
    port map (
            O => \N__15522\,
            I => \N__15519\
        );

    \I__2812\ : Odrv4
    port map (
            O => \N__15519\,
            I => \Lab_UT.dictrl.next_state_RNINV3PZ0Z_2\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15510\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__15515\,
            I => \N__15507\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__15514\,
            I => \N__15501\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__15513\,
            I => \N__15498\
        );

    \I__2807\ : InMux
    port map (
            O => \N__15510\,
            I => \N__15495\
        );

    \I__2806\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15482\
        );

    \I__2805\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15482\
        );

    \I__2804\ : InMux
    port map (
            O => \N__15505\,
            I => \N__15482\
        );

    \I__2803\ : InMux
    port map (
            O => \N__15504\,
            I => \N__15482\
        );

    \I__2802\ : InMux
    port map (
            O => \N__15501\,
            I => \N__15482\
        );

    \I__2801\ : InMux
    port map (
            O => \N__15498\,
            I => \N__15482\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15495\,
            I => \N__15477\
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__15482\,
            I => \N__15477\
        );

    \I__2798\ : Span4Mux_s2_v
    port map (
            O => \N__15477\,
            I => \N__15474\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__15474\,
            I => \Lab_UT.min2_3\
        );

    \I__2796\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15468\,
            I => \uu2.bitmapZ0Z_203\
        );

    \I__2794\ : InMux
    port map (
            O => \N__15465\,
            I => \N__15462\
        );

    \I__2793\ : LocalMux
    port map (
            O => \N__15462\,
            I => \N__15459\
        );

    \I__2792\ : Odrv4
    port map (
            O => \N__15459\,
            I => \uu2.bitmapZ0Z_200\
        );

    \I__2791\ : InMux
    port map (
            O => \N__15456\,
            I => \N__15453\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__15453\,
            I => \N__15449\
        );

    \I__2789\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15446\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__15449\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__15446\,
            I => \Lab_UT.dictrl.next_state_0_0\
        );

    \I__2786\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__15438\,
            I => \Lab_UT.dictrl.N_8\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__15435\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_\
        );

    \I__2783\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15429\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__15429\,
            I => \Lab_UT.dictrl.N_20_0\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__15426\,
            I => \Lab_UT.dictrl.N_18_0_cascade_\
        );

    \I__2780\ : CascadeMux
    port map (
            O => \N__15423\,
            I => \N__15418\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \N__15415\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15421\,
            I => \N__15401\
        );

    \I__2777\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15401\
        );

    \I__2776\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15401\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15401\
        );

    \I__2774\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15390\
        );

    \I__2773\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15390\
        );

    \I__2772\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15390\
        );

    \I__2771\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15390\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15401\,
            I => \N__15387\
        );

    \I__2769\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15382\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15382\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__15390\,
            I => \N__15377\
        );

    \I__2766\ : Span4Mux_s2_v
    port map (
            O => \N__15387\,
            I => \N__15377\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15382\,
            I => \N__15374\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__15377\,
            I => \N__15371\
        );

    \I__2763\ : Odrv12
    port map (
            O => \N__15374\,
            I => \Lab_UT.dictrl.state_fast_3\
        );

    \I__2762\ : Odrv4
    port map (
            O => \N__15371\,
            I => \Lab_UT.dictrl.state_fast_3\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15361\
        );

    \I__2760\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15356\
        );

    \I__2759\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15356\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15361\,
            I => \N__15353\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__15356\,
            I => \N__15348\
        );

    \I__2756\ : Span4Mux_h
    port map (
            O => \N__15353\,
            I => \N__15348\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__15348\,
            I => \N__15345\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__15345\,
            I => \Lab_UT.dictrl.state_fast_2\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__15342\,
            I => \N__15337\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__15341\,
            I => \N__15333\
        );

    \I__2751\ : CascadeMux
    port map (
            O => \N__15340\,
            I => \N__15330\
        );

    \I__2750\ : InMux
    port map (
            O => \N__15337\,
            I => \N__15325\
        );

    \I__2749\ : InMux
    port map (
            O => \N__15336\,
            I => \N__15325\
        );

    \I__2748\ : InMux
    port map (
            O => \N__15333\,
            I => \N__15320\
        );

    \I__2747\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15320\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__15325\,
            I => \N__15317\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__15320\,
            I => \N__15314\
        );

    \I__2744\ : Odrv4
    port map (
            O => \N__15317\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__15314\,
            I => \Lab_UT.dictrl.state_1_rep1\
        );

    \I__2742\ : InMux
    port map (
            O => \N__15309\,
            I => \N__15306\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__15306\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_3_2\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__15303\,
            I => \N__15300\
        );

    \I__2739\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15297\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__15297\,
            I => \Lab_UT.dictrl.N_11_1\
        );

    \I__2737\ : InMux
    port map (
            O => \N__15294\,
            I => \N__15291\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__15291\,
            I => \N__15288\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__15288\,
            I => \N__15285\
        );

    \I__2734\ : Odrv4
    port map (
            O => \N__15285\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_4_6\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__15282\,
            I => \Lab_UT.dictrl.N_22_0_cascade_\
        );

    \I__2732\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15276\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__15276\,
            I => \N__15273\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__15273\,
            I => \N__15270\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__15270\,
            I => \Lab_UT.dictrl.g0_i_m2_0_a7_4_7\
        );

    \I__2728\ : InMux
    port map (
            O => \N__15267\,
            I => \N__15264\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__15264\,
            I => \N__15261\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__15261\,
            I => \Lab_UT.dictrl.N_1110_1\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__15258\,
            I => \N__15254\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__15257\,
            I => \N__15250\
        );

    \I__2723\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15237\
        );

    \I__2722\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15237\
        );

    \I__2721\ : InMux
    port map (
            O => \N__15250\,
            I => \N__15237\
        );

    \I__2720\ : InMux
    port map (
            O => \N__15249\,
            I => \N__15237\
        );

    \I__2719\ : InMux
    port map (
            O => \N__15248\,
            I => \N__15237\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__15237\,
            I => \N__15234\
        );

    \I__2717\ : Odrv4
    port map (
            O => \N__15234\,
            I => \Lab_UT.dictrl.N_1459_1\
        );

    \I__2716\ : InMux
    port map (
            O => \N__15231\,
            I => \N__15228\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__15228\,
            I => \Lab_UT.dictrl.N_40_8\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__15225\,
            I => \Lab_UT.dictrl.N_40_3_cascade_\
        );

    \I__2713\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15219\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__15219\,
            I => \Lab_UT.dictrl.N_1102_2\
        );

    \I__2711\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15213\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__15213\,
            I => \N__15210\
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__15210\,
            I => \Lab_UT.dictrl.g2_1_2\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__15207\,
            I => \Lab_UT.dictrl.N_1462_2_cascade_\
        );

    \I__2707\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15201\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__15201\,
            I => \N__15197\
        );

    \I__2705\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15194\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__15197\,
            I => \N__15189\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__15194\,
            I => \N__15189\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__15189\,
            I => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4\
        );

    \I__2701\ : CascadeMux
    port map (
            O => \N__15186\,
            I => \Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_\
        );

    \I__2700\ : InMux
    port map (
            O => \N__15183\,
            I => \N__15177\
        );

    \I__2699\ : InMux
    port map (
            O => \N__15182\,
            I => \N__15177\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__15177\,
            I => \N__15174\
        );

    \I__2697\ : Odrv4
    port map (
            O => \N__15174\,
            I => \Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__15171\,
            I => \Lab_UT.dictrl.N_11_0_cascade_\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__15168\,
            I => \N__15165\
        );

    \I__2694\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15162\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__15162\,
            I => \N__15159\
        );

    \I__2692\ : Odrv12
    port map (
            O => \N__15159\,
            I => \Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1\
        );

    \I__2691\ : InMux
    port map (
            O => \N__15156\,
            I => \N__15138\
        );

    \I__2690\ : InMux
    port map (
            O => \N__15155\,
            I => \N__15138\
        );

    \I__2689\ : InMux
    port map (
            O => \N__15154\,
            I => \N__15138\
        );

    \I__2688\ : InMux
    port map (
            O => \N__15153\,
            I => \N__15138\
        );

    \I__2687\ : InMux
    port map (
            O => \N__15152\,
            I => \N__15138\
        );

    \I__2686\ : InMux
    port map (
            O => \N__15151\,
            I => \N__15138\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__15138\,
            I => \Lab_UT.dictrl.m27_1\
        );

    \I__2684\ : InMux
    port map (
            O => \N__15135\,
            I => \N__15125\
        );

    \I__2683\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15125\
        );

    \I__2682\ : InMux
    port map (
            O => \N__15133\,
            I => \N__15116\
        );

    \I__2681\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15116\
        );

    \I__2680\ : InMux
    port map (
            O => \N__15131\,
            I => \N__15116\
        );

    \I__2679\ : InMux
    port map (
            O => \N__15130\,
            I => \N__15116\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__15125\,
            I => \N__15111\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__15116\,
            I => \N__15111\
        );

    \I__2676\ : Odrv4
    port map (
            O => \N__15111\,
            I => \Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83\
        );

    \I__2675\ : InMux
    port map (
            O => \N__15108\,
            I => \N__15105\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__15105\,
            I => \N__15102\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__15102\,
            I => \Lab_UT.dictrl.N_61\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__15099\,
            I => \Lab_UT.dictrl.N_62_cascade_\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__15096\,
            I => \N__15093\
        );

    \I__2670\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15090\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__15090\,
            I => \N__15087\
        );

    \I__2668\ : Span4Mux_h
    port map (
            O => \N__15087\,
            I => \N__15083\
        );

    \I__2667\ : InMux
    port map (
            O => \N__15086\,
            I => \N__15080\
        );

    \I__2666\ : Span4Mux_v
    port map (
            O => \N__15083\,
            I => \N__15077\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__15080\,
            I => \N__15074\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__15077\,
            I => \Lab_UT.dictrl.N_9_0\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__15074\,
            I => \Lab_UT.dictrl.N_9_0\
        );

    \I__2662\ : InMux
    port map (
            O => \N__15069\,
            I => \N__15063\
        );

    \I__2661\ : InMux
    port map (
            O => \N__15068\,
            I => \N__15063\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__15063\,
            I => \Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1\
        );

    \I__2659\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15057\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__15057\,
            I => \N__15054\
        );

    \I__2657\ : Span4Mux_s2_v
    port map (
            O => \N__15054\,
            I => \N__15051\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__15051\,
            I => \Lab_UT.dictrl.state_fast_1\
        );

    \I__2655\ : InMux
    port map (
            O => \N__15048\,
            I => \N__15033\
        );

    \I__2654\ : InMux
    port map (
            O => \N__15047\,
            I => \N__15033\
        );

    \I__2653\ : InMux
    port map (
            O => \N__15046\,
            I => \N__15033\
        );

    \I__2652\ : InMux
    port map (
            O => \N__15045\,
            I => \N__15033\
        );

    \I__2651\ : InMux
    port map (
            O => \N__15044\,
            I => \N__15033\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__15033\,
            I => \N__15030\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__15030\,
            I => \N__15027\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__15027\,
            I => \N__15024\
        );

    \I__2647\ : Odrv4
    port map (
            O => \N__15024\,
            I => \Lab_UT.dictrl.N_62_1\
        );

    \I__2646\ : CascadeMux
    port map (
            O => \N__15021\,
            I => \N__15018\
        );

    \I__2645\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15015\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__15015\,
            I => \N__15012\
        );

    \I__2643\ : Span12Mux_v
    port map (
            O => \N__15012\,
            I => \N__15009\
        );

    \I__2642\ : Odrv12
    port map (
            O => \N__15009\,
            I => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\
        );

    \I__2641\ : InMux
    port map (
            O => \N__15006\,
            I => \N__15003\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__15003\,
            I => \N__14999\
        );

    \I__2639\ : InMux
    port map (
            O => \N__15002\,
            I => \N__14996\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__14999\,
            I => \N__14993\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__14996\,
            I => \N__14990\
        );

    \I__2636\ : Odrv4
    port map (
            O => \N__14993\,
            I => \Lab_UT.dictrl.N_79\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__14990\,
            I => \Lab_UT.dictrl.N_79\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14985\,
            I => \N__14982\
        );

    \I__2633\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14979\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__14979\,
            I => \Lab_UT.dictrl.state_i_4_1\
        );

    \I__2631\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14973\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__14973\,
            I => \N__14970\
        );

    \I__2629\ : Span12Mux_s11_v
    port map (
            O => \N__14970\,
            I => \N__14967\
        );

    \I__2628\ : Odrv12
    port map (
            O => \N__14967\,
            I => \Lab_UT.dictrl.N_99\
        );

    \I__2627\ : InMux
    port map (
            O => \N__14964\,
            I => \N__14961\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__14961\,
            I => \N__14954\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14947\
        );

    \I__2624\ : InMux
    port map (
            O => \N__14959\,
            I => \N__14944\
        );

    \I__2623\ : InMux
    port map (
            O => \N__14958\,
            I => \N__14941\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14957\,
            I => \N__14938\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__14954\,
            I => \N__14935\
        );

    \I__2620\ : InMux
    port map (
            O => \N__14953\,
            I => \N__14932\
        );

    \I__2619\ : InMux
    port map (
            O => \N__14952\,
            I => \N__14929\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14926\
        );

    \I__2617\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14923\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14947\,
            I => \N__14914\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__14944\,
            I => \N__14914\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__14941\,
            I => \N__14914\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__14938\,
            I => \N__14914\
        );

    \I__2612\ : Sp12to4
    port map (
            O => \N__14935\,
            I => \N__14907\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__14932\,
            I => \N__14907\
        );

    \I__2610\ : LocalMux
    port map (
            O => \N__14929\,
            I => \N__14907\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14926\,
            I => \buart__rx_bitcount_3\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__14923\,
            I => \buart__rx_bitcount_3\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__14914\,
            I => \buart__rx_bitcount_3\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__14907\,
            I => \buart__rx_bitcount_3\
        );

    \I__2605\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14895\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14895\,
            I => \N__14890\
        );

    \I__2603\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14887\
        );

    \I__2602\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14884\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__14890\,
            I => \N__14879\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__14887\,
            I => \N__14874\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14884\,
            I => \N__14874\
        );

    \I__2598\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14869\
        );

    \I__2597\ : InMux
    port map (
            O => \N__14882\,
            I => \N__14869\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__14879\,
            I => \N__14866\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__14874\,
            I => \N__14863\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__14869\,
            I => \buart__rx_valid_3\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__14866\,
            I => \buart__rx_valid_3\
        );

    \I__2592\ : Odrv4
    port map (
            O => \N__14863\,
            I => \buart__rx_valid_3\
        );

    \I__2591\ : CascadeMux
    port map (
            O => \N__14856\,
            I => \Lab_UT.dictrl.g0_0_2_1_cascade_\
        );

    \I__2590\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__14850\,
            I => \Lab_UT.dictrl.g2_1_0\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__14847\,
            I => \Lab_UT.dictrl.g0_0_2_cascade_\
        );

    \I__2587\ : CascadeMux
    port map (
            O => \N__14844\,
            I => \N__14841\
        );

    \I__2586\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14838\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__14838\,
            I => \Lab_UT.dictrl.g0_12_a6_0_1\
        );

    \I__2584\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14829\
        );

    \I__2583\ : CascadeMux
    port map (
            O => \N__14834\,
            I => \N__14821\
        );

    \I__2582\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14818\
        );

    \I__2581\ : InMux
    port map (
            O => \N__14832\,
            I => \N__14815\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__14829\,
            I => \N__14812\
        );

    \I__2579\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14803\
        );

    \I__2578\ : InMux
    port map (
            O => \N__14827\,
            I => \N__14803\
        );

    \I__2577\ : InMux
    port map (
            O => \N__14826\,
            I => \N__14803\
        );

    \I__2576\ : InMux
    port map (
            O => \N__14825\,
            I => \N__14803\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14798\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14821\,
            I => \N__14798\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__14818\,
            I => \N__14793\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__14815\,
            I => \N__14793\
        );

    \I__2571\ : Span4Mux_s3_v
    port map (
            O => \N__14812\,
            I => \N__14786\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14803\,
            I => \N__14786\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__14798\,
            I => \N__14786\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__14793\,
            I => \N__14783\
        );

    \I__2567\ : Span4Mux_v
    port map (
            O => \N__14786\,
            I => \N__14780\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__14783\,
            I => \Lab_UT.dictrl.state_2_rep1\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__14780\,
            I => \Lab_UT.dictrl.state_2_rep1\
        );

    \I__2564\ : CEMux
    port map (
            O => \N__14775\,
            I => \N__14772\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__14772\,
            I => \N__14769\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__14769\,
            I => \N__14766\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__14766\,
            I => \N__14763\
        );

    \I__2560\ : Odrv4
    port map (
            O => \N__14763\,
            I => \Lab_UT.didp.regrce4.LdAMtens_0\
        );

    \I__2559\ : CascadeMux
    port map (
            O => \N__14760\,
            I => \Lab_UT.didp.countrce4.q_5_3_cascade_\
        );

    \I__2558\ : InMux
    port map (
            O => \N__14757\,
            I => \N__14752\
        );

    \I__2557\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14747\
        );

    \I__2556\ : InMux
    port map (
            O => \N__14755\,
            I => \N__14747\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__14752\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__14747\,
            I => \Lab_UT.di_AMtens_3\
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__14742\,
            I => \N__14739\
        );

    \I__2552\ : InMux
    port map (
            O => \N__14739\,
            I => \N__14736\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__14736\,
            I => \Lab_UT.didp.countrce4.un20_qPone\
        );

    \I__2550\ : InMux
    port map (
            O => \N__14733\,
            I => \N__14730\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__14730\,
            I => \uu2.bitmap_pmux_15_ns_1\
        );

    \I__2548\ : InMux
    port map (
            O => \N__14727\,
            I => \N__14723\
        );

    \I__2547\ : InMux
    port map (
            O => \N__14726\,
            I => \N__14719\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__14723\,
            I => \N__14715\
        );

    \I__2545\ : InMux
    port map (
            O => \N__14722\,
            I => \N__14712\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__14719\,
            I => \N__14709\
        );

    \I__2543\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14706\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__14715\,
            I => \o_One_Sec_Pulse\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__14712\,
            I => \o_One_Sec_Pulse\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__14709\,
            I => \o_One_Sec_Pulse\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__14706\,
            I => \o_One_Sec_Pulse\
        );

    \I__2538\ : InMux
    port map (
            O => \N__14697\,
            I => \N__14691\
        );

    \I__2537\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14691\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__14691\,
            I => \N__14688\
        );

    \I__2535\ : Odrv4
    port map (
            O => \N__14688\,
            I => \uu2.bitmapZ0Z_111\
        );

    \I__2534\ : InMux
    port map (
            O => \N__14685\,
            I => \N__14680\
        );

    \I__2533\ : InMux
    port map (
            O => \N__14684\,
            I => \N__14677\
        );

    \I__2532\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14674\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__14680\,
            I => \N__14671\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__14677\,
            I => \N__14668\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__14674\,
            I => \N__14662\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__14671\,
            I => \N__14662\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__14668\,
            I => \N__14659\
        );

    \I__2526\ : InMux
    port map (
            O => \N__14667\,
            I => \N__14656\
        );

    \I__2525\ : Span4Mux_v
    port map (
            O => \N__14662\,
            I => \N__14653\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__14659\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__14656\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__14653\,
            I => \uu2.vram_rd_clkZ0\
        );

    \I__2521\ : InMux
    port map (
            O => \N__14646\,
            I => \N__14643\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__14643\,
            I => \uu2.bitmapZ0Z_194\
        );

    \I__2519\ : CascadeMux
    port map (
            O => \N__14640\,
            I => \N__14637\
        );

    \I__2518\ : InMux
    port map (
            O => \N__14637\,
            I => \N__14634\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__14634\,
            I => \N__14631\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__14631\,
            I => \uu2.bitmapZ0Z_34\
        );

    \I__2515\ : InMux
    port map (
            O => \N__14628\,
            I => \N__14625\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__14625\,
            I => \uu2.bitmapZ0Z_290\
        );

    \I__2513\ : InMux
    port map (
            O => \N__14622\,
            I => \N__14619\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__14619\,
            I => \uu2.bitmapZ0Z_40\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__14616\,
            I => \N__14613\
        );

    \I__2510\ : InMux
    port map (
            O => \N__14613\,
            I => \N__14610\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__14610\,
            I => \uu2.bitmapZ0Z_296\
        );

    \I__2508\ : InMux
    port map (
            O => \N__14607\,
            I => \N__14604\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__14604\,
            I => \uu2.N_207\
        );

    \I__2506\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14598\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__14598\,
            I => \uu2.bitmapZ0Z_168\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__14595\,
            I => \N__14592\
        );

    \I__2503\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14589\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__14589\,
            I => \N__14586\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__14586\,
            I => \uu2.N_195\
        );

    \I__2500\ : InMux
    port map (
            O => \N__14583\,
            I => \N__14580\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__14580\,
            I => \uu2.bitmapZ0Z_66\
        );

    \I__2498\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14574\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__14574\,
            I => \N__14571\
        );

    \I__2496\ : Odrv4
    port map (
            O => \N__14571\,
            I => \uu2.bitmapZ0Z_162\
        );

    \I__2495\ : CascadeMux
    port map (
            O => \N__14568\,
            I => \N__14564\
        );

    \I__2494\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14556\
        );

    \I__2493\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14556\
        );

    \I__2492\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14556\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__14556\,
            I => \uu2.N_91\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__14553\,
            I => \uu2.N_28_cascade_\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__14550\,
            I => \uu2.bitmap_pmux_26_i_m2_1_cascade_\
        );

    \I__2488\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14544\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__14544\,
            I => \N__14541\
        );

    \I__2486\ : Odrv4
    port map (
            O => \N__14541\,
            I => \uu2.bitmap_pmux_sn_N_20\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__14538\,
            I => \uu2.N_55_cascade_\
        );

    \I__2484\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14532\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__14532\,
            I => \uu2.bitmap_pmux_sn_i7_mux_0\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__14529\,
            I => \uu2.N_406_cascade_\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__14526\,
            I => \N__14523\
        );

    \I__2480\ : InMux
    port map (
            O => \N__14523\,
            I => \N__14517\
        );

    \I__2479\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14517\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__14517\,
            I => \uu2.bitmap_pmux\
        );

    \I__2477\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14511\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__14511\,
            I => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\
        );

    \I__2475\ : InMux
    port map (
            O => \N__14508\,
            I => \N__14505\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14502\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__14502\,
            I => \Lab_UT.dictrl.next_state_RNO_3Z0Z_0\
        );

    \I__2472\ : CascadeMux
    port map (
            O => \N__14499\,
            I => \Lab_UT.dictrl.m67_am_1_0_cascade_\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__14496\,
            I => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\
        );

    \I__2470\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14490\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__14490\,
            I => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\
        );

    \I__2468\ : InMux
    port map (
            O => \N__14487\,
            I => \N__14484\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__14484\,
            I => \Lab_UT.dictrl.G_17_i_a5_0\
        );

    \I__2466\ : InMux
    port map (
            O => \N__14481\,
            I => \N__14477\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__14480\,
            I => \N__14474\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__14477\,
            I => \N__14471\
        );

    \I__2463\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14468\
        );

    \I__2462\ : Span4Mux_h
    port map (
            O => \N__14471\,
            I => \N__14465\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__14468\,
            I => \Lab_UT.dictrl.N_65\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__14465\,
            I => \Lab_UT.dictrl.N_65\
        );

    \I__2459\ : CascadeMux
    port map (
            O => \N__14460\,
            I => \Lab_UT.dictrl.N_65_cascade_\
        );

    \I__2458\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14454\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__14454\,
            I => \Lab_UT.dictrl.N_101\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__14451\,
            I => \N__14448\
        );

    \I__2455\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14445\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__14445\,
            I => \N__14442\
        );

    \I__2453\ : Odrv12
    port map (
            O => \N__14442\,
            I => \uu2.mem0.w_addr_5\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__14439\,
            I => \N__14436\
        );

    \I__2451\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14433\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__14433\,
            I => \N__14430\
        );

    \I__2449\ : Span4Mux_h
    port map (
            O => \N__14430\,
            I => \N__14427\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__14427\,
            I => \uu2.mem0.w_addr_6\
        );

    \I__2447\ : InMux
    port map (
            O => \N__14424\,
            I => \N__14421\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__14421\,
            I => \N__14417\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__14420\,
            I => \N__14412\
        );

    \I__2444\ : Span4Mux_s1_v
    port map (
            O => \N__14417\,
            I => \N__14409\
        );

    \I__2443\ : InMux
    port map (
            O => \N__14416\,
            I => \N__14402\
        );

    \I__2442\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14402\
        );

    \I__2441\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14402\
        );

    \I__2440\ : Odrv4
    port map (
            O => \N__14409\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14402\,
            I => \uu2.w_addr_userZ0Z_7\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__14397\,
            I => \N__14394\
        );

    \I__2437\ : InMux
    port map (
            O => \N__14394\,
            I => \N__14391\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__14391\,
            I => \N__14388\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__14388\,
            I => \N__14385\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__14385\,
            I => \uu2.mem0.w_addr_7\
        );

    \I__2433\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14379\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__14379\,
            I => \Lab_UT.dictrl.g2_0_3_3\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__14376\,
            I => \Lab_UT.dictrl.g2_0_4_3_cascade_\
        );

    \I__2430\ : InMux
    port map (
            O => \N__14373\,
            I => \N__14363\
        );

    \I__2429\ : InMux
    port map (
            O => \N__14372\,
            I => \N__14363\
        );

    \I__2428\ : InMux
    port map (
            O => \N__14371\,
            I => \N__14360\
        );

    \I__2427\ : InMux
    port map (
            O => \N__14370\,
            I => \N__14357\
        );

    \I__2426\ : InMux
    port map (
            O => \N__14369\,
            I => \N__14352\
        );

    \I__2425\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14352\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__14363\,
            I => \N__14347\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__14360\,
            I => \N__14342\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14342\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__14352\,
            I => \N__14339\
        );

    \I__2420\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14334\
        );

    \I__2419\ : InMux
    port map (
            O => \N__14350\,
            I => \N__14334\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__14347\,
            I => \N__14326\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__14342\,
            I => \N__14323\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14318\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__14334\,
            I => \N__14318\
        );

    \I__2414\ : InMux
    port map (
            O => \N__14333\,
            I => \N__14315\
        );

    \I__2413\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14306\
        );

    \I__2412\ : InMux
    port map (
            O => \N__14331\,
            I => \N__14306\
        );

    \I__2411\ : InMux
    port map (
            O => \N__14330\,
            I => \N__14306\
        );

    \I__2410\ : InMux
    port map (
            O => \N__14329\,
            I => \N__14306\
        );

    \I__2409\ : Odrv4
    port map (
            O => \N__14326\,
            I => \Lab_UT.dictrl.m12Z0Z_1\
        );

    \I__2408\ : Odrv4
    port map (
            O => \N__14323\,
            I => \Lab_UT.dictrl.m12Z0Z_1\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__14318\,
            I => \Lab_UT.dictrl.m12Z0Z_1\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__14315\,
            I => \Lab_UT.dictrl.m12Z0Z_1\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__14306\,
            I => \Lab_UT.dictrl.m12Z0Z_1\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__14295\,
            I => \Lab_UT.dictrl.N_11_1_cascade_\
        );

    \I__2403\ : InMux
    port map (
            O => \N__14292\,
            I => \N__14289\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__14289\,
            I => \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__14286\,
            I => \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_\
        );

    \I__2400\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14273\
        );

    \I__2399\ : InMux
    port map (
            O => \N__14282\,
            I => \N__14270\
        );

    \I__2398\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14261\
        );

    \I__2397\ : InMux
    port map (
            O => \N__14280\,
            I => \N__14261\
        );

    \I__2396\ : InMux
    port map (
            O => \N__14279\,
            I => \N__14261\
        );

    \I__2395\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14261\
        );

    \I__2394\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14258\
        );

    \I__2393\ : InMux
    port map (
            O => \N__14276\,
            I => \N__14255\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__14273\,
            I => bu_rx_data_fast_6
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__14270\,
            I => bu_rx_data_fast_6
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__14261\,
            I => bu_rx_data_fast_6
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__14258\,
            I => bu_rx_data_fast_6
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__14255\,
            I => bu_rx_data_fast_6
        );

    \I__2387\ : CEMux
    port map (
            O => \N__14244\,
            I => \N__14220\
        );

    \I__2386\ : CEMux
    port map (
            O => \N__14243\,
            I => \N__14220\
        );

    \I__2385\ : CEMux
    port map (
            O => \N__14242\,
            I => \N__14220\
        );

    \I__2384\ : CEMux
    port map (
            O => \N__14241\,
            I => \N__14220\
        );

    \I__2383\ : CEMux
    port map (
            O => \N__14240\,
            I => \N__14220\
        );

    \I__2382\ : CEMux
    port map (
            O => \N__14239\,
            I => \N__14220\
        );

    \I__2381\ : CEMux
    port map (
            O => \N__14238\,
            I => \N__14220\
        );

    \I__2380\ : CEMux
    port map (
            O => \N__14237\,
            I => \N__14220\
        );

    \I__2379\ : GlobalMux
    port map (
            O => \N__14220\,
            I => \N__14217\
        );

    \I__2378\ : gio2CtrlBuf
    port map (
            O => \N__14217\,
            I => \buart.Z_rx.sample_g\
        );

    \I__2377\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14211\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__14211\,
            I => \N__14208\
        );

    \I__2375\ : Odrv12
    port map (
            O => \N__14208\,
            I => \Lab_UT.dictrl.N_100\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__14205\,
            I => \N__14202\
        );

    \I__2373\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14199\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__14199\,
            I => \N__14196\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__14196\,
            I => \Lab_UT.dictrl.next_state_RNO_8Z0Z_0\
        );

    \I__2370\ : InMux
    port map (
            O => \N__14193\,
            I => \N__14190\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__14190\,
            I => \N__14187\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__14187\,
            I => \Lab_UT.dictrl.m63_d_0_ns_1\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__14184\,
            I => \Lab_UT.dictrl.m59_3_cascade_\
        );

    \I__2366\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14178\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__14178\,
            I => \Lab_UT.dictrl.g2_0_3_4\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__14175\,
            I => \Lab_UT.dictrl.g2_0_4_4_cascade_\
        );

    \I__2363\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14169\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__14169\,
            I => \Lab_UT.dictrl.g2_0_3_2\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__14166\,
            I => \Lab_UT.dictrl.g2_0_4_2_cascade_\
        );

    \I__2360\ : InMux
    port map (
            O => \N__14163\,
            I => \N__14160\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__14160\,
            I => \Lab_UT.dictrl.g2_0_3\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__14157\,
            I => \Lab_UT.dictrl.g2_0_4_cascade_\
        );

    \I__2357\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14140\
        );

    \I__2356\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14140\
        );

    \I__2355\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14140\
        );

    \I__2354\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14140\
        );

    \I__2353\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14137\
        );

    \I__2352\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14134\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14129\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__14137\,
            I => \N__14129\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__14134\,
            I => bu_rx_data_fast_0
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__14129\,
            I => bu_rx_data_fast_0
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__14124\,
            I => \N__14118\
        );

    \I__2346\ : CascadeMux
    port map (
            O => \N__14123\,
            I => \N__14115\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__14122\,
            I => \N__14112\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__14121\,
            I => \N__14109\
        );

    \I__2343\ : InMux
    port map (
            O => \N__14118\,
            I => \N__14098\
        );

    \I__2342\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14098\
        );

    \I__2341\ : InMux
    port map (
            O => \N__14112\,
            I => \N__14098\
        );

    \I__2340\ : InMux
    port map (
            O => \N__14109\,
            I => \N__14098\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__14108\,
            I => \N__14095\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__14107\,
            I => \N__14091\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14088\
        );

    \I__2336\ : InMux
    port map (
            O => \N__14095\,
            I => \N__14085\
        );

    \I__2335\ : InMux
    port map (
            O => \N__14094\,
            I => \N__14082\
        );

    \I__2334\ : InMux
    port map (
            O => \N__14091\,
            I => \N__14079\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__14088\,
            I => \N__14076\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__14085\,
            I => \N__14073\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__14082\,
            I => \N__14070\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__14079\,
            I => bu_rx_data_fast_4
        );

    \I__2329\ : Odrv4
    port map (
            O => \N__14076\,
            I => bu_rx_data_fast_4
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__14073\,
            I => bu_rx_data_fast_4
        );

    \I__2327\ : Odrv4
    port map (
            O => \N__14070\,
            I => bu_rx_data_fast_4
        );

    \I__2326\ : InMux
    port map (
            O => \N__14061\,
            I => \N__14047\
        );

    \I__2325\ : InMux
    port map (
            O => \N__14060\,
            I => \N__14047\
        );

    \I__2324\ : InMux
    port map (
            O => \N__14059\,
            I => \N__14047\
        );

    \I__2323\ : InMux
    port map (
            O => \N__14058\,
            I => \N__14047\
        );

    \I__2322\ : InMux
    port map (
            O => \N__14057\,
            I => \N__14042\
        );

    \I__2321\ : InMux
    port map (
            O => \N__14056\,
            I => \N__14039\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__14047\,
            I => \N__14036\
        );

    \I__2319\ : InMux
    port map (
            O => \N__14046\,
            I => \N__14031\
        );

    \I__2318\ : InMux
    port map (
            O => \N__14045\,
            I => \N__14031\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__14042\,
            I => \N__14026\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__14039\,
            I => \N__14026\
        );

    \I__2315\ : Span4Mux_v
    port map (
            O => \N__14036\,
            I => \N__14023\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__14031\,
            I => \N__14018\
        );

    \I__2313\ : Span4Mux_v
    port map (
            O => \N__14026\,
            I => \N__14018\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__14023\,
            I => bu_rx_data_3_rep1
        );

    \I__2311\ : Odrv4
    port map (
            O => \N__14018\,
            I => bu_rx_data_3_rep1
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__14013\,
            I => \N__14010\
        );

    \I__2309\ : InMux
    port map (
            O => \N__14010\,
            I => \N__14007\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__14007\,
            I => \N__14003\
        );

    \I__2307\ : InMux
    port map (
            O => \N__14006\,
            I => \N__14000\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__14003\,
            I => \Lab_UT.dictrl.m15Z0Z_1\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__14000\,
            I => \Lab_UT.dictrl.m15Z0Z_1\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13995\,
            I => \N__13992\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13992\,
            I => \N__13987\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13991\,
            I => \N__13984\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13990\,
            I => \N__13981\
        );

    \I__2300\ : Odrv4
    port map (
            O => \N__13987\,
            I => \Lab_UT.dictrl.N_88_mux\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13984\,
            I => \Lab_UT.dictrl.N_88_mux\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13981\,
            I => \Lab_UT.dictrl.N_88_mux\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \Lab_UT.dictrl.g2_0_4_1_cascade_\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__13971\,
            I => \Lab_UT.dictrl.m53_d_1_2_cascade_\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__13968\,
            I => \Lab_UT.dictrl.N_45_cascade_\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13960\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13951\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13963\,
            I => \N__13948\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13960\,
            I => \N__13945\
        );

    \I__2290\ : InMux
    port map (
            O => \N__13959\,
            I => \N__13936\
        );

    \I__2289\ : InMux
    port map (
            O => \N__13958\,
            I => \N__13936\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13936\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13956\,
            I => \N__13936\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13931\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13954\,
            I => \N__13931\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__13951\,
            I => \N__13928\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__13948\,
            I => \N__13919\
        );

    \I__2282\ : Span4Mux_v
    port map (
            O => \N__13945\,
            I => \N__13919\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13936\,
            I => \N__13919\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__13931\,
            I => \N__13916\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__13928\,
            I => \N__13913\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13908\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13908\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__13919\,
            I => \N__13905\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__13916\,
            I => \N__13902\
        );

    \I__2274\ : Odrv4
    port map (
            O => \N__13913\,
            I => bu_rx_data_1_rep2
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13908\,
            I => bu_rx_data_1_rep2
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__13905\,
            I => bu_rx_data_1_rep2
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__13902\,
            I => bu_rx_data_1_rep2
        );

    \I__2270\ : InMux
    port map (
            O => \N__13893\,
            I => \N__13890\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__13890\,
            I => \Lab_UT.dictrl.g2_0_3_1\
        );

    \I__2268\ : CascadeMux
    port map (
            O => \N__13887\,
            I => \N__13878\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__13886\,
            I => \N__13872\
        );

    \I__2266\ : CascadeMux
    port map (
            O => \N__13885\,
            I => \N__13869\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__13884\,
            I => \N__13866\
        );

    \I__2264\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13863\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13882\,
            I => \N__13860\
        );

    \I__2262\ : InMux
    port map (
            O => \N__13881\,
            I => \N__13853\
        );

    \I__2261\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13853\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13877\,
            I => \N__13853\
        );

    \I__2259\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13850\
        );

    \I__2258\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13847\
        );

    \I__2257\ : InMux
    port map (
            O => \N__13872\,
            I => \N__13840\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13869\,
            I => \N__13840\
        );

    \I__2255\ : InMux
    port map (
            O => \N__13866\,
            I => \N__13840\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__13863\,
            I => \N__13835\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__13860\,
            I => \N__13830\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__13853\,
            I => \N__13830\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__13850\,
            I => \N__13827\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13824\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__13840\,
            I => \N__13821\
        );

    \I__2248\ : InMux
    port map (
            O => \N__13839\,
            I => \N__13816\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13838\,
            I => \N__13816\
        );

    \I__2246\ : Span4Mux_h
    port map (
            O => \N__13835\,
            I => \N__13811\
        );

    \I__2245\ : Span4Mux_h
    port map (
            O => \N__13830\,
            I => \N__13811\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__13827\,
            I => \N__13804\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__13824\,
            I => \N__13804\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__13821\,
            I => \N__13804\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__13816\,
            I => bu_rx_data_2_rep2
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__13811\,
            I => bu_rx_data_2_rep2
        );

    \I__2239\ : Odrv4
    port map (
            O => \N__13804\,
            I => bu_rx_data_2_rep2
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__13797\,
            I => \N__13794\
        );

    \I__2237\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13791\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13791\,
            I => \N__13787\
        );

    \I__2235\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \N__13784\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__13787\,
            I => \N__13781\
        );

    \I__2233\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13778\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__13781\,
            I => \Lab_UT_dictrl_m59_1\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__13778\,
            I => \Lab_UT_dictrl_m59_1\
        );

    \I__2230\ : InMux
    port map (
            O => \N__13773\,
            I => \N__13770\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__13770\,
            I => \N__13767\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__13767\,
            I => \Lab_UT.dictrl.g0_12_a6_3_6\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13761\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13758\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__13758\,
            I => \Lab_UT.dictrl.N_10\
        );

    \I__2224\ : InMux
    port map (
            O => \N__13755\,
            I => \N__13752\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__13752\,
            I => \Lab_UT.dictrl.g0_12_1\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__13749\,
            I => \Lab_UT.dictrl.m15Z0Z_1_cascade_\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13746\,
            I => \N__13743\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__13743\,
            I => \N__13740\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__13740\,
            I => \Lab_UT.dictrl.N_8_0\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__13737\,
            I => \Lab_UT.dictrl.N_93_cascade_\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__13734\,
            I => \N__13731\
        );

    \I__2216\ : InMux
    port map (
            O => \N__13731\,
            I => \N__13728\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__13728\,
            I => \Lab_UT.dictrl.N_10_0\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13722\
        );

    \I__2213\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13719\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__13719\,
            I => \N__13716\
        );

    \I__2211\ : Span4Mux_h
    port map (
            O => \N__13716\,
            I => \N__13713\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__13713\,
            I => \Lab_UT.dictrl.g0_i_a4_0_1\
        );

    \I__2209\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13707\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__13707\,
            I => \Lab_UT.dictrl.g0_i_a4_0_3\
        );

    \I__2207\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13692\
        );

    \I__2206\ : InMux
    port map (
            O => \N__13703\,
            I => \N__13692\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13692\
        );

    \I__2204\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13689\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \N__13684\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__13699\,
            I => \N__13681\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__13692\,
            I => \N__13673\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__13689\,
            I => \N__13673\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__13688\,
            I => \N__13668\
        );

    \I__2198\ : InMux
    port map (
            O => \N__13687\,
            I => \N__13663\
        );

    \I__2197\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13663\
        );

    \I__2196\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13658\
        );

    \I__2195\ : InMux
    port map (
            O => \N__13680\,
            I => \N__13658\
        );

    \I__2194\ : InMux
    port map (
            O => \N__13679\,
            I => \N__13653\
        );

    \I__2193\ : InMux
    port map (
            O => \N__13678\,
            I => \N__13653\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__13673\,
            I => \N__13650\
        );

    \I__2191\ : InMux
    port map (
            O => \N__13672\,
            I => \N__13647\
        );

    \I__2190\ : InMux
    port map (
            O => \N__13671\,
            I => \N__13642\
        );

    \I__2189\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13642\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__13663\,
            I => \N__13639\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__13658\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__13653\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2185\ : Odrv4
    port map (
            O => \N__13650\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__13647\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__13642\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__13639\,
            I => \Lab_UT.dispString.cntZ0Z_2\
        );

    \I__2181\ : InMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__13623\,
            I => \Lab_UT.dispString.b1_m_1\
        );

    \I__2179\ : CascadeMux
    port map (
            O => \N__13620\,
            I => \Lab_UT.dispString.m67_ns_1_cascade_\
        );

    \I__2178\ : InMux
    port map (
            O => \N__13617\,
            I => \N__13614\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__2176\ : Odrv4
    port map (
            O => \N__13611\,
            I => \Lab_UT.dispString.N_143\
        );

    \I__2175\ : InMux
    port map (
            O => \N__13608\,
            I => \N__13605\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__13605\,
            I => \N__13601\
        );

    \I__2173\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13598\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__13601\,
            I => \Lab_UT.dispString.N_23_0\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__13598\,
            I => \Lab_UT.dispString.N_23_0\
        );

    \I__2170\ : InMux
    port map (
            O => \N__13593\,
            I => \N__13590\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__13590\,
            I => \Lab_UT.dispString.N_158\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__13587\,
            I => \Lab_UT.dispString.m90_ns_1_cascade_\
        );

    \I__2167\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13581\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__13581\,
            I => \N__13578\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__13578\,
            I => \Lab_UT.dispString.N_164\
        );

    \I__2164\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13563\
        );

    \I__2163\ : InMux
    port map (
            O => \N__13574\,
            I => \N__13563\
        );

    \I__2162\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13556\
        );

    \I__2161\ : InMux
    port map (
            O => \N__13572\,
            I => \N__13556\
        );

    \I__2160\ : InMux
    port map (
            O => \N__13571\,
            I => \N__13556\
        );

    \I__2159\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13550\
        );

    \I__2158\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13550\
        );

    \I__2157\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13547\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__13563\,
            I => \N__13530\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__13556\,
            I => \N__13530\
        );

    \I__2154\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13527\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__13550\,
            I => \N__13524\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13521\
        );

    \I__2151\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13514\
        );

    \I__2150\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13514\
        );

    \I__2149\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13514\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13511\
        );

    \I__2147\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13508\
        );

    \I__2146\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13505\
        );

    \I__2145\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13502\
        );

    \I__2144\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13493\
        );

    \I__2143\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13493\
        );

    \I__2142\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13493\
        );

    \I__2141\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13493\
        );

    \I__2140\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13490\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__13530\,
            I => \N__13487\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__13527\,
            I => \N__13484\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__13524\,
            I => \N__13477\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__13521\,
            I => \N__13477\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__13514\,
            I => \N__13477\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__13511\,
            I => \N__13474\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__13508\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__13505\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__13502\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__13493\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__13490\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__13487\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__13484\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2126\ : Odrv4
    port map (
            O => \N__13477\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__13474\,
            I => \Lab_UT.dispString.cntZ0Z_0\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__13455\,
            I => \N__13448\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__13454\,
            I => \N__13444\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__13453\,
            I => \N__13441\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__13452\,
            I => \N__13438\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__13451\,
            I => \N__13435\
        );

    \I__2119\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13426\
        );

    \I__2118\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13426\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13444\,
            I => \N__13426\
        );

    \I__2116\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13423\
        );

    \I__2115\ : InMux
    port map (
            O => \N__13438\,
            I => \N__13416\
        );

    \I__2114\ : InMux
    port map (
            O => \N__13435\,
            I => \N__13416\
        );

    \I__2113\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13416\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__13433\,
            I => \N__13405\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__13426\,
            I => \N__13400\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__13423\,
            I => \N__13395\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__13416\,
            I => \N__13395\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13390\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13390\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13413\,
            I => \N__13387\
        );

    \I__2105\ : InMux
    port map (
            O => \N__13412\,
            I => \N__13382\
        );

    \I__2104\ : InMux
    port map (
            O => \N__13411\,
            I => \N__13382\
        );

    \I__2103\ : InMux
    port map (
            O => \N__13410\,
            I => \N__13375\
        );

    \I__2102\ : InMux
    port map (
            O => \N__13409\,
            I => \N__13375\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13375\
        );

    \I__2100\ : InMux
    port map (
            O => \N__13405\,
            I => \N__13370\
        );

    \I__2099\ : InMux
    port map (
            O => \N__13404\,
            I => \N__13370\
        );

    \I__2098\ : InMux
    port map (
            O => \N__13403\,
            I => \N__13367\
        );

    \I__2097\ : Span4Mux_v
    port map (
            O => \N__13400\,
            I => \N__13360\
        );

    \I__2096\ : Span4Mux_v
    port map (
            O => \N__13395\,
            I => \N__13360\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__13390\,
            I => \N__13360\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__13387\,
            I => \N__13357\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__13382\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__13375\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__13370\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__13367\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__13360\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2088\ : Odrv4
    port map (
            O => \N__13357\,
            I => \Lab_UT.dispString.cntZ0Z_1\
        );

    \I__2087\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13341\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__13341\,
            I => \Lab_UT.dispString.N_166\
        );

    \I__2085\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13335\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__13335\,
            I => \N__13332\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__13332\,
            I => \Lab_UT.dispString.N_167\
        );

    \I__2082\ : InMux
    port map (
            O => \N__13329\,
            I => \N__13326\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__13326\,
            I => \N__13323\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__13323\,
            I => \Lab_UT_dictrl_g1_0_3\
        );

    \I__2079\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13317\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__13317\,
            I => \N__13314\
        );

    \I__2077\ : Span4Mux_s2_v
    port map (
            O => \N__13314\,
            I => \N__13311\
        );

    \I__2076\ : Odrv4
    port map (
            O => \N__13311\,
            I => \uu2.mem0.w_data_2\
        );

    \I__2075\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__13305\,
            I => \Lab_UT.dispString.N_145\
        );

    \I__2073\ : CascadeMux
    port map (
            O => \N__13302\,
            I => \Lab_UT.dispString.N_146_cascade_\
        );

    \I__2072\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13290\
        );

    \I__2071\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13290\
        );

    \I__2070\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13290\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__13290\,
            I => \L3_tx_data_2\
        );

    \I__2068\ : InMux
    port map (
            O => \N__13287\,
            I => \N__13283\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__13286\,
            I => \N__13280\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__13283\,
            I => \N__13276\
        );

    \I__2065\ : InMux
    port map (
            O => \N__13280\,
            I => \N__13271\
        );

    \I__2064\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13271\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__13276\,
            I => \L3_tx_data_0\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__13271\,
            I => \L3_tx_data_0\
        );

    \I__2061\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13262\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13258\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__13262\,
            I => \N__13255\
        );

    \I__2058\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13250\
        );

    \I__2057\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13250\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__13255\,
            I => \L3_tx_data_6\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__13250\,
            I => \L3_tx_data_6\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__13245\,
            I => \Lab_UT.dispString.m82_ns_1_cascade_\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__13242\,
            I => \Lab_UT.dispString.N_156_cascade_\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__13239\,
            I => \N__13235\
        );

    \I__2051\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13231\
        );

    \I__2050\ : InMux
    port map (
            O => \N__13235\,
            I => \N__13226\
        );

    \I__2049\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13226\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__13231\,
            I => \N__13223\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__13226\,
            I => \N__13220\
        );

    \I__2046\ : Odrv12
    port map (
            O => \N__13223\,
            I => \L3_tx_data_3\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__13220\,
            I => \L3_tx_data_3\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__13215\,
            I => \uu2.un1_w_user_lf_0_cascade_\
        );

    \I__2043\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13209\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__13209\,
            I => \uu2.un1_w_user_lfZ0Z_4\
        );

    \I__2041\ : InMux
    port map (
            O => \N__13206\,
            I => \N__13203\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__13203\,
            I => \uu2.un1_w_user_lf_0\
        );

    \I__2039\ : InMux
    port map (
            O => \N__13200\,
            I => \N__13197\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__13197\,
            I => \N__13194\
        );

    \I__2037\ : Span4Mux_s0_v
    port map (
            O => \N__13194\,
            I => \N__13189\
        );

    \I__2036\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13184\
        );

    \I__2035\ : InMux
    port map (
            O => \N__13192\,
            I => \N__13184\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__13189\,
            I => \L3_tx_data_5\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__13184\,
            I => \L3_tx_data_5\
        );

    \I__2032\ : InMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__13176\,
            I => \N__13171\
        );

    \I__2030\ : InMux
    port map (
            O => \N__13175\,
            I => \N__13166\
        );

    \I__2029\ : InMux
    port map (
            O => \N__13174\,
            I => \N__13166\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__13171\,
            I => \L3_tx_data_1\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__13166\,
            I => \L3_tx_data_1\
        );

    \I__2026\ : InMux
    port map (
            O => \N__13161\,
            I => \N__13158\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__13158\,
            I => \N__13153\
        );

    \I__2024\ : InMux
    port map (
            O => \N__13157\,
            I => \N__13148\
        );

    \I__2023\ : InMux
    port map (
            O => \N__13156\,
            I => \N__13148\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__13153\,
            I => \L3_tx_data_4\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__13148\,
            I => \L3_tx_data_4\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__13143\,
            I => \uu2.m35Z0Z_4_cascade_\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__13140\,
            I => \uu2.un1_w_user_cr_0_cascade_\
        );

    \I__2018\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13134\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__13134\,
            I => \N__13131\
        );

    \I__2016\ : Odrv4
    port map (
            O => \N__13131\,
            I => \uu2.mem0.N_69_i\
        );

    \I__2015\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13122\
        );

    \I__2014\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13122\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__13122\,
            I => \uu2.N_96_mux\
        );

    \I__2012\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__13116\,
            I => \N__13113\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__13113\,
            I => \uu2.mem0.N_71_i\
        );

    \I__2009\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13107\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__13107\,
            I => \N__13104\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__13104\,
            I => \uu2.mem0.N_91_mux\
        );

    \I__2006\ : InMux
    port map (
            O => \N__13101\,
            I => \N__13098\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13095\
        );

    \I__2004\ : Span4Mux_s3_h
    port map (
            O => \N__13095\,
            I => \N__13092\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__13092\,
            I => \uu2.mem0.N_50_i\
        );

    \I__2002\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13084\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__13088\,
            I => \N__13081\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__13087\,
            I => \N__13078\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__13084\,
            I => \N__13074\
        );

    \I__1998\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13071\
        );

    \I__1997\ : InMux
    port map (
            O => \N__13078\,
            I => \N__13066\
        );

    \I__1996\ : InMux
    port map (
            O => \N__13077\,
            I => \N__13066\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__13074\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__13071\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__13066\,
            I => \uu2.w_addr_userZ0Z_3\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__13059\,
            I => \N__13056\
        );

    \I__1991\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13053\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__13053\,
            I => \N__13050\
        );

    \I__1989\ : Span4Mux_s1_v
    port map (
            O => \N__13050\,
            I => \N__13047\
        );

    \I__1988\ : Span4Mux_s3_h
    port map (
            O => \N__13047\,
            I => \N__13044\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__13044\,
            I => \uu2.mem0.w_addr_3\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__13041\,
            I => \N__13038\
        );

    \I__1985\ : InMux
    port map (
            O => \N__13038\,
            I => \N__13035\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__13035\,
            I => \N__13032\
        );

    \I__1983\ : Span4Mux_s1_v
    port map (
            O => \N__13032\,
            I => \N__13029\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__13029\,
            I => \uu2.mem0.w_addr_4\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__13026\,
            I => \uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_\
        );

    \I__1980\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13020\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__13020\,
            I => \Lab_UT.dictrl.N_10_1\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__13017\,
            I => \Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__13014\,
            I => \N__13011\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__13011\,
            I => \Lab_UT.dictrl.g0_i_m2_1_1\
        );

    \I__1975\ : InMux
    port map (
            O => \N__13008\,
            I => \N__13005\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__13005\,
            I => \Lab_UT.dictrl.g0_i_m2_1_a6_3_2\
        );

    \I__1973\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12997\
        );

    \I__1972\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12989\
        );

    \I__1971\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12989\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__12997\,
            I => \N__12986\
        );

    \I__1969\ : InMux
    port map (
            O => \N__12996\,
            I => \N__12979\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12995\,
            I => \N__12979\
        );

    \I__1967\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12979\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__12989\,
            I => \N__12976\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__12986\,
            I => bu_rx_data_fast_3
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__12979\,
            I => bu_rx_data_fast_3
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__12976\,
            I => bu_rx_data_fast_3
        );

    \I__1962\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12963\
        );

    \I__1961\ : InMux
    port map (
            O => \N__12968\,
            I => \N__12963\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__12963\,
            I => \Lab_UT.dictrl.N_7_0\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__12960\,
            I => \Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_\
        );

    \I__1958\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12954\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__12954\,
            I => \Lab_UT.dictrl.G_17_i_a5_1\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12948\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12948\,
            I => \N__12945\
        );

    \I__1954\ : Odrv12
    port map (
            O => \N__12945\,
            I => \uu2.mem0.N_66_i\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12939\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__12939\,
            I => \N__12936\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__12936\,
            I => \N__12933\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__12933\,
            I => \uu2.mem0.N_56_i\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__12930\,
            I => \N__12926\
        );

    \I__1948\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12921\
        );

    \I__1947\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12921\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12921\,
            I => \uu2.N_95_mux\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \uu2.N_96_mux_cascade_\
        );

    \I__1944\ : InMux
    port map (
            O => \N__12915\,
            I => \N__12912\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__12912\,
            I => \N__12909\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__12909\,
            I => \N__12906\
        );

    \I__1941\ : Odrv4
    port map (
            O => \N__12906\,
            I => \uu2.mem0.N_63_i\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \N__12900\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12900\,
            I => \N__12897\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__1937\ : Odrv12
    port map (
            O => \N__12894\,
            I => \Lab_UT.dispString.m107_eZ0Z_3\
        );

    \I__1936\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12881\
        );

    \I__1935\ : InMux
    port map (
            O => \N__12890\,
            I => \N__12881\
        );

    \I__1934\ : InMux
    port map (
            O => \N__12889\,
            I => \N__12881\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__12888\,
            I => \N__12878\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__12881\,
            I => \N__12875\
        );

    \I__1931\ : InMux
    port map (
            O => \N__12878\,
            I => \N__12872\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__12875\,
            I => bu_rx_data_fast_5
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__12872\,
            I => bu_rx_data_fast_5
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__12867\,
            I => \Lab_UT.dictrl.N_10_1_cascade_\
        );

    \I__1927\ : InMux
    port map (
            O => \N__12864\,
            I => \N__12861\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__12861\,
            I => \N__12858\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__12858\,
            I => \N__12855\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__12855\,
            I => \Lab_UT.dictrl.N_17_0\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__12852\,
            I => \Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12846\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12846\,
            I => \N__12843\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__12843\,
            I => \N_22\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12837\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__12837\,
            I => \Lab_UT.dictrl.N_1105_0\
        );

    \I__1917\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12830\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__12833\,
            I => \N__12824\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__12830\,
            I => \N__12821\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12818\
        );

    \I__1913\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12811\
        );

    \I__1912\ : InMux
    port map (
            O => \N__12827\,
            I => \N__12811\
        );

    \I__1911\ : InMux
    port map (
            O => \N__12824\,
            I => \N__12811\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__12821\,
            I => bu_rx_data_fast_7
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__12818\,
            I => bu_rx_data_fast_7
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__12811\,
            I => bu_rx_data_fast_7
        );

    \I__1907\ : InMux
    port map (
            O => \N__12804\,
            I => \N__12801\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__12801\,
            I => \buart.Z_rx.G_17_i_a5_2_5\
        );

    \I__1905\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__12795\,
            I => \N__12792\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__12789\,
            I => \buart.Z_rx.G_17_i_a5_2_4\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__12786\,
            I => \G_17_i_a5_2_6_cascade_\
        );

    \I__1900\ : InMux
    port map (
            O => \N__12783\,
            I => \N__12770\
        );

    \I__1899\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12770\
        );

    \I__1898\ : InMux
    port map (
            O => \N__12781\,
            I => \N__12770\
        );

    \I__1897\ : InMux
    port map (
            O => \N__12780\,
            I => \N__12770\
        );

    \I__1896\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12767\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__12770\,
            I => bu_rx_data_fast_1
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__12767\,
            I => bu_rx_data_fast_1
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \N__12758\
        );

    \I__1892\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12755\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12743\
        );

    \I__1890\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12743\
        );

    \I__1889\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12743\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12743\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12740\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__12743\,
            I => bu_rx_data_fast_2
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__12740\,
            I => bu_rx_data_fast_2
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \Lab_UT.dictrl.g2_0_3_0_cascade_\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__12729\,
            I => \Lab_UT.dictrl.g2_0_4_0\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__12726\,
            I => \N__12722\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12718\
        );

    \I__1879\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12713\
        );

    \I__1878\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12713\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12718\,
            I => \N__12705\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__12713\,
            I => \N__12702\
        );

    \I__1875\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12691\
        );

    \I__1874\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12691\
        );

    \I__1873\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12691\
        );

    \I__1872\ : InMux
    port map (
            O => \N__12709\,
            I => \N__12691\
        );

    \I__1871\ : InMux
    port map (
            O => \N__12708\,
            I => \N__12691\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__12705\,
            I => bu_rx_data_1_rep1
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__12702\,
            I => bu_rx_data_1_rep1
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__12691\,
            I => bu_rx_data_1_rep1
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__12684\,
            I => \N__12679\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__12683\,
            I => \N__12674\
        );

    \I__1865\ : CascadeMux
    port map (
            O => \N__12682\,
            I => \N__12671\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12661\
        );

    \I__1863\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12661\
        );

    \I__1862\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12661\
        );

    \I__1861\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12650\
        );

    \I__1860\ : InMux
    port map (
            O => \N__12671\,
            I => \N__12650\
        );

    \I__1859\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12650\
        );

    \I__1858\ : InMux
    port map (
            O => \N__12669\,
            I => \N__12650\
        );

    \I__1857\ : InMux
    port map (
            O => \N__12668\,
            I => \N__12650\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__12661\,
            I => \N__12647\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__12650\,
            I => bu_rx_data_2_rep1
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__12647\,
            I => bu_rx_data_2_rep1
        );

    \I__1853\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12639\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__12639\,
            I => \Lab_UT.dictrl.m27_d_1\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__12636\,
            I => \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_\
        );

    \I__1850\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12627\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__12627\,
            I => \Lab_UT.dictrl.G_17_i_a5_0_0\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__12624\,
            I => \N__12621\
        );

    \I__1846\ : InMux
    port map (
            O => \N__12621\,
            I => \N__12618\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__12618\,
            I => \Lab_UT.dictrl.m71Z0Z_0\
        );

    \I__1844\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12599\
        );

    \I__1843\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12599\
        );

    \I__1842\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12599\
        );

    \I__1841\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12599\
        );

    \I__1840\ : InMux
    port map (
            O => \N__12611\,
            I => \N__12590\
        );

    \I__1839\ : InMux
    port map (
            O => \N__12610\,
            I => \N__12590\
        );

    \I__1838\ : InMux
    port map (
            O => \N__12609\,
            I => \N__12590\
        );

    \I__1837\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12590\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__12599\,
            I => \N__12585\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__12590\,
            I => \N__12585\
        );

    \I__1834\ : Span4Mux_h
    port map (
            O => \N__12585\,
            I => \N__12582\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__12582\,
            I => \N_105_mux\
        );

    \I__1832\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12576\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__12576\,
            I => \Lab_UT.dispString.N_186\
        );

    \I__1830\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12570\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__12570\,
            I => \Lab_UT.dictrl.g0_12_a6_3Z0Z_7\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__12567\,
            I => \Lab_UT.dictrl.g0_12_a6_3_8_cascade_\
        );

    \I__1827\ : InMux
    port map (
            O => \N__12564\,
            I => \N__12561\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__12561\,
            I => \Lab_UT.dictrl.N_16\
        );

    \I__1825\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12555\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__12555\,
            I => \N_10_2\
        );

    \I__1823\ : InMux
    port map (
            O => \N__12552\,
            I => \N__12549\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__12549\,
            I => \Lab_UT.dictrl.N_97_mux_0_0_0\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__12546\,
            I => \Lab_UT.dictrl.g0_10_1_cascade_\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__1819\ : InMux
    port map (
            O => \N__12540\,
            I => \N__12537\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__12534\,
            I => \N__12531\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__12531\,
            I => \Lab_UT.dictrl.m63_d_0_ns_1_1\
        );

    \I__1815\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12524\
        );

    \I__1814\ : InMux
    port map (
            O => \N__12527\,
            I => \N__12521\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__12524\,
            I => \N__12518\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__12521\,
            I => \N__12515\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__12518\,
            I => \Lab_UT.dispString.N_112_mux\
        );

    \I__1810\ : Odrv4
    port map (
            O => \N__12515\,
            I => \Lab_UT.dispString.N_112_mux\
        );

    \I__1809\ : InMux
    port map (
            O => \N__12510\,
            I => \N__12507\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__12507\,
            I => \uu0.sec_clkDZ0\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__12504\,
            I => \Lab_UT.alarmstate_1_0_i_1_cascade_\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__12501\,
            I => \G_215_cascade_\
        );

    \I__1805\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12495\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__12495\,
            I => \G_214\
        );

    \I__1803\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12486\
        );

    \I__1802\ : InMux
    port map (
            O => \N__12491\,
            I => \N__12486\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__12486\,
            I => \G_216\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__12483\,
            I => \G_214_cascade_\
        );

    \I__1799\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12477\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__12477\,
            I => \Lab_UT.m57\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__12474\,
            I => \N__12470\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__12473\,
            I => \N__12464\
        );

    \I__1795\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12455\
        );

    \I__1794\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12455\
        );

    \I__1793\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12455\
        );

    \I__1792\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12455\
        );

    \I__1791\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12447\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__12455\,
            I => \N__12444\
        );

    \I__1789\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12441\
        );

    \I__1788\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12432\
        );

    \I__1787\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12432\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12451\,
            I => \N__12432\
        );

    \I__1785\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12432\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12447\,
            I => \G_213\
        );

    \I__1783\ : Odrv4
    port map (
            O => \N__12444\,
            I => \G_213\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__12441\,
            I => \G_213\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__12432\,
            I => \G_213\
        );

    \I__1780\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12409\
        );

    \I__1779\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12409\
        );

    \I__1778\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12409\
        );

    \I__1777\ : InMux
    port map (
            O => \N__12420\,
            I => \N__12409\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__12419\,
            I => \N__12403\
        );

    \I__1775\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12399\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__12409\,
            I => \N__12396\
        );

    \I__1773\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12393\
        );

    \I__1772\ : InMux
    port map (
            O => \N__12407\,
            I => \N__12384\
        );

    \I__1771\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12384\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12403\,
            I => \N__12384\
        );

    \I__1769\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12384\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__12399\,
            I => \G_215\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__12396\,
            I => \G_215\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__12393\,
            I => \G_215\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__12384\,
            I => \G_215\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__12375\,
            I => \G_213_cascade_\
        );

    \I__1763\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12365\
        );

    \I__1762\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12365\
        );

    \I__1761\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12362\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__12365\,
            I => \N__12359\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__12362\,
            I => \uu0.un88_ci_3\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__12359\,
            I => \uu0.un88_ci_3\
        );

    \I__1757\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12351\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__12351\,
            I => \N__12347\
        );

    \I__1755\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12342\
        );

    \I__1754\ : Span4Mux_h
    port map (
            O => \N__12347\,
            I => \N__12339\
        );

    \I__1753\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12334\
        );

    \I__1752\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12334\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__12342\,
            I => \N__12331\
        );

    \I__1750\ : Odrv4
    port map (
            O => \N__12339\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__12334\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__12331\,
            I => \uu0.l_countZ0Z_6\
        );

    \I__1747\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12321\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__12321\,
            I => \N__12318\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__12318\,
            I => \uu0.un99_ci_0\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__1743\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12309\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__12309\,
            I => \Lab_UT.dispString.dOutP_0_iv_2_tz_1\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__12306\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_\
        );

    \I__1740\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__12300\,
            I => \Lab_UT.dispString.dOutP_0_iv_1_1_1\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__12297\,
            I => \N__12294\
        );

    \I__1737\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12291\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__12291\,
            I => \Lab_UT.dispString.m74_ns_1\
        );

    \I__1735\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12285\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__12285\,
            I => \Lab_UT.dispString.m77_ns_1\
        );

    \I__1733\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12278\
        );

    \I__1732\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12275\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12270\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12270\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__12270\,
            I => \Lab_UT.dispString.N_30_i\
        );

    \I__1728\ : InMux
    port map (
            O => \N__12267\,
            I => \N__12264\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__12264\,
            I => \Lab_UT.dispString.dOutP_0_iv_0_1\
        );

    \I__1726\ : InMux
    port map (
            O => \N__12261\,
            I => \N__12258\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__12258\,
            I => \N__12254\
        );

    \I__1724\ : InMux
    port map (
            O => \N__12257\,
            I => \N__12250\
        );

    \I__1723\ : Span4Mux_h
    port map (
            O => \N__12254\,
            I => \N__12247\
        );

    \I__1722\ : InMux
    port map (
            O => \N__12253\,
            I => \N__12244\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__12250\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1720\ : Odrv4
    port map (
            O => \N__12247\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__12244\,
            I => \uu0.l_countZ0Z_5\
        );

    \I__1718\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12233\
        );

    \I__1717\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12230\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__12233\,
            I => \N__12227\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12222\
        );

    \I__1714\ : Span4Mux_h
    port map (
            O => \N__12227\,
            I => \N__12219\
        );

    \I__1713\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12214\
        );

    \I__1712\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12214\
        );

    \I__1711\ : Odrv12
    port map (
            O => \N__12222\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__12219\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__12214\,
            I => \uu0.l_countZ0Z_4\
        );

    \I__1708\ : InMux
    port map (
            O => \N__12207\,
            I => \N__12201\
        );

    \I__1707\ : InMux
    port map (
            O => \N__12206\,
            I => \N__12201\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__12201\,
            I => \uu2.un284_ci\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__12198\,
            I => \N__12195\
        );

    \I__1704\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12186\
        );

    \I__1703\ : InMux
    port map (
            O => \N__12194\,
            I => \N__12186\
        );

    \I__1702\ : InMux
    port map (
            O => \N__12193\,
            I => \N__12179\
        );

    \I__1701\ : InMux
    port map (
            O => \N__12192\,
            I => \N__12179\
        );

    \I__1700\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12179\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__12186\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__12179\,
            I => \uu2.l_countZ0Z_1\
        );

    \I__1697\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12162\
        );

    \I__1696\ : InMux
    port map (
            O => \N__12173\,
            I => \N__12162\
        );

    \I__1695\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12162\
        );

    \I__1694\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12159\
        );

    \I__1693\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12154\
        );

    \I__1692\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12154\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__12162\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__12159\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__12154\,
            I => \uu2.l_countZ0Z_0\
        );

    \I__1688\ : CEMux
    port map (
            O => \N__12147\,
            I => \N__12144\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12141\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__12141\,
            I => \uu2.un28_w_addr_user_i_0\
        );

    \I__1685\ : InMux
    port map (
            O => \N__12138\,
            I => \N__12134\
        );

    \I__1684\ : InMux
    port map (
            O => \N__12137\,
            I => \N__12131\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__12134\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__12131\,
            I => \uu2.un1_l_count_1_0\
        );

    \I__1681\ : InMux
    port map (
            O => \N__12126\,
            I => \N__12099\
        );

    \I__1680\ : InMux
    port map (
            O => \N__12125\,
            I => \N__12099\
        );

    \I__1679\ : InMux
    port map (
            O => \N__12124\,
            I => \N__12099\
        );

    \I__1678\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12099\
        );

    \I__1677\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12099\
        );

    \I__1676\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12099\
        );

    \I__1675\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12099\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__12119\,
            I => \N__12095\
        );

    \I__1673\ : InMux
    port map (
            O => \N__12118\,
            I => \N__12084\
        );

    \I__1672\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12084\
        );

    \I__1671\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12084\
        );

    \I__1670\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12084\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__12114\,
            I => \N__12081\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__12099\,
            I => \N__12078\
        );

    \I__1667\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12069\
        );

    \I__1666\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12069\
        );

    \I__1665\ : InMux
    port map (
            O => \N__12094\,
            I => \N__12069\
        );

    \I__1664\ : InMux
    port map (
            O => \N__12093\,
            I => \N__12069\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__12084\,
            I => \N__12066\
        );

    \I__1662\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12063\
        );

    \I__1661\ : Span4Mux_h
    port map (
            O => \N__12078\,
            I => \N__12056\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__12069\,
            I => \N__12056\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__12066\,
            I => \N__12056\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__12063\,
            I => vbuf_tx_data_rdy
        );

    \I__1657\ : Odrv4
    port map (
            O => \N__12056\,
            I => vbuf_tx_data_rdy
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__12048\,
            I => \N__12044\
        );

    \I__1654\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12028\
        );

    \I__1653\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12028\
        );

    \I__1652\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12028\
        );

    \I__1651\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12028\
        );

    \I__1650\ : InMux
    port map (
            O => \N__12041\,
            I => \N__12028\
        );

    \I__1649\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12023\
        );

    \I__1648\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12023\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__12028\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__12023\,
            I => \uu2.w_addr_userZ0Z_0\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__12018\,
            I => \uu2.un426_ci_3_cascade_\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__12015\,
            I => \N__12011\
        );

    \I__1643\ : InMux
    port map (
            O => \N__12014\,
            I => \N__12008\
        );

    \I__1642\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12002\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__12008\,
            I => \N__11999\
        );

    \I__1640\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11996\
        );

    \I__1639\ : InMux
    port map (
            O => \N__12006\,
            I => \N__11991\
        );

    \I__1638\ : InMux
    port map (
            O => \N__12005\,
            I => \N__11991\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__12002\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__11999\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__11996\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__11991\,
            I => \uu2.r_addrZ0Z_4\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11982\,
            I => \N__11979\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11979\,
            I => \N__11973\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11970\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11965\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11965\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__11973\,
            I => \uu2.un404_ci_0\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__11970\,
            I => \uu2.un404_ci_0\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__11965\,
            I => \uu2.un404_ci_0\
        );

    \I__1625\ : InMux
    port map (
            O => \N__11958\,
            I => \N__11951\
        );

    \I__1624\ : InMux
    port map (
            O => \N__11957\,
            I => \N__11942\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11956\,
            I => \N__11942\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11942\
        );

    \I__1621\ : InMux
    port map (
            O => \N__11954\,
            I => \N__11942\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11951\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__11942\,
            I => \uu2.trig_rd_is_det\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__11937\,
            I => \N__11934\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11934\,
            I => \N__11931\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__11930\,
            I => \N__11922\
        );

    \I__1614\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11917\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11917\
        );

    \I__1612\ : Span4Mux_s2_v
    port map (
            O => \N__11925\,
            I => \N__11914\
        );

    \I__1611\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11911\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__11917\,
            I => \N__11908\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__11914\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__11911\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__11908\,
            I => \uu2.r_addrZ0Z_5\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__11898\,
            I => \Lab_UT.dictrl.g1_5_0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__11892\,
            I => \Lab_UT.dictrl.N_97_mux_0\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__11889\,
            I => \Lab_UT.dictrl.g0_16_2_cascade_\
        );

    \I__1601\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11883\,
            I => \N__11880\
        );

    \I__1599\ : Span4Mux_v
    port map (
            O => \N__11880\,
            I => \N__11877\
        );

    \I__1598\ : Odrv4
    port map (
            O => \N__11877\,
            I => \Lab_UT.dictrl.N_2446_1\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__11874\,
            I => \N__11871\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11871\,
            I => \N__11868\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__11868\,
            I => \N__11865\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__11865\,
            I => \uu2.mem0.w_addr_0\
        );

    \I__1593\ : IoInMux
    port map (
            O => \N__11862\,
            I => \N__11859\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__1591\ : Span12Mux_s9_v
    port map (
            O => \N__11856\,
            I => \N__11852\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11849\
        );

    \I__1589\ : Odrv12
    port map (
            O => \N__11852\,
            I => clk
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__11849\,
            I => clk
        );

    \I__1587\ : SRMux
    port map (
            O => \N__11844\,
            I => \N__11841\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__11841\,
            I => \N__11837\
        );

    \I__1585\ : CEMux
    port map (
            O => \N__11840\,
            I => \N__11834\
        );

    \I__1584\ : Span4Mux_h
    port map (
            O => \N__11837\,
            I => \N__11831\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11828\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__11831\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__11828\,
            I => \uu2.vram_wr_en_0_iZ0\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__11823\,
            I => \N__11820\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11817\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__11817\,
            I => \N__11814\
        );

    \I__1577\ : Odrv4
    port map (
            O => \N__11814\,
            I => \uu2.mem0.w_addr_1\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__11811\,
            I => \N__11808\
        );

    \I__1575\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11805\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__11805\,
            I => \N__11802\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__11802\,
            I => \uu2.mem0.w_addr_2\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__11799\,
            I => \Lab_UT.dictrl.m40Z0Z_1_cascade_\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11793\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11793\,
            I => \N__11790\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__11790\,
            I => \N__11787\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__11787\,
            I => \Lab_UT.dictrl.N_10_3\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \Lab_UT.dictrl.N_5_0_cascade_\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__1565\ : InMux
    port map (
            O => \N__11778\,
            I => \N__11775\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__11775\,
            I => \Lab_UT.dictrl.g0_9Z0Z_3\
        );

    \I__1563\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__1561\ : Odrv12
    port map (
            O => \N__11766\,
            I => \Lab_UT.dictrl.g1_4\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__11763\,
            I => \Lab_UT.dictrl.N_97_mux_0_cascade_\
        );

    \I__1559\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__1557\ : Span4Mux_s3_h
    port map (
            O => \N__11754\,
            I => \N__11751\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__11751\,
            I => \Lab_UT.dictrl.N_2435_0\
        );

    \I__1555\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11745\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11742\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__11742\,
            I => \N__11737\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11730\
        );

    \I__1551\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11730\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__11737\,
            I => \N__11727\
        );

    \I__1549\ : InMux
    port map (
            O => \N__11736\,
            I => \N__11722\
        );

    \I__1548\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11722\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__11730\,
            I => \N__11719\
        );

    \I__1546\ : Odrv4
    port map (
            O => \N__11727\,
            I => \buart__rx_hh_1\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__11722\,
            I => \buart__rx_hh_1\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__11719\,
            I => \buart__rx_hh_1\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__11706\,
            I => \Lab_UT.dictrl.g0_12_o6_2_2\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__11703\,
            I => \Lab_UT.dictrl.N_13_0_cascade_\
        );

    \I__1539\ : InMux
    port map (
            O => \N__11700\,
            I => \N__11697\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__11697\,
            I => \Lab_UT.dictrl.g0_10Z0Z_3\
        );

    \I__1537\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11691\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__11691\,
            I => \Lab_UT.dictrl.m34_4Z0Z_2\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__11688\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\
        );

    \I__1534\ : CascadeMux
    port map (
            O => \N__11685\,
            I => \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__11682\,
            I => \N__11677\
        );

    \I__1532\ : InMux
    port map (
            O => \N__11681\,
            I => \N__11672\
        );

    \I__1531\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11672\
        );

    \I__1530\ : InMux
    port map (
            O => \N__11677\,
            I => \N__11669\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__11672\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__11669\,
            I => \buart.Z_tx.bitcountZ0Z_2\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \N__11660\
        );

    \I__1526\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11649\
        );

    \I__1525\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11649\
        );

    \I__1524\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11649\
        );

    \I__1523\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11649\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__11649\,
            I => \buart.Z_tx.bitcountZ0Z_1\
        );

    \I__1521\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11639\
        );

    \I__1520\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11636\
        );

    \I__1519\ : InMux
    port map (
            O => \N__11644\,
            I => \N__11629\
        );

    \I__1518\ : InMux
    port map (
            O => \N__11643\,
            I => \N__11629\
        );

    \I__1517\ : InMux
    port map (
            O => \N__11642\,
            I => \N__11629\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__11639\,
            I => \N__11626\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__11636\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__11629\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__11626\,
            I => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\
        );

    \I__1512\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11604\
        );

    \I__1511\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11604\
        );

    \I__1510\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11604\
        );

    \I__1509\ : InMux
    port map (
            O => \N__11616\,
            I => \N__11604\
        );

    \I__1508\ : InMux
    port map (
            O => \N__11615\,
            I => \N__11604\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__11604\,
            I => \buart.Z_tx.bitcountZ0Z_0\
        );

    \I__1506\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11588\
        );

    \I__1505\ : InMux
    port map (
            O => \N__11600\,
            I => \N__11588\
        );

    \I__1504\ : InMux
    port map (
            O => \N__11599\,
            I => \N__11588\
        );

    \I__1503\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11578\
        );

    \I__1502\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11578\
        );

    \I__1501\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11573\
        );

    \I__1500\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11573\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__11588\,
            I => \N__11570\
        );

    \I__1498\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11563\
        );

    \I__1497\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11563\
        );

    \I__1496\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11563\
        );

    \I__1495\ : InMux
    port map (
            O => \N__11584\,
            I => \N__11558\
        );

    \I__1494\ : InMux
    port map (
            O => \N__11583\,
            I => \N__11558\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__11578\,
            I => \N__11555\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__11573\,
            I => \uu0.un4_l_count_0\
        );

    \I__1491\ : Odrv4
    port map (
            O => \N__11570\,
            I => \uu0.un4_l_count_0\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__11563\,
            I => \uu0.un4_l_count_0\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__11558\,
            I => \uu0.un4_l_count_0\
        );

    \I__1488\ : Odrv4
    port map (
            O => \N__11555\,
            I => \uu0.un4_l_count_0\
        );

    \I__1487\ : IoInMux
    port map (
            O => \N__11544\,
            I => \N__11541\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__11541\,
            I => \N__11538\
        );

    \I__1485\ : IoSpan4Mux
    port map (
            O => \N__11538\,
            I => \N__11535\
        );

    \I__1484\ : Span4Mux_s0_h
    port map (
            O => \N__11535\,
            I => \N__11532\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__11532\,
            I => \uu0.un11_l_count_i\
        );

    \I__1482\ : InMux
    port map (
            O => \N__11529\,
            I => \N__11523\
        );

    \I__1481\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11523\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__11523\,
            I => \N__11520\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__11517\,
            I => \uu0.delay_lineZ0Z_0\
        );

    \I__1477\ : InMux
    port map (
            O => \N__11514\,
            I => \N__11511\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__11511\,
            I => \uu0.delay_lineZ0Z_1\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__11508\,
            I => \buart.Z_tx.un1_bitcount_c3_cascade_\
        );

    \I__1474\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11499\
        );

    \I__1473\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11499\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__11499\,
            I => \buart.Z_tx.bitcountZ0Z_3\
        );

    \I__1471\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11493\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__11493\,
            I => \buart.Z_tx.uart_busy_0_0\
        );

    \I__1469\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11484\
        );

    \I__1468\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11477\
        );

    \I__1467\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11477\
        );

    \I__1466\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11477\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11474\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__11477\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1463\ : Odrv4
    port map (
            O => \N__11474\,
            I => \buart.Z_tx.ser_clk\
        );

    \I__1462\ : CascadeMux
    port map (
            O => \N__11469\,
            I => \N__11466\
        );

    \I__1461\ : InMux
    port map (
            O => \N__11466\,
            I => \N__11463\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__11463\,
            I => \uu2.un1_l_count_1_2_0\
        );

    \I__1459\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11455\
        );

    \I__1458\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11452\
        );

    \I__1457\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11449\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__11455\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__11452\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__11449\,
            I => \uu2.l_countZ0Z_5\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__11442\,
            I => \uu2.vbuf_count.un328_ci_3_cascade_\
        );

    \I__1452\ : InMux
    port map (
            O => \N__11439\,
            I => \N__11436\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__11436\,
            I => \N__11431\
        );

    \I__1450\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11428\
        );

    \I__1449\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11425\
        );

    \I__1448\ : Span4Mux_s3_h
    port map (
            O => \N__11431\,
            I => \N__11422\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__11428\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__11425\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__11422\,
            I => \uu2.un1_l_count_2_0\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \uu2.un350_ci_cascade_\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \N__11405\
        );

    \I__1442\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11400\
        );

    \I__1441\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11400\
        );

    \I__1440\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11393\
        );

    \I__1439\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11393\
        );

    \I__1438\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11393\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__11400\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__11393\,
            I => \uu2.l_countZ0Z_4\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__11388\,
            I => \N__11383\
        );

    \I__1434\ : InMux
    port map (
            O => \N__11387\,
            I => \N__11376\
        );

    \I__1433\ : InMux
    port map (
            O => \N__11386\,
            I => \N__11376\
        );

    \I__1432\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11376\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__11376\,
            I => \uu2.l_countZ0Z_9\
        );

    \I__1430\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__11370\,
            I => \uu2.un1_l_count_2_2\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__11367\,
            I => \N__11364\
        );

    \I__1427\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11358\
        );

    \I__1426\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11351\
        );

    \I__1425\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11351\
        );

    \I__1424\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11351\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__11358\,
            I => \uu2.un306_ci\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__11351\,
            I => \uu2.un306_ci\
        );

    \I__1421\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11340\
        );

    \I__1420\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11340\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__11340\,
            I => \uu2.vbuf_count.un328_ci_3\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__11337\,
            I => \N__11334\
        );

    \I__1417\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11319\
        );

    \I__1416\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11319\
        );

    \I__1415\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11319\
        );

    \I__1414\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11319\
        );

    \I__1413\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11319\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__11319\,
            I => \uu2.l_countZ0Z_6\
        );

    \I__1411\ : InMux
    port map (
            O => \N__11316\,
            I => \N__11309\
        );

    \I__1410\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11309\
        );

    \I__1409\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11306\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__11309\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__11306\,
            I => \uu2.l_countZ0Z_7\
        );

    \I__1406\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11298\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__11298\,
            I => \uu2.un350_ci\
        );

    \I__1404\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11290\
        );

    \I__1403\ : InMux
    port map (
            O => \N__11294\,
            I => \N__11287\
        );

    \I__1402\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11284\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__11290\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__11287\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__11284\,
            I => \uu2.l_countZ0Z_8\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__11277\,
            I => \uu2.un1_l_count_1_3_cascade_\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__11274\,
            I => \uu2.un1_l_count_2_0_cascade_\
        );

    \I__1396\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__11268\,
            I => \uu2.un1_l_count_1_3\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__11265\,
            I => \N__11260\
        );

    \I__1393\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11255\
        );

    \I__1392\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11255\
        );

    \I__1391\ : InMux
    port map (
            O => \N__11260\,
            I => \N__11252\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__11255\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__11252\,
            I => \uu2.l_countZ0Z_3\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__11247\,
            I => \N__11240\
        );

    \I__1387\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11229\
        );

    \I__1386\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11229\
        );

    \I__1385\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11229\
        );

    \I__1384\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11229\
        );

    \I__1383\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11229\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__11229\,
            I => \uu2.l_countZ0Z_2\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__11226\,
            I => \uu2.un306_ci_cascade_\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__11223\,
            I => \uu2.un404_ci_0_cascade_\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__11220\,
            I => \N__11217\
        );

    \I__1378\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11211\
        );

    \I__1377\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11204\
        );

    \I__1376\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11204\
        );

    \I__1375\ : InMux
    port map (
            O => \N__11214\,
            I => \N__11204\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__11211\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__11204\,
            I => \uu2.r_addrZ0Z_6\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__11199\,
            I => \N__11194\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11191\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__11197\,
            I => \N__11188\
        );

    \I__1369\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11185\
        );

    \I__1368\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11180\
        );

    \I__1367\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11180\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__11185\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__11180\,
            I => \uu2.r_addrZ0Z_3\
        );

    \I__1364\ : CascadeMux
    port map (
            O => \N__11175\,
            I => \N__11171\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__11174\,
            I => \N__11168\
        );

    \I__1362\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11163\
        );

    \I__1361\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11160\
        );

    \I__1360\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11155\
        );

    \I__1359\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11155\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__11163\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__11160\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__11155\,
            I => \uu2.r_addrZ0Z_2\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__11148\,
            I => \N__11145\
        );

    \I__1354\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11142\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11135\
        );

    \I__1352\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11130\
        );

    \I__1351\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11130\
        );

    \I__1350\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11125\
        );

    \I__1349\ : InMux
    port map (
            O => \N__11138\,
            I => \N__11125\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__11135\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__11130\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__11125\,
            I => \uu2.r_addrZ0Z_1\
        );

    \I__1345\ : CEMux
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__11115\,
            I => \uu2.trig_rd_is_det_0\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__11112\,
            I => \uu2.trig_rd_is_det_cascade_\
        );

    \I__1342\ : CascadeMux
    port map (
            O => \N__11109\,
            I => \N__11105\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11101\
        );

    \I__1340\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11095\
        );

    \I__1339\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11088\
        );

    \I__1338\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11088\
        );

    \I__1337\ : InMux
    port map (
            O => \N__11100\,
            I => \N__11088\
        );

    \I__1336\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11083\
        );

    \I__1335\ : InMux
    port map (
            O => \N__11098\,
            I => \N__11083\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__11095\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__11088\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__11083\,
            I => \uu2.r_addrZ0Z_0\
        );

    \I__1331\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11073\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__11073\,
            I => \uu2.trig_rd_detZ0Z_1\
        );

    \I__1329\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11064\
        );

    \I__1328\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11064\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__11064\,
            I => \uu2.trig_rd_detZ0Z_0\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__1325\ : InMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__11052\,
            I => \Lab_UT.dictrl.g1_6_0\
        );

    \I__1322\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11046\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__11046\,
            I => \uu2.vbuf_raddr.un426_ci_3\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__11043\,
            I => \uu2.vbuf_raddr.un426_ci_3_cascade_\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__11040\,
            I => \N__11037\
        );

    \I__1318\ : InMux
    port map (
            O => \N__11037\,
            I => \N__11033\
        );

    \I__1317\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11030\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__11033\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1315\ : LocalMux
    port map (
            O => \N__11030\,
            I => \uu2.r_addrZ0Z_8\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__11025\,
            I => \N__11021\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__11024\,
            I => \N__11018\
        );

    \I__1312\ : InMux
    port map (
            O => \N__11021\,
            I => \N__11014\
        );

    \I__1311\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11009\
        );

    \I__1310\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11009\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__11014\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__11009\,
            I => \uu2.r_addrZ0Z_7\
        );

    \I__1307\ : InMux
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__11001\,
            I => \uu2.vbuf_raddr.un448_ci_0\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \Lab_UT.dictrl.N_1792_1_cascade_\
        );

    \I__1304\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10992\,
            I => \Lab_UT.dictrl.N_1451_0\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__10989\,
            I => \Lab_UT.dictrl.g0_i_a5_2_4_cascade_\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10986\,
            I => \N__10983\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10983\,
            I => \Lab_UT.dictrl.g0_i_a5_2_5\
        );

    \I__1299\ : CascadeMux
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__1298\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__10974\,
            I => \Lab_UT.dictrl.g0_5_3\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10968\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__10968\,
            I => \N__10965\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__10965\,
            I => \Lab_UT.dictrl.g0_5_4\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10962\,
            I => \Lab_UT.dictrl.g0_69_1_cascade_\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10956\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10956\,
            I => \Lab_UT.dictrl.g1_0_3_1\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__10953\,
            I => \Lab_UT.dictrl.g1_5_1_cascade_\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10950\,
            I => \N__10947\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__10947\,
            I => \Lab_UT.dictrl.N_61_1\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10941\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10941\,
            I => \Lab_UT.dictrl.g1_7_0\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10935\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N_107\
        );

    \I__1283\ : CascadeMux
    port map (
            O => \N__10932\,
            I => \m72_cascade_\
        );

    \I__1282\ : InMux
    port map (
            O => \N__10929\,
            I => \N__10923\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10928\,
            I => \N__10923\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__10923\,
            I => \N_105\
        );

    \I__1279\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10914\
        );

    \I__1278\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10914\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__10914\,
            I => \resetGen.reset_countZ0Z_3\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__10911\,
            I => \N__10906\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10898\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10898\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10891\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10891\
        );

    \I__1271\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10891\
        );

    \I__1270\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10888\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__10898\,
            I => \resetGen_reset_count_4\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__10891\,
            I => \resetGen_reset_count_4\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__10888\,
            I => \resetGen_reset_count_4\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__10881\,
            I => \N__10876\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__10880\,
            I => \N__10872\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__10879\,
            I => \N__10869\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10863\
        );

    \I__1262\ : InMux
    port map (
            O => \N__10875\,
            I => \N__10863\
        );

    \I__1261\ : InMux
    port map (
            O => \N__10872\,
            I => \N__10856\
        );

    \I__1260\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10856\
        );

    \I__1259\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10856\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__10863\,
            I => \resetGen_reset_count_0\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__10856\,
            I => \resetGen_reset_count_0\
        );

    \I__1256\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10848\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__10848\,
            I => \N__10843\
        );

    \I__1254\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10838\
        );

    \I__1253\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10838\
        );

    \I__1252\ : Odrv4
    port map (
            O => \N__10843\,
            I => \buart__rx_hh_0\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__10838\,
            I => \buart__rx_hh_0\
        );

    \I__1250\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10830\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__10830\,
            I => \N__10827\
        );

    \I__1248\ : Odrv12
    port map (
            O => \N__10827\,
            I => vbuf_tx_data_6
        );

    \I__1247\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10821\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__10821\,
            I => \buart.Z_tx.shifterZ0Z_7\
        );

    \I__1245\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10815\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10812\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__10812\,
            I => vbuf_tx_data_7
        );

    \I__1242\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10806\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__10806\,
            I => \buart.Z_tx.shifterZ0Z_8\
        );

    \I__1240\ : CEMux
    port map (
            O => \N__10803\,
            I => \N__10800\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10800\,
            I => \N__10797\
        );

    \I__1238\ : Span4Mux_s1_v
    port map (
            O => \N__10797\,
            I => \N__10793\
        );

    \I__1237\ : CEMux
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__10793\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__10790\,
            I => \buart.Z_tx.un1_uart_wr_i_0_i\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10785\,
            I => \N__10781\
        );

    \I__1233\ : InMux
    port map (
            O => \N__10784\,
            I => \N__10778\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10781\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__10778\,
            I => \uu0.l_countZ0Z_13\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__1229\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10760\
        );

    \I__1228\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10760\
        );

    \I__1227\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10760\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10757\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10752\
        );

    \I__1224\ : Span4Mux_s1_h
    port map (
            O => \N__10757\,
            I => \N__10752\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__10752\,
            I => \uu0.un4_l_count_0_8\
        );

    \I__1222\ : InMux
    port map (
            O => \N__10749\,
            I => \N__10746\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__10746\,
            I => \N__10740\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__10745\,
            I => \N__10737\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__10744\,
            I => \N__10734\
        );

    \I__1218\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10731\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__10740\,
            I => \N__10728\
        );

    \I__1216\ : InMux
    port map (
            O => \N__10737\,
            I => \N__10723\
        );

    \I__1215\ : InMux
    port map (
            O => \N__10734\,
            I => \N__10723\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__10731\,
            I => \uu0.un154_ci_9\
        );

    \I__1213\ : Odrv4
    port map (
            O => \N__10728\,
            I => \uu0.un154_ci_9\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10723\,
            I => \uu0.un154_ci_9\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10709\
        );

    \I__1210\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10709\
        );

    \I__1209\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10706\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10703\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__10706\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__1206\ : Odrv4
    port map (
            O => \N__10703\,
            I => \uu0.l_countZ0Z_12\
        );

    \I__1205\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10695\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__10695\,
            I => \uu0.un165_ci_0\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10679\
        );

    \I__1201\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10679\
        );

    \I__1200\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10679\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__10686\,
            I => \resetGen_reset_count_1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__10679\,
            I => \resetGen_reset_count_1\
        );

    \I__1197\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10671\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__10671\,
            I => \uu0.un44_ci\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__10668\,
            I => \N__10665\
        );

    \I__1194\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10662\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__1192\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10651\
        );

    \I__1191\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10651\
        );

    \I__1190\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10648\
        );

    \I__1189\ : Odrv4
    port map (
            O => \N__10656\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__10651\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__10648\,
            I => \uu0.l_countZ0Z_2\
        );

    \I__1186\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10636\
        );

    \I__1185\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10631\
        );

    \I__1184\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10631\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__10636\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__10631\,
            I => \uu0.l_countZ0Z_3\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__10626\,
            I => \N__10620\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__10625\,
            I => \N__10617\
        );

    \I__1179\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10614\
        );

    \I__1178\ : InMux
    port map (
            O => \N__10623\,
            I => \N__10611\
        );

    \I__1177\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10608\
        );

    \I__1176\ : InMux
    port map (
            O => \N__10617\,
            I => \N__10605\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__10614\,
            I => \uu0.un66_ci\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__10611\,
            I => \uu0.un66_ci\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__10608\,
            I => \uu0.un66_ci\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__10605\,
            I => \uu0.un66_ci\
        );

    \I__1171\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10591\
        );

    \I__1170\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10586\
        );

    \I__1169\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10586\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__10591\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__10586\,
            I => \uu0.l_countZ0Z_7\
        );

    \I__1166\ : InMux
    port map (
            O => \N__10581\,
            I => \N__10578\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__10578\,
            I => \uu0.un220_ci\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__10575\,
            I => \N__10572\
        );

    \I__1163\ : InMux
    port map (
            O => \N__10572\,
            I => \N__10569\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__10569\,
            I => \uu0.un143_ci_0\
        );

    \I__1161\ : CascadeMux
    port map (
            O => \N__10566\,
            I => \N__10563\
        );

    \I__1160\ : InMux
    port map (
            O => \N__10563\,
            I => \N__10558\
        );

    \I__1159\ : InMux
    port map (
            O => \N__10562\,
            I => \N__10553\
        );

    \I__1158\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10553\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__10558\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__10553\,
            I => \uu0.l_countZ0Z_11\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10544\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__10547\,
            I => \N__10541\
        );

    \I__1153\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10536\
        );

    \I__1152\ : InMux
    port map (
            O => \N__10541\,
            I => \N__10536\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__10536\,
            I => \uu0.l_countZ0Z_18\
        );

    \I__1150\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10530\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__10530\,
            I => \uu0.un4_l_count_11\
        );

    \I__1148\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10524\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__10524\,
            I => \N__10521\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__10521\,
            I => \uu0.un4_l_count_12\
        );

    \I__1145\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10515\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__10515\,
            I => \uu0.un4_l_count_13\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__10512\,
            I => \uu0.un4_l_count_16_cascade_\
        );

    \I__1142\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10506\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__10506\,
            I => \N__10503\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__10503\,
            I => \uu0.un4_l_count_18\
        );

    \I__1139\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10489\
        );

    \I__1138\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10489\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__10498\,
            I => \N__10484\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__10497\,
            I => \N__10481\
        );

    \I__1135\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10477\
        );

    \I__1134\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10472\
        );

    \I__1133\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10472\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10469\
        );

    \I__1131\ : InMux
    port map (
            O => \N__10488\,
            I => \N__10466\
        );

    \I__1130\ : InMux
    port map (
            O => \N__10487\,
            I => \N__10457\
        );

    \I__1129\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10457\
        );

    \I__1128\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10457\
        );

    \I__1127\ : InMux
    port map (
            O => \N__10480\,
            I => \N__10457\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__10477\,
            I => \uu0.un110_ci\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__10472\,
            I => \uu0.un110_ci\
        );

    \I__1124\ : Odrv12
    port map (
            O => \N__10469\,
            I => \uu0.un110_ci\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__10466\,
            I => \uu0.un110_ci\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__10457\,
            I => \uu0.un110_ci\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__10446\,
            I => \uu0.un4_l_count_0_cascade_\
        );

    \I__1120\ : CEMux
    port map (
            O => \N__10443\,
            I => \N__10428\
        );

    \I__1119\ : CEMux
    port map (
            O => \N__10442\,
            I => \N__10428\
        );

    \I__1118\ : CEMux
    port map (
            O => \N__10441\,
            I => \N__10428\
        );

    \I__1117\ : CEMux
    port map (
            O => \N__10440\,
            I => \N__10428\
        );

    \I__1116\ : CEMux
    port map (
            O => \N__10439\,
            I => \N__10428\
        );

    \I__1115\ : GlobalMux
    port map (
            O => \N__10428\,
            I => \N__10425\
        );

    \I__1114\ : gio2CtrlBuf
    port map (
            O => \N__10425\,
            I => \uu0.un11_l_count_i_g\
        );

    \I__1113\ : InMux
    port map (
            O => \N__10422\,
            I => \N__10419\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__10419\,
            I => \N__10416\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__10416\,
            I => vbuf_tx_data_5
        );

    \I__1110\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10410\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__10410\,
            I => \N__10407\
        );

    \I__1108\ : Odrv12
    port map (
            O => \N__10407\,
            I => \buart.Z_tx.shifterZ0Z_6\
        );

    \I__1107\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10391\
        );

    \I__1106\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10391\
        );

    \I__1105\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10391\
        );

    \I__1104\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10391\
        );

    \I__1103\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10388\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__10391\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__10388\,
            I => \uu0.l_countZ0Z_0\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__10383\,
            I => \N__10378\
        );

    \I__1099\ : InMux
    port map (
            O => \N__10382\,
            I => \N__10370\
        );

    \I__1098\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10370\
        );

    \I__1097\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10370\
        );

    \I__1096\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10367\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__10370\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__10367\,
            I => \uu0.l_countZ0Z_1\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__10362\,
            I => \uu0.un66_ci_cascade_\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10359\,
            I => \uu0.un110_ci_cascade_\
        );

    \I__1091\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10350\
        );

    \I__1090\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10345\
        );

    \I__1089\ : InMux
    port map (
            O => \N__10354\,
            I => \N__10345\
        );

    \I__1088\ : InMux
    port map (
            O => \N__10353\,
            I => \N__10342\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__10350\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__10345\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__10342\,
            I => \uu0.l_countZ0Z_10\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10330\
        );

    \I__1083\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10323\
        );

    \I__1082\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10323\
        );

    \I__1081\ : InMux
    port map (
            O => \N__10330\,
            I => \N__10318\
        );

    \I__1080\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10318\
        );

    \I__1079\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10314\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10311\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10308\
        );

    \I__1076\ : InMux
    port map (
            O => \N__10317\,
            I => \N__10305\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__10314\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1074\ : Odrv4
    port map (
            O => \N__10311\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__10308\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10305\,
            I => \uu0.l_countZ0Z_8\
        );

    \I__1071\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10287\
        );

    \I__1070\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10287\
        );

    \I__1069\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10280\
        );

    \I__1068\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10280\
        );

    \I__1067\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10280\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__10287\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__10280\,
            I => \uu0.l_countZ0Z_9\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__10275\,
            I => \N__10270\
        );

    \I__1063\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10263\
        );

    \I__1062\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10263\
        );

    \I__1061\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10263\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__10263\,
            I => \uu0.l_countZ0Z_17\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__10260\,
            I => \N__10255\
        );

    \I__1058\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10248\
        );

    \I__1057\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10248\
        );

    \I__1056\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10248\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__10248\,
            I => \uu0.un198_ci_2\
        );

    \I__1054\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10235\
        );

    \I__1053\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10235\
        );

    \I__1052\ : InMux
    port map (
            O => \N__10243\,
            I => \N__10235\
        );

    \I__1051\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10232\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__10235\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__10232\,
            I => \uu0.l_countZ0Z_16\
        );

    \I__1048\ : InMux
    port map (
            O => \N__10227\,
            I => \N__10224\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__10224\,
            I => vbuf_tx_data_1
        );

    \I__1046\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10218\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__10218\,
            I => \buart.Z_tx.shifterZ0Z_2\
        );

    \I__1044\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10212\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__10212\,
            I => vbuf_tx_data_2
        );

    \I__1042\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__10206\,
            I => \buart.Z_tx.shifterZ0Z_3\
        );

    \I__1040\ : InMux
    port map (
            O => \N__10203\,
            I => \N__10200\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__10200\,
            I => vbuf_tx_data_3
        );

    \I__1038\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__10194\,
            I => \buart.Z_tx.shifterZ0Z_4\
        );

    \I__1036\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10188\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__10188\,
            I => vbuf_tx_data_4
        );

    \I__1034\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10182\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__10182\,
            I => \buart.Z_tx.shifterZ0Z_5\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__10179\,
            I => \uu0.un44_ci_cascade_\
        );

    \I__1031\ : InMux
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__10173\,
            I => \uu2.r_data_wire_2\
        );

    \I__1029\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10167\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__10167\,
            I => \uu2.r_data_wire_3\
        );

    \I__1027\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10161\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__10161\,
            I => \uu2.r_data_wire_4\
        );

    \I__1025\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__10155\,
            I => \uu2.r_data_wire_5\
        );

    \I__1023\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10149\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__10149\,
            I => \uu2.r_data_wire_6\
        );

    \I__1021\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__10143\,
            I => \uu2.r_data_wire_7\
        );

    \I__1019\ : InMux
    port map (
            O => \N__10140\,
            I => \N__10137\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__10137\,
            I => vbuf_tx_data_0
        );

    \I__1017\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10131\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__10131\,
            I => \buart.Z_tx.shifterZ0Z_1\
        );

    \I__1015\ : InMux
    port map (
            O => \N__10128\,
            I => \N__10125\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__10125\,
            I => \buart.Z_tx.shifterZ0Z_0\
        );

    \I__1013\ : IoInMux
    port map (
            O => \N__10122\,
            I => \N__10119\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__10119\,
            I => \N__10116\
        );

    \I__1011\ : Span12Mux_s1_h
    port map (
            O => \N__10116\,
            I => \N__10113\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__10113\,
            I => o_serial_data_c
        );

    \I__1009\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10105\
        );

    \I__1008\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10100\
        );

    \I__1007\ : InMux
    port map (
            O => \N__10108\,
            I => \N__10100\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__10105\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__10100\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_1\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__1003\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10086\
        );

    \I__1002\ : InMux
    port map (
            O => \N__10091\,
            I => \N__10079\
        );

    \I__1001\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10079\
        );

    \I__1000\ : InMux
    port map (
            O => \N__10089\,
            I => \N__10079\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__10086\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__10079\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_0\
        );

    \I__997\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10069\
        );

    \I__996\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10064\
        );

    \I__995\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10064\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__10069\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__10064\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_2\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__10059\,
            I => \N__10056\
        );

    \I__991\ : InMux
    port map (
            O => \N__10056\,
            I => \N__10053\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__10053\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\
        );

    \I__989\ : InMux
    port map (
            O => \N__10050\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\
        );

    \I__988\ : InMux
    port map (
            O => \N__10047\,
            I => \N__10043\
        );

    \I__987\ : InMux
    port map (
            O => \N__10046\,
            I => \N__10040\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__10043\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__10040\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_3\
        );

    \I__984\ : InMux
    port map (
            O => \N__10035\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__10032\,
            I => \N__10028\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__10031\,
            I => \N__10024\
        );

    \I__981\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10021\
        );

    \I__980\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10018\
        );

    \I__979\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10015\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__10021\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__10018\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__10015\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_4\
        );

    \I__975\ : InMux
    port map (
            O => \N__10008\,
            I => \N__10005\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__10005\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\
        );

    \I__973\ : InMux
    port map (
            O => \N__10002\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\
        );

    \I__972\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9990\
        );

    \I__971\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9990\
        );

    \I__970\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9985\
        );

    \I__969\ : InMux
    port map (
            O => \N__9996\,
            I => \N__9985\
        );

    \I__968\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9982\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__9990\,
            I => \N__9979\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9985\,
            I => \buart__rx_ser_clk\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9982\,
            I => \buart__rx_ser_clk\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__9979\,
            I => \buart__rx_ser_clk\
        );

    \I__963\ : InMux
    port map (
            O => \N__9972\,
            I => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__9969\,
            I => \N__9966\
        );

    \I__961\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9962\
        );

    \I__960\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9959\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9962\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9959\,
            I => \buart.Z_rx.Z_baudgen.counterZ0Z_5\
        );

    \I__957\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9951\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9951\,
            I => \uu2.r_data_wire_0\
        );

    \I__955\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9945\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9945\,
            I => \uu2.r_data_wire_1\
        );

    \I__953\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9939\,
            I => \uart_RXD\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__9936\,
            I => \N__9932\
        );

    \I__950\ : InMux
    port map (
            O => \N__9935\,
            I => \N__9927\
        );

    \I__949\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9927\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__9927\,
            I => \Lab_UT.dispString.N_115_mux\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__9924\,
            I => \Lab_UT.dispString.N_115_mux_cascade_\
        );

    \I__946\ : InMux
    port map (
            O => \N__9921\,
            I => \N__9914\
        );

    \I__945\ : InMux
    port map (
            O => \N__9920\,
            I => \N__9911\
        );

    \I__944\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9904\
        );

    \I__943\ : InMux
    port map (
            O => \N__9918\,
            I => \N__9904\
        );

    \I__942\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9904\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9914\,
            I => \buart__rx_bitcount_1\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9911\,
            I => \buart__rx_bitcount_1\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__9904\,
            I => \buart__rx_bitcount_1\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__9897\,
            I => \N__9892\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \N__9888\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__9895\,
            I => \N__9885\
        );

    \I__935\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9878\
        );

    \I__934\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9878\
        );

    \I__933\ : InMux
    port map (
            O => \N__9888\,
            I => \N__9878\
        );

    \I__932\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9875\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__9878\,
            I => \N__9872\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__9875\,
            I => \buart__rx_bitcount_4\
        );

    \I__929\ : Odrv4
    port map (
            O => \N__9872\,
            I => \buart__rx_bitcount_4\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__9867\,
            I => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\
        );

    \I__927\ : InMux
    port map (
            O => \N__9864\,
            I => \N__9861\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9861\,
            I => \Lab_UT.dispString.N_177\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \buart__rx_ser_clk_cascade_\
        );

    \I__924\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9851\
        );

    \I__923\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9845\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__9851\,
            I => \N__9842\
        );

    \I__921\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9839\
        );

    \I__920\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9834\
        );

    \I__919\ : InMux
    port map (
            O => \N__9848\,
            I => \N__9834\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9845\,
            I => \buart__rx_bitcount_0\
        );

    \I__917\ : Odrv4
    port map (
            O => \N__9842\,
            I => \buart__rx_bitcount_0\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9839\,
            I => \buart__rx_bitcount_0\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__9834\,
            I => \buart__rx_bitcount_0\
        );

    \I__914\ : IoInMux
    port map (
            O => \N__9825\,
            I => \N__9822\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__9822\,
            I => \N__9819\
        );

    \I__912\ : IoSpan4Mux
    port map (
            O => \N__9819\,
            I => \N__9816\
        );

    \I__911\ : Span4Mux_s0_v
    port map (
            O => \N__9816\,
            I => \N__9813\
        );

    \I__910\ : Span4Mux_v
    port map (
            O => \N__9813\,
            I => \N__9810\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__9810\,
            I => \buart__rx_sample\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__907\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9801\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__9801\,
            I => \buart.Z_rx.bitcount_cry_2_THRU_CO\
        );

    \I__905\ : InMux
    port map (
            O => \N__9798\,
            I => \buart.Z_rx.bitcount_cry_2\
        );

    \I__904\ : InMux
    port map (
            O => \N__9795\,
            I => \buart.Z_rx.bitcount_cry_3\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__9792\,
            I => \Lab_UT_dispString_m103_ns_1_cascade_\
        );

    \I__902\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9786\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__9786\,
            I => \buart.Z_rx.bitcount_cry_0_THRU_CO\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__9783\,
            I => \buart__rx_N_27_0_i_cascade_\
        );

    \I__899\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__9774\,
            I => \N_179\
        );

    \I__896\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9765\
        );

    \I__895\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9758\
        );

    \I__894\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9758\
        );

    \I__893\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9758\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__9765\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__9758\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_0\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__9753\,
            I => \resetGen_reset_count_2_2_cascade_\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__9750\,
            I => \N__9744\
        );

    \I__888\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9735\
        );

    \I__887\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9735\
        );

    \I__886\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9735\
        );

    \I__885\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9735\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__9735\,
            I => \resetGen_reset_count_2\
        );

    \I__883\ : InMux
    port map (
            O => \N__9732\,
            I => \buart.Z_rx.bitcount_cry_0\
        );

    \I__882\ : InMux
    port map (
            O => \N__9729\,
            I => \buart.Z_rx.bitcount_cry_1\
        );

    \I__881\ : InMux
    port map (
            O => \N__9726\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\
        );

    \I__880\ : InMux
    port map (
            O => \N__9723\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\
        );

    \I__879\ : InMux
    port map (
            O => \N__9720\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\
        );

    \I__878\ : InMux
    port map (
            O => \N__9717\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\
        );

    \I__877\ : InMux
    port map (
            O => \N__9714\,
            I => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\
        );

    \I__876\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9705\
        );

    \I__875\ : InMux
    port map (
            O => \N__9710\,
            I => \N__9705\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__9705\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_5\
        );

    \I__873\ : InMux
    port map (
            O => \N__9702\,
            I => \N__9696\
        );

    \I__872\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9696\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__9696\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_4\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__9693\,
            I => \N__9689\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__9692\,
            I => \N__9686\
        );

    \I__868\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9681\
        );

    \I__867\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9681\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__9681\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_6\
        );

    \I__865\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9672\
        );

    \I__864\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9672\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__9672\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_2\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__9669\,
            I => \N__9665\
        );

    \I__861\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9662\
        );

    \I__860\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9659\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__9662\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__9659\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_3\
        );

    \I__857\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9651\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__9651\,
            I => \buart.Z_tx.Z_baudgen.ser_clk_4\
        );

    \I__855\ : CascadeMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__854\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9640\
        );

    \I__853\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9635\
        );

    \I__852\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9635\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__9640\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__9635\,
            I => \buart.Z_tx.Z_baudgen.counterZ0Z_1\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__9630\,
            I => \N__9627\
        );

    \I__848\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9615\
        );

    \I__847\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9615\
        );

    \I__846\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9615\
        );

    \I__845\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9610\
        );

    \I__844\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9610\
        );

    \I__843\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9607\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__9615\,
            I => \N__9602\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__9610\,
            I => \N__9602\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__9607\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__9602\,
            I => \uu0.l_precountZ0Z_0\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__9597\,
            I => \uu0.un4_l_count_14_cascade_\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__9594\,
            I => \uu0.un154_ci_9_cascade_\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__9591\,
            I => \uu0.un187_ci_1_cascade_\
        );

    \I__835\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9576\
        );

    \I__834\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9576\
        );

    \I__833\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9576\
        );

    \I__832\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9576\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__9576\,
            I => \uu0.l_countZ0Z_14\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__9573\,
            I => \N__9568\
        );

    \I__829\ : InMux
    port map (
            O => \N__9572\,
            I => \N__9561\
        );

    \I__828\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9561\
        );

    \I__827\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9561\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__9561\,
            I => \uu0.l_countZ0Z_15\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__9558\,
            I => \N__9553\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__9557\,
            I => \N__9550\
        );

    \I__823\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9543\
        );

    \I__822\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9543\
        );

    \I__821\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9543\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__9543\,
            I => \uu0.l_precountZ0Z_3\
        );

    \I__819\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9525\
        );

    \I__818\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9525\
        );

    \I__817\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9525\
        );

    \I__816\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9525\
        );

    \I__815\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9525\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__9525\,
            I => \uu0.l_precountZ0Z_1\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__9522\,
            I => \N__9516\
        );

    \I__812\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9507\
        );

    \I__811\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9507\
        );

    \I__810\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9507\
        );

    \I__809\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9507\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__9507\,
            I => \uu0.l_precountZ0Z_2\
        );

    \I__807\ : IoInMux
    port map (
            O => \N__9504\,
            I => \N__9501\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9498\
        );

    \I__805\ : IoSpan4Mux
    port map (
            O => \N__9498\,
            I => \N__9495\
        );

    \I__804\ : Odrv4
    port map (
            O => \N__9495\,
            I => clk_in_c
        );

    \INVuu2.bitmap_84C\ : INV
    port map (
            O => \INVuu2.bitmap_84C_net\,
            I => \N__26194\
        );

    \INVuu2.bitmap_212C\ : INV
    port map (
            O => \INVuu2.bitmap_212C_net\,
            I => \N__26200\
        );

    \INVuu2.w_addr_displaying_0C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_0C_net\,
            I => \N__26204\
        );

    \INVuu2.bitmap_87C\ : INV
    port map (
            O => \INVuu2.bitmap_87C_net\,
            I => \N__26186\
        );

    \INVuu2.bitmap_314C\ : INV
    port map (
            O => \INVuu2.bitmap_314C_net\,
            I => \N__26193\
        );

    \INVuu2.w_addr_user_5C\ : INV
    port map (
            O => \INVuu2.w_addr_user_5C_net\,
            I => \N__26203\
        );

    \INVuu2.bitmap_93C\ : INV
    port map (
            O => \INVuu2.bitmap_93C_net\,
            I => \N__26178\
        );

    \INVuu2.bitmap_215C\ : INV
    port map (
            O => \INVuu2.bitmap_215C_net\,
            I => \N__26185\
        );

    \INVuu2.w_addr_displaying_3C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_3C_net\,
            I => \N__26192\
        );

    \INVuu2.w_addr_displaying_nesr_5C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_nesr_5C_net\,
            I => \N__26199\
        );

    \INVuu2.bitmap_197C\ : INV
    port map (
            O => \INVuu2.bitmap_197C_net\,
            I => \N__26177\
        );

    \INVuu2.w_addr_displaying_1C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_1C_net\,
            I => \N__26184\
        );

    \INVuu2.bitmap_203C\ : INV
    port map (
            O => \INVuu2.bitmap_203C_net\,
            I => \N__26191\
        );

    \INVuu2.bitmap_111C\ : INV
    port map (
            O => \INVuu2.bitmap_111C_net\,
            I => \N__26152\
        );

    \INVuu2.bitmap_66C\ : INV
    port map (
            O => \INVuu2.bitmap_66C_net\,
            I => \N__26160\
        );

    \INVuu2.bitmap_296C\ : INV
    port map (
            O => \INVuu2.bitmap_296C_net\,
            I => \N__26169\
        );

    \INVuu2.w_addr_displaying_4C\ : INV
    port map (
            O => \INVuu2.w_addr_displaying_4C_net\,
            I => \N__26163\
        );

    \INVuu2.w_addr_user_nesr_8C\ : INV
    port map (
            O => \INVuu2.w_addr_user_nesr_8C_net\,
            I => \N__26176\
        );

    \INVuu2.w_addr_user_1C\ : INV
    port map (
            O => \INVuu2.w_addr_user_1C_net\,
            I => \N__26183\
        );

    \INVuu2.r_data_reg_0C\ : INV
    port map (
            O => \INVuu2.r_data_reg_0C_net\,
            I => \N__26202\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11862\,
            GLOBALBUFFEROUTPUT => clk_g
        );

    \bu_rx_data_rdy_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25611\,
            GLOBALBUFFEROUTPUT => bu_rx_data_rdy_0_g
        );

    \uu0.delay_line_RNILLLG7_0_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11544\,
            GLOBALBUFFEROUTPUT => \uu0.un11_l_count_i_g\
        );

    \buart.Z_rx.sample_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9825\,
            GLOBALBUFFEROUTPUT => \buart.Z_rx.sample_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \resetGen.rst_RNI4PQ1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__16693\,
            GLOBALBUFFEROUTPUT => rst_g
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \uu2.vram_rd_clk_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14667\,
            in2 => \_gnd_net_\,
            in3 => \N__11439\,
            lcout => \uu2.vram_rd_clkZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => 'H',
            sr => \N__25833\
        );

    \uu0.l_precount_0_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9622\,
            lcout => \uu0.l_precountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26205\,
            ce => 'H',
            sr => \N__25833\
        );

    \uu0.l_count_5_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10624\,
            in1 => \N__12257\,
            in2 => \_gnd_net_\,
            in3 => \N__12236\,
            lcout => \uu0.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__10442\,
            sr => \N__25830\
        );

    \uu0.l_count_8_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10488\,
            in2 => \_gnd_net_\,
            in3 => \N__10328\,
            lcout => \uu0.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26201\,
            ce => \N__10442\,
            sr => \N__25830\
        );

    \uu0.delay_line_0_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9537\,
            in1 => \N__9625\,
            in2 => \N__9558\,
            in3 => \N__9519\,
            lcout => \uu0.delay_lineZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26195\,
            ce => 'H',
            sr => \N__25827\
        );

    \uu0.l_precount_3_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__9521\,
            in1 => \N__9556\,
            in2 => \N__9630\,
            in3 => \N__9540\,
            lcout => \uu0.l_precountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26195\,
            ce => 'H',
            sr => \N__25827\
        );

    \uu0.l_precount_RNI85Q91_3_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__12253\,
            in2 => \N__9557\,
            in3 => \N__10377\,
            lcout => \uu0.un4_l_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_precount_1_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9624\,
            in2 => \_gnd_net_\,
            in3 => \N__9538\,
            lcout => \uu0.l_precountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26195\,
            ce => 'H',
            sr => \N__25827\
        );

    \uu0.l_precount_2_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__9539\,
            in1 => \N__9626\,
            in2 => \_gnd_net_\,
            in3 => \N__9520\,
            lcout => \uu0.l_precountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26195\,
            ce => 'H',
            sr => \N__25827\
        );

    \uu0.l_precount_RNI3Q7K1_2_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10317\,
            in1 => \N__10659\,
            in2 => \N__9522\,
            in3 => \N__10400\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIO2782_16_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9623\,
            in1 => \N__10242\,
            in2 => \N__9597\,
            in3 => \N__10773\,
            lcout => \uu0.un4_l_count_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10770\,
            in1 => \N__9571\,
            in2 => \N__10744\,
            in3 => \N__9586\,
            lcout => \uu0.un198_ci_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10354\,
            in1 => \N__10329\,
            in2 => \N__10566\,
            in3 => \N__10295\,
            lcout => \uu0.un154_ci_9\,
            ltout => \uu0.un154_ci_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10771\,
            in1 => \_gnd_net_\,
            in2 => \N__9594\,
            in3 => \N__9587\,
            lcout => OPEN,
            ltout => \uu0.un187_ci_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_15_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__9572\,
            in1 => \N__10496\,
            in2 => \N__9591\,
            in3 => \N__11595\,
            lcout => \uu0.l_countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26188\,
            ce => \N__10439\,
            sr => \N__25824\
        );

    \uu0.l_count_14_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__10494\,
            in2 => \N__10745\,
            in3 => \N__9588\,
            lcout => \uu0.l_countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26188\,
            ce => \N__10439\,
            sr => \N__25824\
        );

    \uu0.l_count_4_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__10623\,
            in1 => \N__12226\,
            in2 => \_gnd_net_\,
            in3 => \N__11596\,
            lcout => \uu0.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26188\,
            ce => \N__10439\,
            sr => \N__25824\
        );

    \uu0.l_count_10_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__10296\,
            in1 => \N__10495\,
            in2 => \N__10335\,
            in3 => \N__10355\,
            lcout => \uu0.l_countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26188\,
            ce => \N__10439\,
            sr => \N__25824\
        );

    \uu0.l_count_RNIGTCU_15_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9585\,
            in1 => \N__10353\,
            in2 => \N__9573\,
            in3 => \N__12225\,
            lcout => \uu0.un4_l_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9771\,
            in2 => \N__9648\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_2_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9678\,
            in2 => \_gnd_net_\,
            in3 => \N__9726\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_1\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            clk => \N__26180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_3_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11488\,
            in1 => \N__9668\,
            in2 => \_gnd_net_\,
            in3 => \N__9723\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_2\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            clk => \N__26180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_4_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9702\,
            in2 => \_gnd_net_\,
            in3 => \N__9720\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_3\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            clk => \N__26180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_5_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__9711\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \buart.Z_tx.Z_baudgen.un2_counter_cry_4\,
            carryout => \buart.Z_tx.Z_baudgen.un2_counter_cry_5\,
            clk => \N__26180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_6_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11487\,
            in2 => \N__9693\,
            in3 => \N__9714\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9710\,
            in1 => \N__9701\,
            in2 => \N__9692\,
            in3 => \N__9677\,
            lcout => \buart.Z_tx.Z_baudgen.ser_clk_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9643\,
            in1 => \N__9768\,
            in2 => \N__9669\,
            in3 => \N__9654\,
            lcout => \buart.Z_tx.ser_clk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_1_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9770\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.Z_baudgen.counter_0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9769\,
            lcout => \buart.Z_tx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26173\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m75_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10689\,
            in1 => \N__10868\,
            in2 => \N__9750\,
            in3 => \N__12608\,
            lcout => \N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m82_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__12610\,
            in1 => \N__10691\,
            in2 => \N__10880\,
            in3 => \N__9747\,
            lcout => OPEN,
            ltout => \resetGen_reset_count_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_2_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__9749\,
            in1 => \N__10909\,
            in2 => \N__9753\,
            in3 => \N__12611\,
            lcout => \resetGen_reset_count_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m78_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__12609\,
            in1 => \N__10690\,
            in2 => \N__10879\,
            in3 => \N__9748\,
            lcout => \N_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.rst_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10910\,
            lcout => rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_3_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__16250\,
            in1 => \N__16181\,
            in2 => \N__9807\,
            in3 => \N__14951\,
            lcout => \buart__rx_bitcount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26156\,
            ce => \N__16081\,
            sr => \N__25817\
        );

    \buart.Z_rx.bitcount_cry_c_0_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9850\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => \buart.Z_rx.bitcount_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9920\,
            in2 => \_gnd_net_\,
            in3 => \N__9732\,
            lcout => \buart.Z_rx.bitcount_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_0\,
            carryout => \buart.Z_rx.bitcount_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16131\,
            in2 => \_gnd_net_\,
            in3 => \N__9729\,
            lcout => \buart.Z_rx.bitcount_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_1\,
            carryout => \buart.Z_rx.bitcount_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14950\,
            in2 => \_gnd_net_\,
            in3 => \N__9798\,
            lcout => \buart.Z_rx.bitcount_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.bitcount_cry_2\,
            carryout => \buart.Z_rx.bitcount_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_4_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__16249\,
            in1 => \N__16174\,
            in2 => \N__9895\,
            in3 => \N__9795\,
            lcout => \buart__rx_bitcount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26150\,
            ce => \N__16085\,
            sr => \N__25818\
        );

    \Lab_UT.dispString.m103_ns_1_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000111111"
        )
    port map (
            in0 => \N__9998\,
            in1 => \N__14958\,
            in2 => \N__9936\,
            in3 => \N__14882\,
            lcout => OPEN,
            ltout => \Lab_UT_dispString_m103_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_sbtinv_4_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101111001010"
        )
    port map (
            in0 => \N__9780\,
            in1 => \N__9999\,
            in2 => \N__9792\,
            in3 => \N__25924\,
            lcout => \buart.Z_rx.bitcounte_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_0_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__16238\,
            in1 => \N__16173\,
            in2 => \N__16959\,
            in3 => \N__9854\,
            lcout => \buart__rx_bitcount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26144\,
            ce => \N__16077\,
            sr => \N__25819\
        );

    \Lab_UT.dispString.N_27_0_i_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14883\,
            in1 => \N__9935\,
            in2 => \_gnd_net_\,
            in3 => \N__14959\,
            lcout => \buart__rx_N_27_0_i\,
            ltout => \buart__rx_N_27_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_1_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101001101011100"
        )
    port map (
            in0 => \N__16239\,
            in1 => \N__9789\,
            in2 => \N__9783\,
            in3 => \N__9921\,
            lcout => \buart__rx_bitcount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26144\,
            ce => \N__16077\,
            sr => \N__25819\
        );

    \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16128\,
            in1 => \N__9917\,
            in2 => \N__9896\,
            in3 => \N__9848\,
            lcout => \buart__rx_valid_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m103_e_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11740\,
            in2 => \_gnd_net_\,
            in3 => \N__10846\,
            lcout => \N_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_0_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9942\,
            lcout => \buart__rx_hh_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26135\,
            ce => 'H',
            sr => \N__25821\
        );

    \Lab_UT.dispString.m8_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16129\,
            in1 => \N__9919\,
            in2 => \N__9897\,
            in3 => \N__9849\,
            lcout => \Lab_UT.dispString.N_115_mux\,
            ltout => \Lab_UT.dispString.N_115_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m11_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14960\,
            in1 => \N__10847\,
            in2 => \N__9924\,
            in3 => \N__11741\,
            lcout => \buart__rx_startbit\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m97_e_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9918\,
            in1 => \N__9891\,
            in2 => \_gnd_net_\,
            in3 => \N__14957\,
            lcout => \Lab_UT.dispString.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_2_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__10073\,
            in1 => \N__16241\,
            in2 => \N__10059\,
            in3 => \N__9996\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI2GE3_1_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10046\,
            in1 => \N__10072\,
            in2 => \N__10031\,
            in3 => \N__10108\,
            lcout => OPEN,
            ltout => \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_RNI3O55_5_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9965\,
            in2 => \N__9867\,
            in3 => \N__10089\,
            lcout => \buart__rx_ser_clk\,
            ltout => \buart__rx_ser_clk_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m98_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000000000000"
        )
    port map (
            in0 => \N__9864\,
            in1 => \N__16130\,
            in2 => \N__9858\,
            in3 => \N__9855\,
            lcout => \buart__rx_sample\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_4_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__10008\,
            in1 => \N__16242\,
            in2 => \N__10032\,
            in3 => \N__9997\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_1_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__10091\,
            in1 => \_gnd_net_\,
            in2 => \N__16253\,
            in3 => \N__10109\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_0_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16240\,
            in2 => \_gnd_net_\,
            in3 => \N__10090\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26131\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10110\,
            in2 => \N__10095\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10074\,
            in2 => \_gnd_net_\,
            in3 => \N__10050\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_1\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_3_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16252\,
            in1 => \N__10047\,
            in2 => \_gnd_net_\,
            in3 => \N__10035\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_2\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            clk => \N__26128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10027\,
            in2 => \_gnd_net_\,
            in3 => \N__10002\,
            lcout => \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \buart.Z_rx.Z_baudgen.un5_counter_cry_3\,
            carryout => \buart.Z_rx.Z_baudgen.un5_counter_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.Z_baudgen.counter_5_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__9995\,
            in1 => \N__16251\,
            in2 => \N__9969\,
            in3 => \N__9972\,
            lcout => \buart.Z_rx.Z_baudgen.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9954\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9948\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_2_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_3_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10170\,
            lcout => vbuf_tx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_4_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10164\,
            lcout => vbuf_tx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_5_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10158\,
            lcout => vbuf_tx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_6_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10152\,
            lcout => vbuf_tx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \uu2.r_data_reg_7_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vbuf_tx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.r_data_reg_0C_net\,
            ce => \N__16011\,
            sr => \_gnd_net_\
        );

    \buart.Z_tx.shifter_1_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12122\,
            in1 => \N__10221\,
            in2 => \_gnd_net_\,
            in3 => \N__10140\,
            lcout => \buart.Z_tx.shifterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.shifter_0_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10134\,
            in2 => \_gnd_net_\,
            in3 => \N__12120\,
            lcout => \buart.Z_tx.shifterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.uart_tx_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10128\,
            lcout => o_serial_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.shifter_2_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10209\,
            in1 => \N__12123\,
            in2 => \_gnd_net_\,
            in3 => \N__10227\,
            lcout => \buart.Z_tx.shifterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.shifter_3_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12124\,
            in1 => \N__10197\,
            in2 => \_gnd_net_\,
            in3 => \N__10215\,
            lcout => \buart.Z_tx.shifterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.shifter_4_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10185\,
            in1 => \N__12125\,
            in2 => \_gnd_net_\,
            in3 => \N__10203\,
            lcout => \buart.Z_tx.shifterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \buart.Z_tx.shifter_5_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12126\,
            in1 => \N__10413\,
            in2 => \_gnd_net_\,
            in3 => \N__10191\,
            lcout => \buart.Z_tx.shifterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26196\,
            ce => \N__10803\,
            sr => \N__25834\
        );

    \uu0.l_count_6_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__12372\,
            in1 => \N__12346\,
            in2 => \N__10625\,
            in3 => \N__11601\,
            lcout => \uu0.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26189\,
            ce => \N__10443\,
            sr => \N__25832\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10402\,
            lcout => \uu0.un44_ci\,
            ltout => \uu0.un44_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_2_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10179\,
            in3 => \N__10661\,
            lcout => \uu0.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26189\,
            ce => \N__10443\,
            sr => \N__25832\
        );

    \uu0.l_count_1_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__10382\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10404\,
            lcout => \uu0.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26189\,
            ce => \N__10443\,
            sr => \N__25832\
        );

    \uu0.l_count_0_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10403\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11599\,
            lcout => \uu0.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26189\,
            ce => \N__10443\,
            sr => \N__25832\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10660\,
            in1 => \N__10401\,
            in2 => \N__10383\,
            in3 => \N__10641\,
            lcout => \uu0.un66_ci\,
            ltout => \uu0.un66_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12371\,
            in1 => \N__12345\,
            in2 => \N__10362\,
            in3 => \N__10596\,
            lcout => \uu0.un110_ci\,
            ltout => \uu0.un110_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_12_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__11600\,
            in1 => \N__10743\,
            in2 => \N__10359\,
            in3 => \N__10714\,
            lcout => \uu0.l_countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26189\,
            ce => \N__10443\,
            sr => \N__25832\
        );

    \uu0.l_count_RNIRLTJ1_17_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__10594\,
            in2 => \N__10275\,
            in3 => \N__10639\,
            lcout => \uu0.un4_l_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10333\,
            in1 => \N__10356\,
            in2 => \_gnd_net_\,
            in3 => \N__10293\,
            lcout => \uu0.un143_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_9_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__10487\,
            in2 => \_gnd_net_\,
            in3 => \N__10334\,
            lcout => \uu0.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26181\,
            ce => \N__10441\,
            sr => \N__25828\
        );

    \uu0.l_count_17_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__10245\,
            in1 => \N__10259\,
            in2 => \N__10498\,
            in3 => \N__10274\,
            lcout => \uu0.l_countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26181\,
            ce => \N__10441\,
            sr => \N__25828\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10273\,
            in1 => \N__10480\,
            in2 => \N__10260\,
            in3 => \N__10243\,
            lcout => \uu0.un220_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_16_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__10244\,
            in1 => \N__10258\,
            in2 => \N__10497\,
            in3 => \N__11585\,
            lcout => \uu0.l_countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26181\,
            ce => \N__10441\,
            sr => \N__25828\
        );

    \uu0.l_count_3_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__11587\,
            in1 => \N__10674\,
            in2 => \N__10668\,
            in3 => \N__10640\,
            lcout => \uu0.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26181\,
            ce => \N__10441\,
            sr => \N__25828\
        );

    \uu0.l_count_7_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__10595\,
            in1 => \N__12324\,
            in2 => \N__10626\,
            in3 => \N__11586\,
            lcout => \uu0.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26181\,
            ce => \N__10441\,
            sr => \N__25828\
        );

    \uu0.l_count_18_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__11584\,
            in1 => \_gnd_net_\,
            in2 => \N__10548\,
            in3 => \N__10581\,
            lcout => \uu0.l_countZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26174\,
            ce => \N__10440\,
            sr => \N__25825\
        );

    \uu0.l_count_11_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__10499\,
            in1 => \N__10562\,
            in2 => \N__10575\,
            in3 => \N__11583\,
            lcout => \uu0.l_countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26174\,
            ce => \N__10440\,
            sr => \N__25825\
        );

    \uu0.l_count_RNIOIDD2_18_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10561\,
            in1 => \N__12350\,
            in2 => \N__10547\,
            in3 => \N__10533\,
            lcout => OPEN,
            ltout => \uu0.un4_l_count_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNI8ORT6_15_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10527\,
            in1 => \N__10518\,
            in2 => \N__10512\,
            in3 => \N__10509\,
            lcout => \uu0.un4_l_count_0\,
            ltout => \uu0.un4_l_count_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_13_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__10698\,
            in1 => \N__10500\,
            in2 => \N__10446\,
            in3 => \N__10785\,
            lcout => \uu0.l_countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26174\,
            ce => \N__10440\,
            sr => \N__25825\
        );

    \buart.Z_tx.shifter_6_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12117\,
            in1 => \N__10824\,
            in2 => \_gnd_net_\,
            in3 => \N__10422\,
            lcout => \buart.Z_tx.shifterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26166\,
            ce => \N__10796\,
            sr => \N__25823\
        );

    \buart.Z_tx.shifter_7_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10833\,
            in1 => \N__10809\,
            in2 => \_gnd_net_\,
            in3 => \N__12118\,
            lcout => \buart.Z_tx.shifterZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26166\,
            ce => \N__10796\,
            sr => \N__25823\
        );

    \buart.Z_tx.shifter_8_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12116\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10818\,
            lcout => \buart.Z_tx.shifterZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26166\,
            ce => \N__10796\,
            sr => \N__25823\
        );

    \buart.Z_tx.bitcount_RNI22V22_2_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12115\,
            in2 => \_gnd_net_\,
            in3 => \N__11646\,
            lcout => \buart.Z_tx.un1_uart_wr_i_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25876\,
            in2 => \_gnd_net_\,
            in3 => \N__16635\,
            lcout => \Lab_UT.didp.regrce2.LdAStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16665\,
            lcout => \Lab_UT.didp.regrce4.LdAMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.l_count_RNIFAQ9_13_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10784\,
            lcout => \uu0.un4_l_count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10749\,
            in2 => \_gnd_net_\,
            in3 => \N__10716\,
            lcout => \uu0.un165_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010100010000"
        )
    port map (
            in0 => \N__12614\,
            in1 => \N__10905\,
            in2 => \N__10881\,
            in3 => \N__10692\,
            lcout => \resetGen_reset_count_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m72_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10903\,
            in2 => \_gnd_net_\,
            in3 => \N__12612\,
            lcout => OPEN,
            ltout => \m72_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_3_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110110101000"
        )
    port map (
            in0 => \N__10919\,
            in1 => \N__10938\,
            in2 => \N__10932\,
            in3 => \N__10928\,
            lcout => \resetGen.reset_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_4_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__10929\,
            in1 => \N__10920\,
            in2 => \N__10911\,
            in3 => \N__12615\,
            lcout => \resetGen_reset_count_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \resetGen.reset_count_0_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__10904\,
            in1 => \N__10875\,
            in2 => \_gnd_net_\,
            in3 => \N__12613\,
            lcout => \resetGen_reset_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26157\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.hh_1_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10851\,
            lcout => \buart__rx_hh_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26145\,
            ce => 'H',
            sr => \N__25820\
        );

    \buart.Z_rx.shifter_2_rep2_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26389\,
            lcout => bu_rx_data_2_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_3_rep1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18875\,
            lcout => bu_rx_data_3_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_4_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19047\,
            lcout => bu_rx_data_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_3_rep2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18876\,
            lcout => bu_rx_data_3_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_5_rep1_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19212\,
            lcout => bu_rx_data_5_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_7_rep1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11736\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_7_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11735\,
            lcout => bu_rx_data_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \buart.Z_rx.shifter_1_rep2_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26651\,
            lcout => bu_rx_data_1_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26136\,
            ce => \N__14244\,
            sr => \N__25822\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIEGPT_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__18586\,
            in1 => \N__18339\,
            in2 => \N__20503\,
            in3 => \N__19729\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_69_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNIDS133_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010100000101"
        )
    port map (
            in0 => \N__18340\,
            in1 => \N__10959\,
            in2 => \N__10962\,
            in3 => \N__14370\,
            lcout => \Lab_UT.dictrl.N_61_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_0_1_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13927\,
            in1 => \N__13839\,
            in2 => \N__18724\,
            in3 => \N__17117\,
            lcout => \Lab_UT.dictrl.g1_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_10_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__13838\,
            in1 => \N__20489\,
            in2 => \N__18725\,
            in3 => \N__13926\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g1_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_9_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19191\,
            in2 => \N__10953\,
            in3 => \N__19036\,
            lcout => \Lab_UT.dictrl.g1_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNII0HP5_2_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011000"
        )
    port map (
            in0 => \N__22813\,
            in1 => \N__10950\,
            in2 => \N__11061\,
            in3 => \N__10944\,
            lcout => \Lab_UT.dictrl.N_62_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_5_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__24317\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22814\,
            lcout => \Lab_UT.dictrl.g2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_3_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001011"
        )
    port map (
            in0 => \N__22816\,
            in1 => \N__24318\,
            in2 => \N__12543\,
            in3 => \N__11886\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1792_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100101100000"
        )
    port map (
            in0 => \N__24319\,
            in1 => \N__22817\,
            in2 => \N__10998\,
            in3 => \N__10995\,
            lcout => \Lab_UT.dictrl.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIE5JQ_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22812\,
            in2 => \_gnd_net_\,
            in3 => \N__24316\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIE5JQZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_2_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__10971\,
            in1 => \N__22815\,
            in2 => \N__10980\,
            in3 => \N__11760\,
            lcout => \Lab_UT.dictrl.N_1451_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__26616\,
            in1 => \N__24062\,
            in2 => \N__19737\,
            in3 => \N__21710\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_a5_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10986\,
            in2 => \N__10989\,
            in3 => \N__14373\,
            lcout => \Lab_UT.dictrl.N_10_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__26359\,
            in1 => \N__18854\,
            in2 => \N__25439\,
            in3 => \N__19209\,
            lcout => \Lab_UT.dictrl.g0_i_a5_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_8_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__21709\,
            in1 => \N__26358\,
            in2 => \N__18892\,
            in3 => \N__26615\,
            lcout => \Lab_UT.dictrl.g0_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_9_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000010"
        )
    port map (
            in0 => \N__14372\,
            in1 => \N__19208\,
            in2 => \N__25440\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.g0_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_0_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25408\,
            lcout => bu_rx_data_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26124\,
            ce => \N__14242\,
            sr => \N__25831\
        );

    \buart.Z_rx.shifter_1_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26617\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26124\,
            ce => \N__14242\,
            sr => \N__25831\
        );

    \buart.Z_rx.shifter_2_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26360\,
            lcout => bu_rx_data_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26124\,
            ce => \N__14242\,
            sr => \N__25831\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNI1TO01_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__18853\,
            in1 => \N__18234\,
            in2 => \N__18152\,
            in3 => \N__19730\,
            lcout => \Lab_UT.dictrl.g1_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_rep2_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18129\,
            lcout => bu_rx_data_6_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26119\,
            ce => \N__14239\,
            sr => \N__25837\
        );

    \uu2.r_addr_esr_7_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11215\,
            in1 => \N__11049\,
            in2 => \N__11024\,
            in3 => \N__11977\,
            lcout => \uu2.r_addrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26190\,
            ce => \N__11118\,
            sr => \N__25812\
        );

    \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12005\,
            lcout => \uu2.vbuf_raddr.un426_ci_3\,
            ltout => \uu2.vbuf_raddr.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_8_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__11036\,
            in1 => \N__11004\,
            in2 => \N__11043\,
            in3 => \N__11976\,
            lcout => \uu2.r_addrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26190\,
            ce => \N__11118\,
            sr => \N__25812\
        );

    \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11017\,
            in2 => \_gnd_net_\,
            in3 => \N__11214\,
            lcout => \uu2.vbuf_raddr.un448_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11166\,
            in1 => \N__11138\,
            in2 => \N__11197\,
            in3 => \N__11098\,
            lcout => \uu2.un404_ci_0\,
            ltout => \uu2.un404_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_esr_6_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__11929\,
            in1 => \N__11216\,
            in2 => \N__11223\,
            in3 => \N__12006\,
            lcout => \uu2.r_addrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26190\,
            ce => \N__11118\,
            sr => \N__25812\
        );

    \uu2.r_addr_esr_3_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11167\,
            in1 => \N__11139\,
            in2 => \N__11198\,
            in3 => \N__11099\,
            lcout => \uu2.r_addrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26190\,
            ce => \N__11118\,
            sr => \N__25812\
        );

    \uu2.r_addr_2_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__11141\,
            in1 => \N__11104\,
            in2 => \N__11174\,
            in3 => \N__11957\,
            lcout => \uu2.r_addrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.r_addr_1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__11955\,
            in1 => \_gnd_net_\,
            in2 => \N__11108\,
            in3 => \N__11140\,
            lcout => \uu2.r_addrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.trig_rd_det_RNINBDQ_1_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11954\,
            in2 => \_gnd_net_\,
            in3 => \N__25880\,
            lcout => \uu2.trig_rd_is_det_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.trig_rd_det_RNIJIIO_1_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11076\,
            in2 => \_gnd_net_\,
            in3 => \N__11069\,
            lcout => \uu2.trig_rd_is_det\,
            ltout => \uu2.trig_rd_is_det_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_addr_0_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11112\,
            in3 => \N__11100\,
            lcout => \uu2.r_addrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.trig_rd_det_1_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11070\,
            lcout => \uu2.trig_rd_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.trig_rd_det_0_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14683\,
            in2 => \_gnd_net_\,
            in3 => \N__12137\,
            lcout => \uu2.trig_rd_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.r_addr_4_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11956\,
            in1 => \N__12007\,
            in2 => \_gnd_net_\,
            in3 => \N__11978\,
            lcout => \uu2.r_addrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26182\,
            ce => 'H',
            sr => \N__25805\
        );

    \uu2.l_count_RNIFGGK1_3_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11314\,
            in1 => \N__11458\,
            in2 => \N__11265\,
            in3 => \N__11293\,
            lcout => \uu2.un1_l_count_1_3\,
            ltout => \uu2.un1_l_count_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_RNI9S834_1_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11244\,
            in1 => \N__12193\,
            in2 => \N__11277\,
            in3 => \N__11373\,
            lcout => \uu2.un1_l_count_2_0\,
            ltout => \uu2.un1_l_count_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_3_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__12207\,
            in1 => \N__11246\,
            in2 => \N__11274\,
            in3 => \N__11264\,
            lcout => \uu2.l_countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26175\,
            ce => 'H',
            sr => \N__25839\
        );

    \uu2.l_count_2_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11245\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12206\,
            lcout => \uu2.l_countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26175\,
            ce => 'H',
            sr => \N__25839\
        );

    \uu2.l_count_RNI9S834_0_1_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12192\,
            in1 => \N__11271\,
            in2 => \N__11469\,
            in3 => \N__11243\,
            lcout => \uu2.un1_l_count_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11263\,
            in1 => \N__12191\,
            in2 => \N__11247\,
            in3 => \N__12171\,
            lcout => \uu2.un306_ci\,
            ltout => \uu2.un306_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_4_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001001000010010"
        )
    port map (
            in0 => \N__11411\,
            in1 => \N__11434\,
            in2 => \N__11226\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26175\,
            ce => 'H',
            sr => \N__25839\
        );

    \uu2.l_count_5_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11410\,
            in2 => \N__11367\,
            in3 => \N__11460\,
            lcout => \uu2.l_countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26175\,
            ce => 'H',
            sr => \N__25839\
        );

    \uu2.l_count_RNIBCGK1_0_9_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11330\,
            in1 => \N__11408\,
            in2 => \N__11388\,
            in3 => \N__12169\,
            lcout => \uu2.un1_l_count_1_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_6_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__11345\,
            in1 => \N__11333\,
            in2 => \_gnd_net_\,
            in3 => \N__11362\,
            lcout => \uu2.l_countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26167\,
            ce => 'H',
            sr => \N__25836\
        );

    \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11459\,
            in2 => \_gnd_net_\,
            in3 => \N__11409\,
            lcout => \uu2.vbuf_count.un328_ci_3\,
            ltout => \uu2.vbuf_count.un328_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11315\,
            in1 => \N__11332\,
            in2 => \N__11442\,
            in3 => \N__11361\,
            lcout => \uu2.un350_ci\,
            ltout => \uu2.un350_ci_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_9_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__11387\,
            in1 => \N__11435\,
            in2 => \N__11415\,
            in3 => \N__11295\,
            lcout => \uu2.l_countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26167\,
            ce => 'H',
            sr => \N__25836\
        );

    \uu2.l_count_RNIBCGK1_9_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__12170\,
            in1 => \N__11331\,
            in2 => \N__11412\,
            in3 => \N__11386\,
            lcout => \uu2.un1_l_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_7_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__11363\,
            in1 => \N__11346\,
            in2 => \N__11337\,
            in3 => \N__11316\,
            lcout => \uu2.l_countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26167\,
            ce => 'H',
            sr => \N__25836\
        );

    \uu2.l_count_8_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11294\,
            in2 => \_gnd_net_\,
            in3 => \N__11301\,
            lcout => \uu2.l_countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26167\,
            ce => 'H',
            sr => \N__25836\
        );

    \Lab_UT.dispString.cnt_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__13680\,
            in1 => \N__13411\,
            in2 => \N__22070\,
            in3 => \N__13541\,
            lcout => \Lab_UT.dispString.cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26158\,
            ce => 'H',
            sr => \N__25800\
        );

    \Lab_UT.dispString.cnt_1_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13540\,
            lcout => \Lab_UT.dispString.cntZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26158\,
            ce => 'H',
            sr => \N__25800\
        );

    \Lab_UT.dispString.cnt_2_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__12282\,
            in1 => \_gnd_net_\,
            in2 => \N__13699\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dispString.cntZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26158\,
            ce => 'H',
            sr => \N__25800\
        );

    \uu0.sec_clk_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__11598\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14722\,
            lcout => \o_One_Sec_Pulse\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26158\,
            ce => 'H',
            sr => \N__25800\
        );

    \uu0.delay_line_RNILLLG7_1_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__11514\,
            in1 => \N__11528\,
            in2 => \_gnd_net_\,
            in3 => \N__11597\,
            lcout => \uu0.un11_l_count_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.delay_line_1_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__11529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uu0.delay_lineZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26158\,
            ce => 'H',
            sr => \N__25800\
        );

    \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11504\,
            in2 => \_gnd_net_\,
            in3 => \N__11615\,
            lcout => \buart.Z_tx.uart_busy_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_3_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__11617\,
            in1 => \N__11681\,
            in2 => \N__11664\,
            in3 => \N__11642\,
            lcout => OPEN,
            ltout => \buart.Z_tx.un1_bitcount_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_3_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101110111110"
        )
    port map (
            in0 => \N__12098\,
            in1 => \N__11645\,
            in2 => \N__11508\,
            in3 => \N__11505\,
            lcout => \buart.Z_tx.bitcountZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26151\,
            ce => 'H',
            sr => \N__25829\
        );

    \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100000000"
        )
    port map (
            in0 => \N__11658\,
            in1 => \N__11496\,
            in2 => \N__11682\,
            in3 => \N__11490\,
            lcout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2\,
            ltout => \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_RNO_0_2_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__11680\,
            in1 => \N__11659\,
            in2 => \N__11688\,
            in3 => \N__11616\,
            lcout => OPEN,
            ltout => \buart.Z_tx.bitcount_RNO_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_tx.bitcount_2_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11685\,
            in3 => \N__12093\,
            lcout => \buart.Z_tx.bitcountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26151\,
            ce => 'H',
            sr => \N__25829\
        );

    \buart.Z_tx.bitcount_1_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110110"
        )
    port map (
            in0 => \N__11643\,
            in1 => \N__11663\,
            in2 => \N__12119\,
            in3 => \N__11619\,
            lcout => \buart.Z_tx.bitcountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26151\,
            ce => 'H',
            sr => \N__25829\
        );

    \buart.Z_tx.bitcount_0_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__11618\,
            in1 => \N__12094\,
            in2 => \_gnd_net_\,
            in3 => \N__11644\,
            lcout => \buart.Z_tx.bitcountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26151\,
            ce => 'H',
            sr => \N__25829\
        );

    \buart.Z_rx.shifter_2_rep2_RNICDH61_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__18891\,
            in1 => \N__21779\,
            in2 => \N__18141\,
            in3 => \N__13883\,
            lcout => \buart.Z_rx.G_17_i_a5_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13413\,
            in2 => \_gnd_net_\,
            in3 => \N__13543\,
            lcout => \Lab_UT.dispString.N_30_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m4_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14953\,
            in2 => \_gnd_net_\,
            in3 => \N__14894\,
            lcout => bu_rx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m71_0_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18910\,
            in2 => \_gnd_net_\,
            in3 => \N__25503\,
            lcout => \Lab_UT.dictrl.m71Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_12_a6_3_7_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19017\,
            in1 => \N__21749\,
            in2 => \N__19190\,
            in3 => \N__26348\,
            lcout => \Lab_UT.dictrl.g0_12_a6_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_RNIH0Q52_5_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__19157\,
            in1 => \N__13329\,
            in2 => \N__13790\,
            in3 => \N__19018\,
            lcout => \N_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_25_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__26349\,
            in1 => \N__19019\,
            in2 => \N__19192\,
            in3 => \N__11700\,
            lcout => \Lab_UT.dictrl.N_97_mux_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIF4VT_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__19423\,
            in1 => \N__20360\,
            in2 => \N__18585\,
            in3 => \N__16592\,
            lcout => \Lab_UT.dictrl.g0_12_o6_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIMFOD2_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14832\,
            in1 => \N__17096\,
            in2 => \_gnd_net_\,
            in3 => \N__19917\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_13_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNIJT0P3_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__11709\,
            in1 => \N__19710\,
            in2 => \N__11703\,
            in3 => \N__16829\,
            lcout => \Lab_UT.dictrl.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIOEMF_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__16593\,
            in1 => \N__14833\,
            in2 => \N__12684\,
            in3 => \N__12725\,
            lcout => \Lab_UT.dictrl.N_17_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m34_4_2_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__17094\,
            in1 => \N__12677\,
            in2 => \_gnd_net_\,
            in3 => \N__14045\,
            lcout => \Lab_UT.dictrl.m34_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m59_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12721\,
            in2 => \_gnd_net_\,
            in3 => \N__14046\,
            lcout => \Lab_UT_dictrl_m59_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_10_3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__12678\,
            in1 => \N__17095\,
            in2 => \N__12726\,
            in3 => \N__19424\,
            lcout => \Lab_UT.dictrl.g0_10Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIOIIC1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13963\,
            in1 => \N__11694\,
            in2 => \N__20488\,
            in3 => \N__15636\,
            lcout => \Lab_UT.dictrl.m34_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_12_o3_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__18729\,
            in1 => \N__13877\,
            in2 => \_gnd_net_\,
            in3 => \N__13956\,
            lcout => \Lab_UT.dictrl.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_17_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13957\,
            in1 => \N__18730\,
            in2 => \N__13887\,
            in3 => \N__20267\,
            lcout => \Lab_UT.dictrl.g1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_13_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__20268\,
            in1 => \N__13881\,
            in2 => \N__18752\,
            in3 => \N__13959\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_0_o7_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_6_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__19149\,
            in1 => \N__21770\,
            in2 => \N__11712\,
            in3 => \N__14371\,
            lcout => \Lab_UT.dictrl.N_15_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_8_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13882\,
            in1 => \N__13958\,
            in2 => \N__18751\,
            in3 => \N__24011\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_a7_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep2_RNIDJQN_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__18994\,
            in1 => \N__18750\,
            in2 => \N__19150\,
            in3 => \N__13964\,
            lcout => \buart.Z_rx.G_17_i_a5_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_5_1_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19115\,
            in2 => \_gnd_net_\,
            in3 => \N__18995\,
            lcout => \Lab_UT.dictrl.g0_i_a4_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_5_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19116\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_6_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18137\,
            lcout => bu_rx_data_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_fast_5_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_fast_4_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18998\,
            lcout => bu_rx_data_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_4_rep1_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18996\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_4_rep2_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18997\,
            lcout => bu_rx_data_4_rep2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26122\,
            ce => \N__14241\,
            sr => \N__25835\
        );

    \buart.Z_rx.shifter_0_rep1_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_0_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_fast_0_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25456\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_1_rep1_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26649\,
            lcout => bu_rx_data_1_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_fast_1_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26650\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_fast_7_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => bu_rx_data_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_2_rep1_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26330\,
            lcout => bu_rx_data_2_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_3_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18933\,
            lcout => bu_rx_data_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \buart.Z_rx.shifter_fast_2_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26331\,
            lcout => bu_rx_data_fast_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26120\,
            ce => \N__14240\,
            sr => \N__25838\
        );

    \Lab_UT.dictrl.g0_9_3_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__12783\,
            in1 => \N__12829\,
            in2 => \N__12762\,
            in3 => \N__12996\,
            lcout => \Lab_UT.dictrl.g0_9Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_i_m2_1_o6_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12754\,
            in2 => \_gnd_net_\,
            in3 => \N__12781\,
            lcout => \Lab_UT.dictrl.N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m23_a0_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__12782\,
            in1 => \_gnd_net_\,
            in2 => \N__12761\,
            in3 => \N__12995\,
            lcout => \Lab_UT.dictrl.m23_aZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m40_1_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__12994\,
            in1 => \N__12753\,
            in2 => \N__14108\,
            in3 => \N__12780\,
            lcout => \Lab_UT.dictrl.m40Z0Z_1\,
            ltout => \Lab_UT.dictrl.m40Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__18931\,
            in1 => \N__22819\,
            in2 => \N__11799\,
            in3 => \N__20577\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__11796\,
            in1 => \N__17238\,
            in2 => \N__11784\,
            in3 => \N__19473\,
            lcout => \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_3_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18932\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => bu_rx_data_fast_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26118\,
            ce => \N__14238\,
            sr => \N__25840\
        );

    \Lab_UT.dictrl.g0_8_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20296\,
            in1 => \N__18595\,
            in2 => \N__11781\,
            in3 => \N__20406\,
            lcout => \Lab_UT.dictrl.N_97_mux_0\,
            ltout => \Lab_UT.dictrl.N_97_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_10_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111101110"
        )
    port map (
            in0 => \N__11901\,
            in1 => \N__11772\,
            in2 => \N__11763\,
            in3 => \N__19735\,
            lcout => \Lab_UT.dictrl.N_2435_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_18_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__20493\,
            in1 => \N__20402\,
            in2 => \N__20045\,
            in3 => \N__19446\,
            lcout => \Lab_UT.dictrl.g1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_20_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19447\,
            in1 => \N__18594\,
            in2 => \N__20409\,
            in3 => \N__20295\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_16_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_12_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__12840\,
            in1 => \N__11895\,
            in2 => \N__11889\,
            in3 => \N__20576\,
            lcout => \Lab_UT.dictrl.N_2446_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__23606\,
            in1 => \N__12041\,
            in2 => \N__23692\,
            in3 => \N__23381\,
            lcout => \uu2.mem0.w_addr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_wr_en_0_i_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011101"
        )
    port map (
            in0 => \N__11855\,
            in1 => \N__23668\,
            in2 => \_gnd_net_\,
            in3 => \N__23603\,
            lcout => \uu2.vram_wr_en_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_0_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__23604\,
            in1 => \N__17551\,
            in2 => \N__23691\,
            in3 => \N__23490\,
            lcout => \uu2.mem0.w_addr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_1_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20959\,
            in1 => \_gnd_net_\,
            in2 => \N__12048\,
            in3 => \N__17555\,
            lcout => \uu2.w_addr_userZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__20843\
        );

    \uu2.w_addr_user_2_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__17556\,
            in1 => \N__12047\,
            in2 => \N__17522\,
            in3 => \N__20960\,
            lcout => \uu2.w_addr_userZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__20843\
        );

    \uu2.mem0.ram512X8_inst_RNO_1_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__17513\,
            in1 => \N__23669\,
            in2 => \N__17376\,
            in3 => \N__23605\,
            lcout => \uu2.mem0.w_addr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12043\,
            in2 => \_gnd_net_\,
            in3 => \N__20958\,
            lcout => \uu2.w_addr_userZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_1C_net\,
            ce => 'H',
            sr => \N__20843\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_5_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12042\,
            in1 => \N__17514\,
            in2 => \N__17559\,
            in3 => \N__13089\,
            lcout => \uu2.un404_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI1VU6_3_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__21050\,
            in1 => \N__13077\,
            in2 => \N__14420\,
            in3 => \N__12039\,
            lcout => \uu2.un3_w_addr_user_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14415\,
            in2 => \_gnd_net_\,
            in3 => \N__20882\,
            lcout => OPEN,
            ltout => \uu2.vbuf_w_addr_user.un448_ci_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_8_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__23533\,
            in1 => \N__20921\,
            in2 => \N__12051\,
            in3 => \N__20894\,
            lcout => \uu2.w_addr_userZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12147\,
            sr => \N__20842\
        );

    \uu2.w_addr_user_nesr_3_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12040\,
            in1 => \N__17518\,
            in2 => \N__13087\,
            in3 => \N__17557\,
            lcout => \uu2.w_addr_userZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12147\,
            sr => \N__20842\
        );

    \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21014\,
            lcout => \uu2.un426_ci_3\,
            ltout => \uu2.un426_ci_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_7_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__20920\,
            in1 => \N__14416\,
            in2 => \N__12018\,
            in3 => \N__20883\,
            lcout => \uu2.w_addr_userZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_nesr_8C_net\,
            ce => \N__12147\,
            sr => \N__20842\
        );

    \uu2.r_addr_5_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__12014\,
            in1 => \N__11982\,
            in2 => \N__11930\,
            in3 => \N__11958\,
            lcout => \uu2.r_addrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26168\,
            ce => 'H',
            sr => \N__25806\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12261\,
            in2 => \_gnd_net_\,
            in3 => \N__12237\,
            lcout => \uu0.un88_ci_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12194\,
            in2 => \_gnd_net_\,
            in3 => \N__12172\,
            lcout => \uu2.un284_ci\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.l_count_1_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__12174\,
            in1 => \_gnd_net_\,
            in2 => \N__12198\,
            in3 => \_gnd_net_\,
            lcout => \uu2.l_countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26168\,
            ce => 'H',
            sr => \N__25806\
        );

    \uu2.l_count_0_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12173\,
            lcout => \uu2.l_countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26168\,
            ce => 'H',
            sr => \N__25806\
        );

    \uu2.w_addr_displaying_nesr_RNO_0_5_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16726\,
            in2 => \_gnd_net_\,
            in3 => \N__25019\,
            lcout => \uu2.un21_w_addr_displaying_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNID65PE_2_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20947\,
            in2 => \_gnd_net_\,
            in3 => \N__20823\,
            lcout => \uu2.un28_w_addr_user_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.r_data_rdy_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010001000"
        )
    port map (
            in0 => \N__14684\,
            in1 => \N__12138\,
            in2 => \N__12114\,
            in3 => \N__25881\,
            lcout => vbuf_tx_data_rdy,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000111111111"
        )
    port map (
            in0 => \N__13409\,
            in1 => \N__13542\,
            in2 => \N__12315\,
            in3 => \N__12303\,
            lcout => \L3_tx_data_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_4_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111100101"
        )
    port map (
            in0 => \N__13678\,
            in1 => \N__22069\,
            in2 => \N__12297\,
            in3 => \N__13410\,
            lcout => \L3_tx_data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12370\,
            in2 => \_gnd_net_\,
            in3 => \N__12354\,
            lcout => \uu0.un99_ci_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_5_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111001110111"
        )
    port map (
            in0 => \N__13408\,
            in1 => \N__13679\,
            in2 => \N__22090\,
            in3 => \N__12288\,
            lcout => \L3_tx_data_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26159\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_1_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011101110111"
        )
    port map (
            in0 => \N__13672\,
            in1 => \N__21195\,
            in2 => \N__22065\,
            in3 => \N__16287\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_2_tz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__13671\,
            in1 => \N__12468\,
            in2 => \_gnd_net_\,
            in3 => \N__12421\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.dOutP_0_iv_1_tz_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_1_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__13403\,
            in1 => \N__13538\,
            in2 => \N__12306\,
            in3 => \N__12267\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_2_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__13536\,
            in1 => \N__12467\,
            in2 => \_gnd_net_\,
            in3 => \N__12420\,
            lcout => \Lab_UT.dispString.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_4_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000101"
        )
    port map (
            in0 => \N__13537\,
            in1 => \N__12469\,
            in2 => \N__13433\,
            in3 => \N__12423\,
            lcout => \Lab_UT.dispString.m74_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_5_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__12422\,
            in1 => \N__13404\,
            in2 => \N__12474\,
            in3 => \N__13539\,
            lcout => \Lab_UT.dispString.m77_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_1_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__12281\,
            in1 => \N__13626\,
            in2 => \N__13688\,
            in3 => \N__21225\,
            lcout => \Lab_UT.dispString.dOutP_0_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_RNISDHD_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12510\,
            in2 => \_gnd_net_\,
            in3 => \N__14718\,
            lcout => \oneSecStrb\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.cnt_RNI7F27_0_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__13535\,
            in1 => \N__12454\,
            in2 => \_gnd_net_\,
            in3 => \N__12408\,
            lcout => \Lab_UT.dispString.N_23_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu0.sec_clkD_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14727\,
            lcout => \uu0.sec_clkDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m57_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100001100"
        )
    port map (
            in0 => \N__17865\,
            in1 => \N__12528\,
            in2 => \N__12419\,
            in3 => \N__12452\,
            lcout => \Lab_UT.m57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m60_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12451\,
            in1 => \N__16720\,
            in2 => \_gnd_net_\,
            in3 => \N__12402\,
            lcout => \G_216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.alarmstate_1_0_i_1_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001000100010"
        )
    port map (
            in0 => \N__12407\,
            in1 => \N__12579\,
            in2 => \N__12473\,
            in3 => \N__17864\,
            lcout => OPEN,
            ltout => \Lab_UT.alarmstate_1_0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_1_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__12418\,
            in1 => \N__12492\,
            in2 => \N__12504\,
            in3 => \N__12498\,
            lcout => \G_215\,
            ltout => \G_215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.alarmstate_1_sqmuxa_1_i_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16719\,
            in2 => \N__12501\,
            in3 => \N__12450\,
            lcout => \G_214\,
            ltout => \G_214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.alarmstate_latch_0_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__12453\,
            in1 => \N__12491\,
            in2 => \N__12483\,
            in3 => \N__12480\,
            lcout => \G_213\,
            ltout => \G_213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_3_0_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101111"
        )
    port map (
            in0 => \N__12406\,
            in1 => \_gnd_net_\,
            in2 => \N__12375\,
            in3 => \N__13555\,
            lcout => \Lab_UT.dispString.N_166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m71_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__25899\,
            in1 => \N__26693\,
            in2 => \N__12624\,
            in3 => \N__13995\,
            lcout => \N_105_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m54_e_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__14952\,
            in1 => \N__14893\,
            in2 => \_gnd_net_\,
            in3 => \N__12527\,
            lcout => \Lab_UT.dispString.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNI0RBN1_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__19720\,
            in1 => \N__13773\,
            in2 => \N__18157\,
            in3 => \N__22977\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_12_a6_3_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNI70I48_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__12573\,
            in1 => \N__17193\,
            in2 => \N__12567\,
            in3 => \N__12564\,
            lcout => \Lab_UT.dictrl.g0_12_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI0UI65_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011001000"
        )
    port map (
            in0 => \N__12558\,
            in1 => \N__12633\,
            in2 => \N__24547\,
            in3 => \N__12552\,
            lcout => \Lab_UT.dictrl.N_23_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_esr_RNINKC83_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__12642\,
            in1 => \N__18630\,
            in2 => \N__15096\,
            in3 => \N__16833\,
            lcout => \Lab_UT.dictrl.state_ret_10_esr_RNINKCZ0Z83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_19_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19422\,
            in1 => \N__15627\,
            in2 => \N__20375\,
            in3 => \N__20283\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_11_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110000"
        )
    port map (
            in0 => \N__18650\,
            in1 => \N__26371\,
            in2 => \N__12546\,
            in3 => \N__18559\,
            lcout => \Lab_UT.dictrl.m63_d_0_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m107_e_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19421\,
            in1 => \N__20282\,
            in2 => \N__12903\,
            in3 => \N__18649\,
            lcout => \Lab_UT.dispString.N_112_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_RNI3S8S_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15336\,
            in1 => \N__15628\,
            in2 => \N__14834\,
            in3 => \N__14057\,
            lcout => \Lab_UT.dictrl.g0_12_a6_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_12_o6_1_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__25501\,
            in1 => \N__26667\,
            in2 => \N__18919\,
            in3 => \N__13990\,
            lcout => \Lab_UT.dictrl.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_1_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000101110011"
        )
    port map (
            in0 => \N__26668\,
            in1 => \N__26372\,
            in2 => \N__22820\,
            in3 => \N__25502\,
            lcout => \Lab_UT.dictrl.N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFP8P_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__15629\,
            in1 => \N__14824\,
            in2 => \_gnd_net_\,
            in3 => \N__17093\,
            lcout => \Lab_UT.dictrl.m27_d_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_7_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__19445\,
            in1 => \N__15630\,
            in2 => \N__15342\,
            in3 => \N__18232\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_a7_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000101"
        )
    port map (
            in0 => \N__16832\,
            in1 => \N__18346\,
            in2 => \N__24053\,
            in3 => \N__14828\,
            lcout => \Lab_UT.dictrl.N_1110_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0H5_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__14825\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24003\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_2_rep1_esr_RNIO0HZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDC4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__15528\,
            in1 => \N__18347\,
            in2 => \N__12636\,
            in3 => \N__14481\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2HDCZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_1_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14826\,
            in1 => \N__24004\,
            in2 => \N__18348\,
            in3 => \N__16830\,
            lcout => \Lab_UT.dictrl.G_17_i_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_RNI2B7F_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16831\,
            in1 => \N__18345\,
            in2 => \N__24054\,
            in3 => \N__14827\,
            lcout => OPEN,
            ltout => \G_17_i_a5_2_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_1_rep2_RNI1CHAB_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__12804\,
            in1 => \N__12798\,
            in2 => \N__12786\,
            in3 => \N__12849\,
            lcout => \G_17_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_e_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12779\,
            in2 => \_gnd_net_\,
            in3 => \N__12752\,
            lcout => \Lab_UT.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_9_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__12710\,
            in1 => \N__12670\,
            in2 => \_gnd_net_\,
            in3 => \N__15411\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_7_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110001"
        )
    port map (
            in0 => \N__14333\,
            in1 => \N__18337\,
            in2 => \N__12735\,
            in3 => \N__12732\,
            lcout => \Lab_UT.dictrl.m53_d_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_10_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__14149\,
            in1 => \N__13002\,
            in2 => \N__14107\,
            in3 => \N__14282\,
            lcout => \Lab_UT.dictrl.g2_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_9_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__15412\,
            in1 => \_gnd_net_\,
            in2 => \N__12682\,
            in3 => \N__12711\,
            lcout => \Lab_UT.dictrl.g2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_9_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__12709\,
            in1 => \N__12669\,
            in2 => \_gnd_net_\,
            in3 => \N__15410\,
            lcout => \Lab_UT.dictrl.g2_0_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_9_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__15413\,
            in1 => \_gnd_net_\,
            in2 => \N__12683\,
            in3 => \N__12712\,
            lcout => \Lab_UT.dictrl.g2_0_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIMUEI_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__12708\,
            in1 => \N__12668\,
            in2 => \_gnd_net_\,
            in3 => \N__15606\,
            lcout => \Lab_UT.dictrl.g2_0_3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m107_e_3_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14150\,
            in1 => \N__14056\,
            in2 => \N__12888\,
            in3 => \N__14276\,
            lcout => \Lab_UT.dispString.m107_eZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m18_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__12827\,
            in1 => \N__12889\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.N_19_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m12_1_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__12891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12828\,
            lcout => \Lab_UT.dictrl.m12Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_i_m2_1_o6_0_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__14094\,
            in1 => \N__12890\,
            in2 => \N__12833\,
            in3 => \N__14277\,
            lcout => \Lab_UT.dictrl.N_10_1\,
            ltout => \Lab_UT.dictrl.N_10_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNI5GLB2_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15631\,
            in1 => \N__18759\,
            in2 => \N__12867\,
            in3 => \N__24002\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_1_a6_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI60US8_0_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__12864\,
            in1 => \N__13014\,
            in2 => \N__12852\,
            in3 => \N__12957\,
            lcout => \N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_21_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__15632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18341\,
            lcout => \Lab_UT.dictrl.N_1105_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI12QU_3_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__20394\,
            in1 => \N__12834\,
            in2 => \N__18603\,
            in3 => \N__15421\,
            lcout => \Lab_UT.dictrl.state_0_fast_esr_RNI12QUZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIB5Q7_0_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__24000\,
            in1 => \_gnd_net_\,
            in2 => \N__15422\,
            in3 => \N__16601\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_1_a6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIF3PO3_0_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110100000"
        )
    port map (
            in0 => \N__13023\,
            in1 => \N__12968\,
            in2 => \N__13017\,
            in3 => \N__13008\,
            lcout => \Lab_UT.dictrl.g0_i_m2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNITRQM_2_LC_5_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__23999\,
            in1 => \N__13001\,
            in2 => \N__15423\,
            in3 => \N__15366\,
            lcout => \Lab_UT.dictrl.g0_i_m2_1_a6_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIO0FK_3_LC_5_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13000\,
            in1 => \N__15414\,
            in2 => \_gnd_net_\,
            in3 => \N__24001\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_1_a6_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIQTO82_0_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12969\,
            in1 => \N__16602\,
            in2 => \N__12960\,
            in3 => \N__14487\,
            lcout => \Lab_UT.dictrl.G_17_i_a5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_11_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__13238\,
            in1 => \N__15775\,
            in2 => \N__12930\,
            in3 => \N__14522\,
            lcout => \uu2.mem0.N_66_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_13_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__15773\,
            in1 => \N__12929\,
            in2 => \_gnd_net_\,
            in3 => \N__13200\,
            lcout => \uu2.mem0.N_56_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI1R353_0_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__23488\,
            in1 => \N__23362\,
            in2 => \N__14568\,
            in3 => \N__23403\,
            lcout => \uu2.N_95_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI1R353_0_0_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__23402\,
            in1 => \N__14563\,
            in2 => \N__23373\,
            in3 => \N__23489\,
            lcout => \uu2.N_96_mux\,
            ltout => \uu2.N_96_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_12_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13161\,
            in1 => \_gnd_net_\,
            in2 => \N__12918\,
            in3 => \N__15774\,
            lcout => \uu2.mem0.N_63_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_9_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111001010100"
        )
    port map (
            in0 => \N__15776\,
            in1 => \N__13128\,
            in2 => \N__14526\,
            in3 => \N__13179\,
            lcout => \uu2.mem0.N_69_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__13127\,
            in1 => \N__13287\,
            in2 => \_gnd_net_\,
            in3 => \N__15777\,
            lcout => \uu2.mem0.N_71_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_15_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23404\,
            in1 => \N__14567\,
            in2 => \_gnd_net_\,
            in3 => \N__23487\,
            lcout => \uu2.mem0.N_91_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_14_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__23592\,
            in1 => \N__13110\,
            in2 => \N__23706\,
            in3 => \N__13266\,
            lcout => \uu2.mem0.N_50_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_2_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__20762\,
            in1 => \N__23697\,
            in2 => \N__13088\,
            in3 => \N__23590\,
            lcout => \uu2.mem0.w_addr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_3_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__23591\,
            in1 => \N__21013\,
            in2 => \N__23705\,
            in3 => \N__17413\,
            lcout => \uu2.mem0.w_addr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIB6L01_4_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__20761\,
            in1 => \_gnd_net_\,
            in2 => \N__17420\,
            in3 => \N__17374\,
            lcout => \uu2.N_75_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNO_0_4_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__23473\,
            in1 => \N__20763\,
            in2 => \N__23380\,
            in3 => \N__25028\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_4_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__17414\,
            in1 => \_gnd_net_\,
            in2 => \N__13026\,
            in3 => \N__17375\,
            lcout => \uu2.w_addr_displayingZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__25767\
        );

    \uu2.w_addr_displaying_RNI2HHB1_4_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011100000"
        )
    port map (
            in0 => \N__23472\,
            in1 => \N__17409\,
            in2 => \N__17381\,
            in3 => \N__20760\,
            lcout => \uu2.bitmap_pmux_sn_N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_2_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__25029\,
            in1 => \N__23474\,
            in2 => \N__17377\,
            in3 => \N__23372\,
            lcout => \uu2.w_addr_displayingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_4C_net\,
            ce => 'H',
            sr => \N__25767\
        );

    \uu2.un1_w_user_lf_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13193\,
            in1 => \N__13212\,
            in2 => \N__13239\,
            in3 => \N__13175\,
            lcout => \uu2.un1_w_user_lf_0\,
            ltout => \uu2.un1_w_user_lf_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI93NG7_2_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23642\,
            in1 => \N__17468\,
            in2 => \N__13215\,
            in3 => \N__23578\,
            lcout => \uu2.un28_w_addr_user_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un1_w_user_lf_4_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13261\,
            in1 => \N__13157\,
            in2 => \N__13286\,
            in3 => \N__13298\,
            lcout => \uu2.un1_w_user_lfZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNI43E87_2_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__25872\,
            in1 => \N__13206\,
            in2 => \N__17472\,
            in3 => \N__23579\,
            lcout => \uu2.w_addr_user_RNI43E87Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.m35_4_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__13192\,
            in1 => \N__13297\,
            in2 => \N__13265\,
            in3 => \N__13174\,
            lcout => OPEN,
            ltout => \uu2.m35Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.m35_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__13156\,
            in1 => \N__13234\,
            in2 => \N__13143\,
            in3 => \N__13279\,
            lcout => \uu2.un1_w_user_cr_0\,
            ltout => \uu2.un1_w_user_cr_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.un4_w_user_data_rdy_0_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13140\,
            in3 => \N__23641\,
            lcout => \uu2.un4_w_user_data_rdyZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_10_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13299\,
            in1 => \N__23662\,
            in2 => \_gnd_net_\,
            in3 => \N__23580\,
            lcout => \uu2.mem0.w_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_2_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001111"
        )
    port map (
            in0 => \N__13569\,
            in1 => \N__13308\,
            in2 => \N__13454\,
            in3 => \N__17832\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_2_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13701\,
            in2 => \N__13302\,
            in3 => \N__13617\,
            lcout => \L3_tx_data_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.rdy_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13570\,
            in1 => \N__22089\,
            in2 => \N__13455\,
            in3 => \N__13704\,
            lcout => \L3_tx_data_rdy\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_0_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111011101"
        )
    port map (
            in0 => \N__13584\,
            in1 => \N__13703\,
            in2 => \_gnd_net_\,
            in3 => \N__13338\,
            lcout => \L3_tx_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_6_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__13702\,
            in1 => \N__13447\,
            in2 => \_gnd_net_\,
            in3 => \N__13608\,
            lcout => \L3_tx_data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26149\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_3_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101001110111"
        )
    port map (
            in0 => \N__13545\,
            in1 => \N__21852\,
            in2 => \N__16347\,
            in3 => \N__13415\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m82_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_3_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__14757\,
            in1 => \N__13546\,
            in2 => \N__13245\,
            in3 => \N__22052\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.N_156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_3_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13687\,
            in2 => \N__13242\,
            in3 => \N__13593\,
            lcout => \L3_tx_data_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_4_1_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__13414\,
            in1 => \N__13544\,
            in2 => \N__13700\,
            in3 => \N__21624\,
            lcout => \Lab_UT.dispString.b1_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_2_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010100101111"
        )
    port map (
            in0 => \N__13574\,
            in1 => \N__17850\,
            in2 => \N__13451\,
            in3 => \N__21650\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m67_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_2_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000001010"
        )
    port map (
            in0 => \N__13573\,
            in1 => \N__22035\,
            in2 => \N__13620\,
            in3 => \N__16307\,
            lcout => \Lab_UT.dispString.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_3_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011001111"
        )
    port map (
            in0 => \N__13575\,
            in1 => \N__13604\,
            in2 => \N__13452\,
            in3 => \N__15996\,
            lcout => \Lab_UT.dispString.N_158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_2_0_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001011111"
        )
    port map (
            in0 => \N__13571\,
            in1 => \N__21375\,
            in2 => \N__16500\,
            in3 => \N__13434\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m90_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_0_0_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001111110011"
        )
    port map (
            in0 => \N__22034\,
            in1 => \N__13572\,
            in2 => \N__13587\,
            in3 => \N__16471\,
            lcout => \Lab_UT.dispString.N_164\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.dOut_RNO_1_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100001011"
        )
    port map (
            in0 => \N__13568\,
            in1 => \N__18003\,
            in2 => \N__13453\,
            in3 => \N__13344\,
            lcout => \Lab_UT.dispString.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_6_rep1_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18151\,
            lcout => bu_rx_data_6_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26127\,
            ce => \N__14243\,
            sr => \N__25826\
        );

    \Lab_UT.dictrl.g1_0_3_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__20487\,
            in1 => \N__17111\,
            in2 => \N__13885\,
            in3 => \N__19439\,
            lcout => \Lab_UT_dictrl_g1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_8_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14006\,
            in1 => \N__17631\,
            in2 => \_gnd_net_\,
            in3 => \N__14369\,
            lcout => \Lab_UT.dictrl.next_state_RNO_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI6DFS_0_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__13954\,
            in1 => \N__17112\,
            in2 => \N__13884\,
            in3 => \N__16600\,
            lcout => \Lab_UT.dictrl.g0_12_a6_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep2_esr_RNIGV0QF_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__16449\,
            in1 => \N__13764\,
            in2 => \N__14844\,
            in3 => \N__13755\,
            lcout => \Lab_UT.dictrl.g2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m15_1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__13955\,
            in1 => \_gnd_net_\,
            in2 => \N__13886\,
            in3 => \N__17113\,
            lcout => \Lab_UT.dictrl.m15Z0Z_1\,
            ltout => \Lab_UT.dictrl.m15Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_esr_RNIMOKF2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__15086\,
            in1 => \N__17630\,
            in2 => \N__13749\,
            in3 => \N__14368\,
            lcout => \Lab_UT.dictrl.m27_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_1_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__13746\,
            in1 => \N__18960\,
            in2 => \N__13734\,
            in3 => \N__13710\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_1_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23083\,
            in2 => \N__13737\,
            in3 => \N__15002\,
            lcout => \Lab_UT.dictrl.next_state_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26121\,
            ce => \N__16884\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_3_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__24484\,
            in1 => \N__22750\,
            in2 => \_gnd_net_\,
            in3 => \N__24278\,
            lcout => \Lab_UT.dictrl.N_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_1_1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18909\,
            in1 => \N__18150\,
            in2 => \N__13725\,
            in3 => \N__24279\,
            lcout => \Lab_UT.dictrl.g0_i_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep2_esr_RNISOI03_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19331\,
            in1 => \N__24458\,
            in2 => \N__14013\,
            in3 => \N__13991\,
            lcout => \Lab_UT.dictrl.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m12_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__20498\,
            in1 => \N__20075\,
            in2 => \N__18763\,
            in3 => \N__14350\,
            lcout => \Lab_UT.dictrl.N_88_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_11_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__18740\,
            in1 => \N__20497\,
            in2 => \N__20091\,
            in3 => \N__20310\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_9_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__13893\,
            in1 => \N__14351\,
            in2 => \N__13974\,
            in3 => \N__19332\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m53_d_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_6_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001110011"
        )
    port map (
            in0 => \N__22818\,
            in1 => \N__24459\,
            in2 => \N__13971\,
            in3 => \N__24345\,
            lcout => \Lab_UT.dictrl.N_1102_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_10_0_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18626\,
            in1 => \N__18920\,
            in2 => \_gnd_net_\,
            in3 => \N__24521\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_5_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__24522\,
            in1 => \N__24292\,
            in2 => \N__13968\,
            in3 => \N__19366\,
            lcout => \Lab_UT.dictrl.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_10_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__13875\,
            in1 => \N__13965\,
            in2 => \_gnd_net_\,
            in3 => \N__15624\,
            lcout => \Lab_UT.dictrl.g2_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_9_0_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__13876\,
            in1 => \N__20502\,
            in2 => \N__13797\,
            in3 => \N__20297\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m59_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_3_0_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100111111"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__19380\,
            in2 => \N__14184\,
            in3 => \N__24524\,
            lcout => \Lab_UT.dictrl.next_state_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_7_0_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__24523\,
            in1 => \_gnd_net_\,
            in2 => \N__18937\,
            in3 => \N__18625\,
            lcout => \Lab_UT.dictrl.m63_d_0_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g2_0_10_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__14278\,
            in1 => \N__14153\,
            in2 => \N__14121\,
            in3 => \N__14060\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_4_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNI2LLA3_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000110011"
        )
    port map (
            in0 => \N__14181\,
            in1 => \N__18321\,
            in2 => \N__14175\,
            in3 => \N__14329\,
            lcout => \Lab_UT.dictrl.m53_d_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_10_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__14279\,
            in1 => \N__14152\,
            in2 => \N__14122\,
            in3 => \N__14059\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_4_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_7_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__18322\,
            in1 => \N__14172\,
            in2 => \N__14166\,
            in3 => \N__14330\,
            lcout => \Lab_UT.dictrl.m53_d_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_10_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__14280\,
            in1 => \N__14151\,
            in2 => \N__14123\,
            in3 => \N__14058\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_7_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__18323\,
            in1 => \N__14163\,
            in2 => \N__14157\,
            in3 => \N__14331\,
            lcout => \Lab_UT.dictrl.m53_d_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_10_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__14281\,
            in1 => \N__14154\,
            in2 => \N__14124\,
            in3 => \N__14061\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_7_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__18324\,
            in1 => \N__14382\,
            in2 => \N__14376\,
            in3 => \N__14332\,
            lcout => \Lab_UT.dictrl.m53_d_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNIMGCH_0_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16599\,
            in2 => \_gnd_net_\,
            in3 => \N__14283\,
            lcout => \Lab_UT.dictrl.N_11_1\,
            ltout => \Lab_UT.dictrl.N_11_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_12_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__14835\,
            in1 => \N__15625\,
            in2 => \N__14295\,
            in3 => \N__24048\,
            lcout => \Lab_UT.dictrl.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_4_0_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19368\,
            in1 => \_gnd_net_\,
            in2 => \N__15700\,
            in3 => \N__14292\,
            lcout => \Lab_UT.dictrl.next_state_RNO_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOF_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18338\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15626\,
            lcout => \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0\,
            ltout => \Lab_UT.dictrl.state_0_3_rep1_esr_RNIBOOFZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNI4DA69_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__15692\,
            in1 => \N__24588\,
            in2 => \N__14286\,
            in3 => \N__22978\,
            lcout => \Lab_UT.dictrl.N_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.shifter_fast_6_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18156\,
            lcout => bu_rx_data_fast_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26117\,
            ce => \N__14237\,
            sr => \N__25841\
        );

    \Lab_UT.dictrl.next_state_RNO_1_0_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14457\,
            in1 => \N__22821\,
            in2 => \_gnd_net_\,
            in3 => \N__14214\,
            lcout => \Lab_UT.dictrl.next_state_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_0_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100011001"
        )
    port map (
            in0 => \N__22822\,
            in1 => \N__24324\,
            in2 => \N__14205\,
            in3 => \N__14193\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.m67_am_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_0_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110101"
        )
    port map (
            in0 => \N__14514\,
            in1 => \N__14508\,
            in2 => \N__14499\,
            in3 => \N__22823\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_0_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__23138\,
            in1 => \_gnd_net_\,
            in2 => \N__14496\,
            in3 => \N__14493\,
            lcout => \Lab_UT.dictrl.next_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26115\,
            ce => \N__16899\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_1_2_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110100000"
        )
    port map (
            in0 => \N__24321\,
            in1 => \N__24552\,
            in2 => \N__14480\,
            in3 => \N__22824\,
            lcout => \Lab_UT.dictrl.next_state_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI2USJ_1_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101000100"
        )
    port map (
            in0 => \N__15452\,
            in1 => \N__24040\,
            in2 => \_gnd_net_\,
            in3 => \N__15060\,
            lcout => \Lab_UT.dictrl.G_17_i_a5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_RNIVHI53_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15623\,
            in1 => \N__19951\,
            in2 => \N__18604\,
            in3 => \N__20143\,
            lcout => \Lab_UT.dictrl.N_65\,
            ltout => \Lab_UT.dictrl.N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_6_0_LC_6_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__24551\,
            in1 => \N__15701\,
            in2 => \N__14460\,
            in3 => \N__24320\,
            lcout => \Lab_UT.dictrl.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__23680\,
            in1 => \N__23607\,
            in2 => \N__21049\,
            in3 => \N__23291\,
            lcout => \uu2.mem0.w_addr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__23608\,
            in1 => \N__23676\,
            in2 => \N__20881\,
            in3 => \N__24957\,
            lcout => \uu2.mem0.w_addr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__25101\,
            in1 => \N__14424\,
            in2 => \N__23693\,
            in3 => \N__23609\,
            lcout => \uu2.mem0.w_addr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI90ME1_0_6_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23290\,
            in1 => \N__25100\,
            in2 => \N__25173\,
            in3 => \N__24955\,
            lcout => \uu2.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI90ME1_6_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111111111"
        )
    port map (
            in0 => \N__24956\,
            in1 => \N__25167\,
            in2 => \N__25104\,
            in3 => \N__23289\,
            lcout => OPEN,
            ltout => \uu2.N_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNIASN45_LC_7_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110100001001"
        )
    port map (
            in0 => \N__17322\,
            in1 => \N__17433\,
            in2 => \N__14553\,
            in3 => \N__15732\,
            lcout => \uu2.bitmap_pmux_sn_i7_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIQBDM1_111_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111011"
        )
    port map (
            in0 => \N__14696\,
            in1 => \N__25076\,
            in2 => \N__14595\,
            in3 => \N__15720\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_26_i_m2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI3JIM3_111_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110000101100"
        )
    port map (
            in0 => \N__25077\,
            in1 => \N__14697\,
            in2 => \N__14550\,
            in3 => \N__14607\,
            lcout => OPEN,
            ltout => \uu2.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIE0KH9_111_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14547\,
            in2 => \N__14538\,
            in3 => \N__20799\,
            lcout => OPEN,
            ltout => \uu2.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIPFVGP_0_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__14535\,
            in1 => \N__17664\,
            in2 => \N__14529\,
            in3 => \N__15726\,
            lcout => \uu2.bitmap_pmux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_296_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__16533\,
            in1 => \N__15504\,
            in2 => \N__16422\,
            in3 => \N__16376\,
            lcout => \uu2.bitmapZ0Z_296\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_200_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__16375\,
            in1 => \N__16408\,
            in2 => \N__15514\,
            in3 => \N__16532\,
            lcout => \uu2.bitmapZ0Z_200\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_72_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__16535\,
            in1 => \N__15506\,
            in2 => \N__16424\,
            in3 => \N__16378\,
            lcout => \uu2.bitmapZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_168_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001011000011110"
        )
    port map (
            in0 => \N__16374\,
            in1 => \N__16407\,
            in2 => \N__15513\,
            in3 => \N__16531\,
            lcout => \uu2.bitmapZ0Z_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_40_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011001111101"
        )
    port map (
            in0 => \N__16534\,
            in1 => \N__15505\,
            in2 => \N__16423\,
            in3 => \N__16377\,
            lcout => \uu2.bitmapZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_RNIQS1B1_40_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__20673\,
            in1 => \N__14622\,
            in2 => \N__14616\,
            in3 => \N__14733\,
            lcout => \uu2.N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNISSSN_162_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14577\,
            in1 => \N__20672\,
            in2 => \_gnd_net_\,
            in3 => \N__14601\,
            lcout => \uu2.N_195\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_75_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110101010111"
        )
    port map (
            in0 => \N__16379\,
            in1 => \N__16418\,
            in2 => \N__15515\,
            in3 => \N__16536\,
            lcout => \uu2.bitmapZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_296C_net\,
            ce => 'H',
            sr => \N__25768\
        );

    \uu2.bitmap_66_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000111101"
        )
    port map (
            in0 => \N__15826\,
            in1 => \N__15964\,
            in2 => \N__15881\,
            in3 => \N__15924\,
            lcout => \uu2.bitmapZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_66C_net\,
            ce => 'H',
            sr => \N__25766\
        );

    \uu2.bitmap_RNIIGUI_66_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14583\,
            in1 => \N__21126\,
            in2 => \_gnd_net_\,
            in3 => \N__14646\,
            lcout => \uu2.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_162_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100111100"
        )
    port map (
            in0 => \N__15825\,
            in1 => \N__15963\,
            in2 => \N__15880\,
            in3 => \N__15923\,
            lcout => \uu2.bitmapZ0Z_162\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_66C_net\,
            ce => 'H',
            sr => \N__25766\
        );

    \uu2.bitmap_RNIHL2N_34_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__24889\,
            in1 => \N__20676\,
            in2 => \N__14640\,
            in3 => \N__14628\,
            lcout => \uu2.bitmap_pmux_15_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_69_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011100011111"
        )
    port map (
            in0 => \N__15925\,
            in1 => \N__15874\,
            in2 => \N__15971\,
            in3 => \N__15827\,
            lcout => \uu2.bitmapZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_66C_net\,
            ce => 'H',
            sr => \N__25766\
        );

    \uu2.bitmap_111_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14726\,
            lcout => \uu2.bitmapZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \uu2.vram_rd_clk_det_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14685\,
            lcout => \uu2.vram_rd_clk_detZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \uu2.vram_rd_clk_det_1_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16023\,
            lcout => \uu2.vram_rd_clk_detZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \uu2.bitmap_194_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__15960\,
            in1 => \N__15918\,
            in2 => \N__15878\,
            in3 => \N__15822\,
            lcout => \uu2.bitmapZ0Z_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \uu2.bitmap_34_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__15962\,
            in1 => \N__15922\,
            in2 => \N__15879\,
            in3 => \N__15824\,
            lcout => \uu2.bitmapZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \uu2.bitmap_290_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__15823\,
            in1 => \N__15864\,
            in2 => \N__15929\,
            in3 => \N__15961\,
            lcout => \uu2.bitmapZ0Z_290\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_111C_net\,
            ce => 'H',
            sr => \N__25765\
        );

    \Lab_UT.didp.regrce4.q_esr_0_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_AMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26146\,
            ce => \N__14775\,
            sr => \N__25804\
        );

    \Lab_UT.didp.regrce4.q_esr_1_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25521\,
            lcout => \Lab_UT.di_AMtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26146\,
            ce => \N__14775\,
            sr => \N__25804\
        );

    \Lab_UT.didp.regrce4.q_esr_2_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26723\,
            lcout => \Lab_UT.di_AMtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26146\,
            ce => \N__14775\,
            sr => \N__25804\
        );

    \Lab_UT.didp.regrce4.q_esr_3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_AMtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26146\,
            ce => \N__14775\,
            sr => \N__25804\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__18411\,
            in1 => \N__26420\,
            in2 => \N__14742\,
            in3 => \N__22213\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_3_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__22178\,
            in1 => \N__22209\,
            in2 => \N__14760\,
            in3 => \N__18372\,
            lcout => \Lab_UT.di_Mtens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__26231\,
            in1 => \N__21847\,
            in2 => \N__22214\,
            in3 => \N__14755\,
            lcout => \Lab_UT.dispString.m49Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNITK144_3_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14756\,
            in1 => \N__22208\,
            in2 => \_gnd_net_\,
            in3 => \N__21344\,
            lcout => \Lab_UT.min1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNIR6J44_3_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21343\,
            in1 => \_gnd_net_\,
            in2 => \N__26235\,
            in3 => \N__21848\,
            lcout => \Lab_UT.min2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__21914\,
            in1 => \N__22281\,
            in2 => \_gnd_net_\,
            in3 => \N__21971\,
            lcout => \Lab_UT.didp.countrce4.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__22425\,
            in1 => \N__22380\,
            in2 => \N__22467\,
            in3 => \N__22968\,
            lcout => \Lab_UT.dictrl.state_1_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26132\,
            ce => \N__22487\,
            sr => \N__25799\
        );

    \Lab_UT.dictrl.state_0_2_rep2_esr_RNI3AA01_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__19779\,
            in1 => \_gnd_net_\,
            in2 => \N__19330\,
            in3 => \N__23084\,
            lcout => \Lab_UT.dictrl.g0_12_a6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_4_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19317\,
            in2 => \_gnd_net_\,
            in3 => \N__19778\,
            lcout => \Lab_UT.dictrl.g2_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNINE144_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16475\,
            in1 => \N__21301\,
            in2 => \_gnd_net_\,
            in3 => \N__21970\,
            lcout => \Lab_UT.min1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIPG144_1_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21302\,
            in1 => \N__22279\,
            in2 => \_gnd_net_\,
            in3 => \N__16282\,
            lcout => \Lab_UT.min1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce4.q_esr_RNIRI144_2_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21326\,
            in1 => \N__21907\,
            in2 => \_gnd_net_\,
            in3 => \N__16308\,
            lcout => \Lab_UT.min1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI56JGE_1_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__15044\,
            in1 => \N__24032\,
            in2 => \N__23163\,
            in3 => \N__15248\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110001"
        )
    port map (
            in0 => \N__24034\,
            in1 => \N__23152\,
            in2 => \N__15258\,
            in3 => \N__15048\,
            lcout => \Lab_UT.dictrl.state_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_0_2_rep1_esr_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__15045\,
            in1 => \N__24037\,
            in2 => \N__23164\,
            in3 => \N__15249\,
            lcout => \Lab_UT.dictrl.state_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_0_2_rep2_esr_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000011110001"
        )
    port map (
            in0 => \N__24033\,
            in1 => \N__23148\,
            in2 => \N__15257\,
            in3 => \N__15046\,
            lcout => \Lab_UT.dictrl.state_2_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_0_esr_2_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__15047\,
            in1 => \N__24038\,
            in2 => \N__23165\,
            in3 => \N__15253\,
            lcout => \Lab_UT.dictrl.stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_ret_1_ess_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000111000011111"
        )
    port map (
            in0 => \N__24035\,
            in1 => \N__23153\,
            in2 => \N__15021\,
            in3 => \N__15006\,
            lcout => \Lab_UT.dictrl.state_i_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNI7ECM_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__18199\,
            in1 => \N__19767\,
            in2 => \N__14985\,
            in3 => \N__19617\,
            lcout => \Lab_UT.LdASones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0001111100001110"
        )
    port map (
            in0 => \N__24036\,
            in1 => \N__23154\,
            in2 => \N__15168\,
            in3 => \N__14976\,
            lcout => \Lab_UT.state_i_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26129\,
            ce => \N__22488\,
            sr => \N__25802\
        );

    \Lab_UT.dictrl.state_ret_12_RNIRIHQ6_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100111000"
        )
    port map (
            in0 => \N__15151\,
            in1 => \N__16978\,
            in2 => \N__24049\,
            in3 => \N__15130\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNI2MD42_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25874\,
            in1 => \N__14964\,
            in2 => \N__24052\,
            in3 => \N__14898\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNIROSR8_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010000000"
        )
    port map (
            in0 => \N__15152\,
            in1 => \N__16979\,
            in2 => \N__14856\,
            in3 => \N__15131\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI71KU22_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__22587\,
            in1 => \N__14853\,
            in2 => \N__14847\,
            in3 => \N__23191\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNI71KU22Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100111000"
        )
    port map (
            in0 => \N__15156\,
            in1 => \N__16987\,
            in2 => \N__24051\,
            in3 => \N__15133\,
            lcout => \Lab_UT.dictrl.state_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26125\,
            ce => \N__22490\,
            sr => \N__25803\
        );

    \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101001010"
        )
    port map (
            in0 => \N__23997\,
            in1 => \N__15153\,
            in2 => \N__16988\,
            in3 => \N__15134\,
            lcout => \Lab_UT.dictrl.state_3_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26125\,
            ce => \N__22490\,
            sr => \N__25803\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100111000"
        )
    port map (
            in0 => \N__15154\,
            in1 => \N__16983\,
            in2 => \N__24050\,
            in3 => \N__15132\,
            lcout => \Lab_UT.dictrl.state_3_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26125\,
            ce => \N__22490\,
            sr => \N__25803\
        );

    \Lab_UT.dictrl.state_0_esr_3_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101001010"
        )
    port map (
            in0 => \N__23998\,
            in1 => \N__15155\,
            in2 => \N__16989\,
            in3 => \N__15135\,
            lcout => \Lab_UT.state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26125\,
            ce => \N__22490\,
            sr => \N__25803\
        );

    \Lab_UT.dictrl.state_ret_2_ess_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__15068\,
            in1 => \N__15182\,
            in2 => \_gnd_net_\,
            in3 => \N__15665\,
            lcout => \Lab_UT.dictrl.state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26123\,
            ce => \N__22491\,
            sr => \N__25807\
        );

    \Lab_UT.dictrl.state_0_esr_RNIS4PO5_2_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011101"
        )
    port map (
            in0 => \N__22775\,
            in1 => \N__15108\,
            in2 => \N__16440\,
            in3 => \N__24144\,
            lcout => \Lab_UT.dictrl.N_62\,
            ltout => \Lab_UT.dictrl.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_10_esr_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000100000000"
        )
    port map (
            in0 => \N__15069\,
            in1 => \N__15183\,
            in2 => \N__15099\,
            in3 => \N__22551\,
            lcout => \Lab_UT.dictrl.N_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26123\,
            ce => \N__22491\,
            sr => \N__25807\
        );

    \Lab_UT.dictrl.state_0_esr_RNIP2CG_1_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23082\,
            in2 => \_gnd_net_\,
            in3 => \N__23911\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNIP2CGZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_1_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__22420\,
            in1 => \N__22372\,
            in2 => \N__22463\,
            in3 => \N__22945\,
            lcout => \Lab_UT.dictrl.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26123\,
            ce => \N__22491\,
            sr => \N__25807\
        );

    \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__22943\,
            in1 => \N__22421\,
            in2 => \N__22379\,
            in3 => \N__22458\,
            lcout => \Lab_UT.dictrl.state_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26123\,
            ce => \N__22491\,
            sr => \N__25807\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__22419\,
            in1 => \N__22371\,
            in2 => \N__22462\,
            in3 => \N__22944\,
            lcout => \Lab_UT.dictrl.state_1_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26123\,
            ce => \N__22491\,
            sr => \N__25807\
        );

    \Lab_UT.dictrl.state_0_esr_RNIQ2M68_3_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__15267\,
            in1 => \N__15231\,
            in2 => \N__24533\,
            in3 => \N__15200\,
            lcout => \Lab_UT.dictrl.N_1459_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_71_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__18935\,
            in1 => \N__20597\,
            in2 => \N__19193\,
            in3 => \N__20196\,
            lcout => \Lab_UT.dictrl.N_40_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_35_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20197\,
            in1 => \N__19164\,
            in2 => \N__20601\,
            in3 => \N__18936\,
            lcout => \Lab_UT.dictrl.N_40_3\,
            ltout => \Lab_UT.dictrl.N_40_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__24030\,
            in1 => \N__19532\,
            in2 => \N__15225\,
            in3 => \N__24489\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1462_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_2_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__15222\,
            in1 => \N__15216\,
            in2 => \N__15207\,
            in3 => \N__24031\,
            lcout => \Lab_UT.dictrl.N_1460_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNI78VA1_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001111"
        )
    port map (
            in0 => \N__24304\,
            in1 => \N__22777\,
            in2 => \N__24058\,
            in3 => \N__23119\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_esr_RNI78VA1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNITVS29_3_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000111010"
        )
    port map (
            in0 => \N__15204\,
            in1 => \N__15693\,
            in2 => \N__15186\,
            in3 => \N__24491\,
            lcout => \Lab_UT.dictrl.state_0_esr_RNITVS29Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_7_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__24303\,
            in1 => \N__19959\,
            in2 => \N__24057\,
            in3 => \N__22776\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__15441\,
            in1 => \N__17250\,
            in2 => \N__15171\,
            in3 => \N__17292\,
            lcout => \Lab_UT.dictrl.state_ret_5_ess_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_5_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__24490\,
            in1 => \N__15456\,
            in2 => \_gnd_net_\,
            in3 => \N__24017\,
            lcout => \Lab_UT.dictrl.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m23_0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20159\,
            in1 => \N__20580\,
            in2 => \N__20094\,
            in3 => \N__20325\,
            lcout => \Lab_UT.dictrl.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_15_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15399\,
            in1 => \N__15364\,
            in2 => \N__15340\,
            in3 => \N__23963\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_0_a7_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_11_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__20157\,
            in1 => \N__20578\,
            in2 => \N__15435\,
            in3 => \N__20323\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_18_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_4_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__15543\,
            in1 => \N__15432\,
            in2 => \N__15426\,
            in3 => \N__23964\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_18_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__20158\,
            in1 => \N__20579\,
            in2 => \N__18605\,
            in3 => \N__20324\,
            lcout => \Lab_UT.dictrl.N_40_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_14_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15400\,
            in1 => \N__15365\,
            in2 => \N__15341\,
            in3 => \N__23962\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_a7_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__15309\,
            in1 => \N__20215\,
            in2 => \N__15303\,
            in3 => \N__19952\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_22_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_3_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__20232\,
            in1 => \N__15294\,
            in2 => \N__15282\,
            in3 => \N__15279\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_8_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20031\,
            in1 => \N__20214\,
            in2 => \_gnd_net_\,
            in3 => \N__19953\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_97_mux_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_5_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101111"
        )
    port map (
            in0 => \N__15714\,
            in1 => \N__19844\,
            in2 => \N__15705\,
            in3 => \N__19725\,
            lcout => \Lab_UT.dictrl.N_1102_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_2_2_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__24534\,
            in1 => \N__15702\,
            in2 => \N__23166\,
            in3 => \N__15666\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_RNO_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__15642\,
            in1 => \N__23159\,
            in2 => \N__15651\,
            in3 => \N__15648\,
            lcout => \Lab_UT.dictrl.next_state_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26116\,
            ce => \N__16895\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_0_2_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22801\,
            in2 => \_gnd_net_\,
            in3 => \N__24322\,
            lcout => \Lab_UT.dictrl.next_state_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNINV3P_2_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__15607\,
            in1 => \N__15539\,
            in2 => \_gnd_net_\,
            in3 => \N__24041\,
            lcout => \Lab_UT.dictrl.next_state_RNINV3PZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_203_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__16383\,
            in1 => \N__16425\,
            in2 => \N__15516\,
            in3 => \N__16530\,
            lcout => \uu2.bitmapZ0Z_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__25774\
        );

    \uu2.bitmap_RNIPJHV_200_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15471\,
            in1 => \N__17797\,
            in2 => \_gnd_net_\,
            in3 => \N__15465\,
            lcout => \uu2.N_199\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__17800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25020\,
            lcout => \uu2.w_addr_displaying_0_repZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_203C_net\,
            ce => 'H',
            sr => \N__25774\
        );

    \uu2.w_addr_displaying_0_rep1_RNIDASJ_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20742\,
            in2 => \_gnd_net_\,
            in3 => \N__17798\,
            lcout => \uu2.w_addr_displaying_0_rep1_RNIDASJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_rep1_RNI8NUT1_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000100"
        )
    port map (
            in0 => \N__17799\,
            in1 => \N__17565\,
            in2 => \N__17382\,
            in3 => \N__20754\,
            lcout => \uu2.bitmap_pmux_sn_N_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIBTRT7_0_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000011111001"
        )
    port map (
            in0 => \N__23328\,
            in1 => \N__23462\,
            in2 => \N__17751\,
            in3 => \N__17586\,
            lcout => \uu2.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIBP86_2_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20628\,
            in2 => \_gnd_net_\,
            in3 => \N__20661\,
            lcout => \uu2.N_24_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_1_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001100110"
        )
    port map (
            in0 => \N__23330\,
            in1 => \N__23464\,
            in2 => \_gnd_net_\,
            in3 => \N__24999\,
            lcout => \uu2.w_addr_displayingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__25771\
        );

    \uu2.w_addr_displaying_fast_2_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111101000000"
        )
    port map (
            in0 => \N__25001\,
            in1 => \N__23334\,
            in2 => \N__23485\,
            in3 => \N__20629\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__25771\
        );

    \uu2.w_addr_displaying_fast_1_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__20784\,
            in1 => \_gnd_net_\,
            in2 => \N__23343\,
            in3 => \N__25000\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__25771\
        );

    \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000010001"
        )
    port map (
            in0 => \N__20633\,
            in1 => \N__20662\,
            in2 => \_gnd_net_\,
            in3 => \N__20783\,
            lcout => \uu2.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIU1AF7_0_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__23329\,
            in1 => \N__23463\,
            in2 => \_gnd_net_\,
            in3 => \N__24998\,
            lcout => \uu2.w_addr_displaying_RNIU1AF7Z0Z_0\,
            ltout => \uu2.w_addr_displaying_RNIU1AF7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_3_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17654\,
            in2 => \N__15975\,
            in3 => \N__20663\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_1C_net\,
            ce => 'H',
            sr => \N__25771\
        );

    \uu2.bitmap_197_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__15972\,
            in1 => \N__15930\,
            in2 => \N__15885\,
            in3 => \N__15831\,
            lcout => \uu2.bitmapZ0Z_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__25769\
        );

    \uu2.bitmap_RNIOMUI_69_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15789\,
            in1 => \N__21127\,
            in2 => \_gnd_net_\,
            in3 => \N__15783\,
            lcout => \uu2.N_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_7_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110001100110"
        )
    port map (
            in0 => \N__23252\,
            in1 => \N__21132\,
            in2 => \N__25162\,
            in3 => \N__15772\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__25769\
        );

    \uu2.w_addr_displaying_7_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101001100110"
        )
    port map (
            in0 => \N__25088\,
            in1 => \N__23250\,
            in2 => \N__25169\,
            in3 => \N__15769\,
            lcout => \uu2.w_addr_displayingZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__25769\
        );

    \uu2.w_addr_displaying_8_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001011110000"
        )
    port map (
            in0 => \N__23251\,
            in1 => \N__15770\,
            in2 => \N__25163\,
            in3 => \N__25089\,
            lcout => \uu2.w_addr_displayingZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__25769\
        );

    \uu2.w_addr_displaying_RNIHDHP6_8_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__25087\,
            in1 => \N__23249\,
            in2 => \N__25168\,
            in3 => \N__15768\,
            lcout => \uu2.w_addr_displaying_RNIHDHP6Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_8_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100100000"
        )
    port map (
            in0 => \N__25079\,
            in1 => \N__15771\,
            in2 => \N__23256\,
            in3 => \N__24890\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_197C_net\,
            ce => 'H',
            sr => \N__25769\
        );

    \uu2.w_addr_displaying_RNIR2PL_8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25078\,
            in2 => \_gnd_net_\,
            in3 => \N__25136\,
            lcout => \uu2.w_addr_displaying_RNIR2PLZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buart.Z_rx.bitcount_es_2_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100011101110100"
        )
    port map (
            in0 => \N__16254\,
            in1 => \N__16191\,
            in2 => \N__16152\,
            in3 => \N__16103\,
            lcout => \buart__rx_bitcount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26170\,
            ce => \N__16089\,
            sr => \N__25842\
        );

    \uu2.bitmap_RNI71NJ_72_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__16044\,
            in2 => \_gnd_net_\,
            in3 => \N__16038\,
            lcout => \uu2.N_196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.vram_rd_clk_det_RNI95711_1_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16032\,
            in1 => \N__16022\,
            in2 => \_gnd_net_\,
            in3 => \N__25873\,
            lcout => \uu2.vram_rd_clk_det_RNI95711Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_0_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__25222\,
            in1 => \N__16336\,
            in2 => \N__17715\,
            in3 => \N__15988\,
            lcout => \Lab_UT.dispString.m49Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNINAM54_3_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__15989\,
            in1 => \N__21340\,
            in2 => \_gnd_net_\,
            in3 => \N__17711\,
            lcout => \Lab_UT.sec2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNIPO4L3_3_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21341\,
            in1 => \_gnd_net_\,
            in2 => \N__25227\,
            in3 => \N__16337\,
            lcout => \Lab_UT.sec1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26413\,
            lcout => \Lab_UT.di_ASones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26161\,
            ce => \N__18021\,
            sr => \N__25813\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIJ6M54_1_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21336\,
            in1 => \N__21255\,
            in2 => \_gnd_net_\,
            in3 => \N__21190\,
            lcout => \Lab_UT.sec2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_1_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25523\,
            lcout => \Lab_UT.di_ASones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26161\,
            ce => \N__18021\,
            sr => \N__25813\
        );

    \Lab_UT.didp.regrce3.q_esr_RNIN2J44_1_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__21620\,
            in1 => \_gnd_net_\,
            in2 => \N__21348\,
            in3 => \N__26577\,
            lcout => \Lab_UT.min2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNIP4J44_2_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21342\,
            in1 => \N__26499\,
            in2 => \_gnd_net_\,
            in3 => \N__21651\,
            lcout => \Lab_UT.min2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_1_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25522\,
            lcout => \Lab_UT.di_AStens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26153\,
            ce => \N__16323\,
            sr => \N__25809\
        );

    \Lab_UT.didp.regrce2.q_esr_2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26724\,
            lcout => \Lab_UT.di_AStens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26153\,
            ce => \N__16323\,
            sr => \N__25809\
        );

    \Lab_UT.didp.regrce2.q_esr_3_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__26422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_AStens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26153\,
            ce => \N__16323\,
            sr => \N__25809\
        );

    \Lab_UT.didp.regrce2.q_esr_0_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21775\,
            lcout => \Lab_UT.di_AStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26153\,
            ce => \N__16323\,
            sr => \N__25809\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_2_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__18407\,
            in1 => \N__26715\,
            in2 => \N__16677\,
            in3 => \N__21905\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__21906\,
            in1 => \N__22177\,
            in2 => \N__16311\,
            in3 => \N__18371\,
            lcout => \Lab_UT.di_Mtens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_3_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__16303\,
            in1 => \N__22269\,
            in2 => \N__16286\,
            in3 => \N__21904\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m49Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_12_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16557\,
            in1 => \N__16548\,
            in2 => \N__16542\,
            in3 => \N__21588\,
            lcout => \Lab_UT.dispString.m49Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21805\,
            lcout => \Lab_UT.di_AMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26139\,
            ce => \N__21821\,
            sr => \N__25801\
        );

    \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__16644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25878\,
            lcout => \Lab_UT.didp.regrce3.LdAMones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNILRDD3_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18032\,
            in1 => \N__16655\,
            in2 => \N__16628\,
            in3 => \N__16643\,
            lcout => \Lab_UT.loadalarm_0\,
            ltout => \Lab_UT.loadalarm_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_RNIL0J44_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110010101100"
        )
    port map (
            in0 => \N__26538\,
            in1 => \N__16490\,
            in2 => \N__16539\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.min2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_7_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__16489\,
            in1 => \N__26537\,
            in2 => \N__16476\,
            in3 => \N__21948\,
            lcout => \Lab_UT.dispString.m49Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNIAOPO_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__22948\,
            in1 => \N__18287\,
            in2 => \N__19048\,
            in3 => \N__16797\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_12_a6_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNIK3DC4_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__18155\,
            in1 => \N__19198\,
            in2 => \N__16452\,
            in3 => \N__18780\,
            lcout => \Lab_UT.dictrl.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_14_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__19040\,
            in1 => \_gnd_net_\,
            in2 => \N__19210\,
            in3 => \N__18153\,
            lcout => \Lab_UT.dictrl.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNIG5AU_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__18154\,
            in1 => \N__19041\,
            in2 => \N__18224\,
            in3 => \N__19197\,
            lcout => \Lab_UT.dictrl.m35_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22266\,
            in2 => \_gnd_net_\,
            in3 => \N__21952\,
            lcout => \Lab_UT.didp.countrce4.un13_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNI9E421_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__19615\,
            in1 => \N__18170\,
            in2 => \_gnd_net_\,
            in3 => \N__19271\,
            lcout => \Lab_UT.LdAMtens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNI79EL_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__22947\,
            in1 => \N__19616\,
            in2 => \N__18217\,
            in3 => \N__16795\,
            lcout => \Lab_UT.LdAMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNIULEV_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16796\,
            in1 => \N__22946\,
            in2 => \N__19310\,
            in3 => \N__19618\,
            lcout => \Lab_UT.LdAStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000110101"
        )
    port map (
            in0 => \N__16611\,
            in1 => \N__22878\,
            in2 => \N__17229\,
            in3 => \N__22588\,
            lcout => \Lab_UT.dicRun_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__17016\,
            in1 => \N__16860\,
            in2 => \N__17046\,
            in3 => \N__17148\,
            lcout => \Lab_UT.dictrl.state_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__17145\,
            in1 => \N__17037\,
            in2 => \N__16862\,
            in3 => \N__17013\,
            lcout => \Lab_UT.dictrl.state_0_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.state_0_0_rep2_esr_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__17014\,
            in1 => \N__16856\,
            in2 => \N__17045\,
            in3 => \N__17146\,
            lcout => \Lab_UT.dictrl.state_0_rep2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.state_0_esr_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__17147\,
            in1 => \N__17041\,
            in2 => \N__16863\,
            in3 => \N__17015\,
            lcout => \Lab_UT.dictrl.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNIN23OR_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__17144\,
            in1 => \N__17036\,
            in2 => \N__16861\,
            in3 => \N__17012\,
            lcout => \Lab_UT.dictrl.next_stateZ0Z_0\,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__22589\,
            in1 => \N__22552\,
            in2 => \N__16992\,
            in3 => \N__17214\,
            lcout => \Lab_UT.LdStens_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26130\,
            ce => \N__22489\,
            sr => \N__25808\
        );

    \Lab_UT.dictrl.next_state_RNICLDV_3_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__23905\,
            in1 => \N__19305\,
            in2 => \N__16908\,
            in3 => \N__16834\,
            lcout => \Lab_UT.dictrl.next_state_latmux_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_3_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dictrl.next_state_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26126\,
            ce => \N__16894\,
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_RNI4JJN_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__19850\,
            in1 => \N__19306\,
            in2 => \N__24012\,
            in3 => \N__16836\,
            lcout => \Lab_UT.dictrl.G_17_i_a5_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_5_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__16835\,
            in1 => \N__19851\,
            in2 => \N__19329\,
            in3 => \N__23909\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_0_a7_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_2_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__16770\,
            in1 => \N__16761\,
            in2 => \N__16749\,
            in3 => \N__16746\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25926\,
            in1 => \N__16733\,
            in2 => \N__16737\,
            in3 => \N__22550\,
            lcout => \Lab_UT.dictrl.state_ret_12and_0_ns_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_0_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__23910\,
            in1 => \N__25925\,
            in2 => \N__22560\,
            in3 => \N__16734\,
            lcout => \Lab_UT.dictrl.state_ret_12and_0_ns_rn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep1_esr_RNI6TSE1_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__25494\,
            in1 => \N__26687\,
            in2 => \_gnd_net_\,
            in3 => \N__17205\,
            lcout => \Lab_UT.dictrl.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_7_1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__26688\,
            in1 => \N__18927\,
            in2 => \N__26391\,
            in3 => \N__25497\,
            lcout => \Lab_UT.dictrl.g0_i_a4_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_16_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110001111"
        )
    port map (
            in0 => \N__25496\,
            in1 => \N__26370\,
            in2 => \N__18938\,
            in3 => \N__26689\,
            lcout => \Lab_UT.dictrl.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_i_m2_5_N_3L3_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100000000"
        )
    port map (
            in0 => \N__26686\,
            in1 => \N__25495\,
            in2 => \N__26390\,
            in3 => \N__17107\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_5_N_3LZ0Z3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3_3_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011101110111"
        )
    port map (
            in0 => \N__18243\,
            in1 => \N__17165\,
            in2 => \N__17181\,
            in3 => \N__17178\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.state_0_fast_esr_RNI3MHO3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNII5BFA_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__17166\,
            in1 => \N__17244\,
            in2 => \N__17151\,
            in3 => \N__17052\,
            lcout => \Lab_UT.dictrl.N_1792_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep2_esr_RNIQV2R6_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101111"
        )
    port map (
            in0 => \N__19830\,
            in1 => \N__17127\,
            in2 => \N__18432\,
            in3 => \N__19700\,
            lcout => \Lab_UT.dictrl.N_1102_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_16_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20595\,
            in1 => \N__17118\,
            in2 => \N__18606\,
            in3 => \N__20217\,
            lcout => \Lab_UT.dictrl.N_40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_13_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100010001"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__24016\,
            in2 => \N__18939\,
            in3 => \N__19831\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000010100000"
        )
    port map (
            in0 => \N__17262\,
            in1 => \N__20596\,
            in2 => \N__17253\,
            in3 => \N__19316\,
            lcout => \Lab_UT.dictrl.g0_i_m2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_17_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__20218\,
            in2 => \_gnd_net_\,
            in3 => \N__19958\,
            lcout => \Lab_UT.dictrl.N_97_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__24271\,
            in1 => \N__20205\,
            in2 => \N__19211\,
            in3 => \N__23981\,
            lcout => \Lab_UT.dictrl.g0_i_a5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_36_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__19956\,
            in1 => \_gnd_net_\,
            in2 => \N__20221\,
            in3 => \N__19199\,
            lcout => \Lab_UT.dictrl.N_97_mux_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_65_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__20198\,
            in2 => \_gnd_net_\,
            in3 => \N__19954\,
            lcout => \Lab_UT.dictrl.N_97_mux_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m40_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__19955\,
            in1 => \_gnd_net_\,
            in2 => \N__20220\,
            in3 => \N__20078\,
            lcout => \Lab_UT.dictrl.N_97_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_0_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23123\,
            in2 => \_gnd_net_\,
            in3 => \N__23983\,
            lcout => \Lab_UT.dictrl.g2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_2_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__23982\,
            in1 => \_gnd_net_\,
            in2 => \N__23155\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_0_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__17268\,
            in1 => \N__17310\,
            in2 => \N__17217\,
            in3 => \N__22979\,
            lcout => \Lab_UT.dictrl.next_state_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__24294\,
            in1 => \N__19227\,
            in2 => \N__24555\,
            in3 => \N__24578\,
            lcout => \Lab_UT.dictrl.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_4_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__19822\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19314\,
            lcout => \Lab_UT.dictrl.g2_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19311\,
            in2 => \_gnd_net_\,
            in3 => \N__19819\,
            lcout => \Lab_UT.dictrl.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_15_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__19823\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24013\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_m2_i_a6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNO_6_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__19357\,
            in1 => \N__17304\,
            in2 => \N__17295\,
            in3 => \N__24293\,
            lcout => \Lab_UT.dictrl.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_4_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__19821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19313\,
            lcout => \Lab_UT.dictrl.g2_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_4_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19312\,
            in2 => \_gnd_net_\,
            in3 => \N__19820\,
            lcout => \Lab_UT.dictrl.g2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_6_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000001"
        )
    port map (
            in0 => \N__19226\,
            in1 => \N__24014\,
            in2 => \N__19736\,
            in3 => \N__19538\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1462_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_7_ess_RNO_3_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__24015\,
            in1 => \N__17283\,
            in2 => \N__17277\,
            in3 => \N__17274\,
            lcout => \Lab_UT.dictrl.N_1460_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_8_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__20090\,
            in1 => \N__20216\,
            in2 => \_gnd_net_\,
            in3 => \N__19957\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_97_mux_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_5_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101111"
        )
    port map (
            in0 => \N__17580\,
            in1 => \N__19824\,
            in2 => \N__17568\,
            in3 => \N__19724\,
            lcout => \Lab_UT.dictrl.N_1102_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI316V_8_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000001010"
        )
    port map (
            in0 => \N__24894\,
            in1 => \N__23277\,
            in2 => \N__24954\,
            in3 => \N__21135\,
            lcout => \uu2.bitmap_pmux_sn_N_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_nesr_RNI9006_8_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__23543\,
            in1 => \N__20872\,
            in2 => \_gnd_net_\,
            in3 => \N__17558\,
            lcout => OPEN,
            ltout => \uu2.un3_w_addr_user_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_RNIINVH_2_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21015\,
            in1 => \N__17523\,
            in2 => \N__17487\,
            in3 => \N__17484\,
            lcout => \uu2.un3_w_addr_user\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_nesr_5_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__23278\,
            in1 => \N__23418\,
            in2 => \N__23385\,
            in3 => \N__23471\,
            lcout => \uu2.w_addr_displayingZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_nesr_5C_net\,
            ce => \N__17448\,
            sr => \N__25778\
        );

    \uu2.w_addr_displaying_fast_RNI3FPC1_1_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001000010"
        )
    port map (
            in0 => \N__20789\,
            in1 => \N__17367\,
            in2 => \N__17421\,
            in3 => \N__17687\,
            lcout => \uu2.w_addr_displaying_fast_RNI3FPC1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIUO0E_1_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17415\,
            in2 => \_gnd_net_\,
            in3 => \N__20788\,
            lcout => \uu2.bitmap_pmux_sn_N_33\,
            ltout => \uu2.bitmap_pmux_sn_N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIRB2A1_4_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001101010011"
        )
    port map (
            in0 => \N__17419\,
            in1 => \N__17653\,
            in2 => \N__17385\,
            in3 => \N__17366\,
            lcout => \uu2.bitmap_pmux_sn_m15_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIMLNS2_1_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000010000000"
        )
    port map (
            in0 => \N__17688\,
            in1 => \N__20610\,
            in2 => \N__17679\,
            in3 => \N__17670\,
            lcout => \uu2.bitmap_pmux_29_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_3_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17655\,
            in1 => \N__20755\,
            in2 => \_gnd_net_\,
            in3 => \N__17637\,
            lcout => \uu2.w_addr_displayingZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_3C_net\,
            ce => 'H',
            sr => \N__25775\
        );

    \Lab_UT.dictrl.m12_2_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__18764\,
            in1 => \N__20508\,
            in2 => \_gnd_net_\,
            in3 => \N__18587\,
            lcout => \Lab_UT.dictrl.m12Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_215_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111101011011"
        )
    port map (
            in0 => \N__24768\,
            in1 => \N__24741\,
            in2 => \N__24693\,
            in3 => \N__24636\,
            lcout => \uu2.bitmapZ0Z_215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_215C_net\,
            ce => 'H',
            sr => \N__25772\
        );

    \uu2.bitmap_RNIE8OP_212_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__24909\,
            in1 => \N__24828\,
            in2 => \_gnd_net_\,
            in3 => \N__17613\,
            lcout => OPEN,
            ltout => \uu2.N_198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI0SET1_3_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101100111"
        )
    port map (
            in0 => \N__25090\,
            in1 => \N__20743\,
            in2 => \N__17607\,
            in3 => \N__24804\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_27_i_m2_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNIPTJR3_3_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001111010"
        )
    port map (
            in0 => \N__20744\,
            in1 => \N__17604\,
            in2 => \N__17595\,
            in3 => \N__17592\,
            lcout => \uu2.bitmap_pmux_27_i_m2_ns_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_93_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011110011111"
        )
    port map (
            in0 => \N__21409\,
            in1 => \N__21504\,
            in2 => \N__21457\,
            in3 => \N__21550\,
            lcout => \uu2.bitmapZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__25770\
        );

    \uu2.bitmap_221_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100111101"
        )
    port map (
            in0 => \N__21549\,
            in1 => \N__21447\,
            in2 => \N__21513\,
            in3 => \N__21408\,
            lcout => \uu2.bitmapZ0Z_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_93C_net\,
            ce => 'H',
            sr => \N__25770\
        );

    \uu2.w_addr_displaying_0_rep1_RNINHPP1_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__20756\,
            in1 => \N__17805\,
            in2 => \N__17772\,
            in3 => \N__17760\,
            lcout => OPEN,
            ltout => \uu2.bitmap_pmux_25_i_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI5BFC3_3_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__20757\,
            in1 => \N__21147\,
            in2 => \N__17754\,
            in3 => \N__17727\,
            lcout => \uu2.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI95TJ_93_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__17739\,
            in1 => \N__17733\,
            in2 => \_gnd_net_\,
            in3 => \N__21131\,
            lcout => \uu2.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m43_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__21361\,
            in1 => \N__25560\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.dispString.N_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIL8M54_2_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21347\,
            in1 => \N__17900\,
            in2 => \_gnd_net_\,
            in3 => \N__17828\,
            lcout => \Lab_UT.sec2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNI28771_3_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__21256\,
            in1 => \N__17901\,
            in2 => \N__17954\,
            in3 => \N__17712\,
            lcout => \Lab_UT.didp.un18_ce\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_3_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__17902\,
            in1 => \N__17953\,
            in2 => \_gnd_net_\,
            in3 => \N__21258\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110111011000"
        )
    port map (
            in0 => \N__22523\,
            in1 => \N__26412\,
            in2 => \N__17721\,
            in3 => \N__17713\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_3_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__21998\,
            in1 => \N__22643\,
            in2 => \N__17718\,
            in3 => \N__17714\,
            lcout => \Lab_UT.di_Sones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_1_2_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__21257\,
            in1 => \_gnd_net_\,
            in2 => \N__17955\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_2_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__17903\,
            in1 => \N__22522\,
            in2 => \N__17910\,
            in3 => \N__26730\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_2_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__17904\,
            in1 => \N__22642\,
            in2 => \N__17907\,
            in3 => \N__21997\,
            lcout => \Lab_UT.di_Sones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_1_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__22641\,
            in1 => \N__18048\,
            in2 => \N__21999\,
            in3 => \N__21259\,
            lcout => \Lab_UT.di_Sones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_4_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__17899\,
            in1 => \N__17845\,
            in2 => \N__25599\,
            in3 => \N__17821\,
            lcout => OPEN,
            ltout => \Lab_UT.dispString.m49Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17874\,
            in1 => \N__21171\,
            in2 => \N__17868\,
            in3 => \N__17964\,
            lcout => \Lab_UT.dispString.N_128_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNINM4L3_2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__25598\,
            in1 => \N__21327\,
            in2 => \_gnd_net_\,
            in3 => \N__17846\,
            lcout => \Lab_UT.sec1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26722\,
            lcout => \Lab_UT.di_ASones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26154\,
            ce => \N__18014\,
            sr => \N__25810\
        );

    \Lab_UT.didp.regrce1.q_esr_RNIH4M54_0_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21303\,
            in1 => \N__17939\,
            in2 => \_gnd_net_\,
            in3 => \N__17999\,
            lcout => \Lab_UT.sec2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_0_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21802\,
            lcout => \Lab_UT.di_ASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26154\,
            ce => \N__18014\,
            sr => \N__25810\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__21263\,
            in1 => \N__25520\,
            in2 => \N__22524\,
            in3 => \N__17936\,
            lcout => \Lab_UT.didp.countrce1.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25879\,
            in2 => \_gnd_net_\,
            in3 => \N__18039\,
            lcout => \Lab_UT.didp.regrce1.LdASones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_11_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__17935\,
            in1 => \N__17998\,
            in2 => \N__17982\,
            in3 => \N__17970\,
            lcout => \Lab_UT.dispString.m49Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__17937\,
            in1 => \N__22521\,
            in2 => \_gnd_net_\,
            in3 => \N__21804\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce1.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce1.q_0_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__21986\,
            in1 => \N__22644\,
            in2 => \N__17958\,
            in3 => \N__17938\,
            lcout => \Lab_UT.di_Sones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24536\,
            in1 => \N__22766\,
            in2 => \N__23162\,
            in3 => \N__18225\,
            lcout => \Lab_UT.LdMtens\,
            ltout => \Lab_UT.LdMtens_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNIDJKH1_3_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17913\,
            in3 => \N__22334\,
            lcout => \Lab_UT.didp.un1_dicLdMtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__18395\,
            in1 => \N__21803\,
            in2 => \_gnd_net_\,
            in3 => \N__21959\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000001"
        )
    port map (
            in0 => \N__22184\,
            in1 => \N__18399\,
            in2 => \N__18414\,
            in3 => \N__22335\,
            lcout => \Lab_UT.di_Mtens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__25519\,
            in1 => \N__22267\,
            in2 => \N__18406\,
            in3 => \N__21960\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce4.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce4.q_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__22185\,
            in1 => \N__22268\,
            in2 => \N__18375\,
            in3 => \N__18359\,
            lcout => \Lab_UT.di_Mtens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010001"
        )
    port map (
            in0 => \N__24368\,
            in1 => \N__23984\,
            in2 => \N__19527\,
            in3 => \N__19666\,
            lcout => \Lab_UT.dictrl.N_1462_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJ_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18271\,
            in2 => \_gnd_net_\,
            in3 => \N__19665\,
            lcout => \Lab_UT.dictrl.state_0_0_rep1_esr_RNICSUJZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__18233\,
            in1 => \N__24485\,
            in2 => \N__22113\,
            in3 => \N__18171\,
            lcout => \Lab_UT.didp.ceZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26133\,
            ce => 'H',
            sr => \N__25814\
        );

    \Lab_UT.didp.ce_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__22143\,
            in1 => \N__22108\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.ceZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26133\,
            ce => 'H',
            sr => \N__25814\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_8_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__19203\,
            in1 => \N__18158\,
            in2 => \_gnd_net_\,
            in3 => \N__19049\,
            lcout => \Lab_UT.dictrl.g1_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_6_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18159\,
            in1 => \N__21786\,
            in2 => \_gnd_net_\,
            in3 => \N__19712\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g0_i_a4_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNO_4_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__19204\,
            in1 => \N__19059\,
            in2 => \N__19053\,
            in3 => \N__19050\,
            lcout => \Lab_UT.dictrl.N_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_3_rep2_esr_RNITVU03_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__18948\,
            in1 => \N__19961\,
            in2 => \N__18934\,
            in3 => \N__19711\,
            lcout => \Lab_UT.dictrl.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m22_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000100"
        )
    port map (
            in0 => \N__18569\,
            in1 => \N__20191\,
            in2 => \N__18771\,
            in3 => \N__18651\,
            lcout => \Lab_UT.dictrl.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_8_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__18570\,
            in1 => \N__20192\,
            in2 => \_gnd_net_\,
            in3 => \N__19960\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_97_mux_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_5_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101111"
        )
    port map (
            in0 => \N__18471\,
            in1 => \N__19833\,
            in2 => \N__18459\,
            in3 => \N__19716\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1102_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_3_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__18456\,
            in1 => \N__18444\,
            in2 => \N__18435\,
            in3 => \N__24039\,
            lcout => \Lab_UT.dictrl.N_1460_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__18431\,
            in1 => \N__24146\,
            in2 => \N__19458\,
            in3 => \N__19328\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1106_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIDHBB9_0_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__24544\,
            in1 => \N__20532\,
            in2 => \N__18417\,
            in3 => \N__24277\,
            lcout => \Lab_UT.dictrl.g1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g1_1_0_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20070\,
            in1 => \N__20395\,
            in2 => \_gnd_net_\,
            in3 => \N__19448\,
            lcout => \Lab_UT.dictrl.g1_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.m28_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__19449\,
            in1 => \_gnd_net_\,
            in2 => \N__20407\,
            in3 => \N__20071\,
            lcout => \Lab_UT.dictrl.N_59\,
            ltout => \Lab_UT.dictrl.N_59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5_0_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011000000"
        )
    port map (
            in0 => \N__19351\,
            in1 => \N__24145\,
            in2 => \N__19335\,
            in3 => \N__19326\,
            lcout => \Lab_UT.dictrl.state_0_0_rep2_esr_RNI3PHI5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_2_rep2_esr_RNICN0J_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19327\,
            in2 => \_gnd_net_\,
            in3 => \N__19832\,
            lcout => \Lab_UT.dictrl.g2_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_50_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20322\,
            in1 => \N__20086\,
            in2 => \N__20223\,
            in3 => \N__20594\,
            lcout => \Lab_UT.dictrl.N_40_5\,
            ltout => \Lab_UT.dictrl.N_40_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_6_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__23966\,
            in1 => \N__19528\,
            in2 => \N__19230\,
            in3 => \N__19714\,
            lcout => \Lab_UT.dictrl.N_1462_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_43_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__20321\,
            in1 => \N__20082\,
            in2 => \N__20222\,
            in3 => \N__20592\,
            lcout => \Lab_UT.dictrl.N_40_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_26_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20593\,
            in1 => \N__20207\,
            in2 => \N__20093\,
            in3 => \N__20320\,
            lcout => \Lab_UT.dictrl.N_40_2\,
            ltout => \Lab_UT.dictrl.N_40_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_6_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000101"
        )
    port map (
            in0 => \N__19713\,
            in1 => \N__19534\,
            in2 => \N__19215\,
            in3 => \N__23965\,
            lcout => \Lab_UT.dictrl.N_1462_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.g0_64_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__20591\,
            in1 => \N__20206\,
            in2 => \N__20092\,
            in3 => \N__20319\,
            lcout => \Lab_UT.dictrl.N_40_7\,
            ltout => \Lab_UT.dictrl.N_40_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.next_state_RNIIKGR3_1_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000101"
        )
    port map (
            in0 => \N__19715\,
            in1 => \N__19533\,
            in2 => \N__20526\,
            in3 => \N__23967\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1462_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNIQRMCB_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__23968\,
            in1 => \N__20523\,
            in2 => \N__20517\,
            in3 => \N__20514\,
            lcout => \Lab_UT.dictrl.N_1460_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_RNO_9_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__20504\,
            in1 => \N__20408\,
            in2 => \N__20076\,
            in3 => \N__20318\,
            lcout => \Lab_UT.dictrl.g0_i_m2_0_a7_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_8_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__20219\,
            in1 => \N__20049\,
            in2 => \_gnd_net_\,
            in3 => \N__19962\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_97_mux_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_5_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011101111"
        )
    port map (
            in0 => \N__19863\,
            in1 => \N__19843\,
            in2 => \N__19740\,
            in3 => \N__19734\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1102_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__19572\,
            in1 => \N__19557\,
            in2 => \N__19551\,
            in3 => \N__24055\,
            lcout => \Lab_UT.dictrl.N_1460_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__19548\,
            in1 => \N__24546\,
            in2 => \N__19542\,
            in3 => \N__24063\,
            lcout => \Lab_UT.dictrl.g0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_user_5_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20972\,
            in1 => \N__20930\,
            in2 => \N__21012\,
            in3 => \N__21037\,
            lcout => \uu2.w_addr_userZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__20844\
        );

    \uu2.w_addr_user_4_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__20929\,
            in1 => \N__20999\,
            in2 => \_gnd_net_\,
            in3 => \N__20971\,
            lcout => \uu2.w_addr_userZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__20844\
        );

    \uu2.w_addr_user_6_LC_11_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__20973\,
            in1 => \N__20931\,
            in2 => \N__20907\,
            in3 => \N__20871\,
            lcout => \uu2.w_addr_userZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_user_5C_net\,
            ce => 'H',
            sr => \N__20844\
        );

    \uu2.w_addr_displaying_RNIMNI42_3_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__25102\,
            in1 => \N__20759\,
            in2 => \N__20685\,
            in3 => \N__24843\,
            lcout => OPEN,
            ltout => \uu2.w_addr_displaying_RNIMNI42Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNI9SFF4_1_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20691\,
            in2 => \N__20802\,
            in3 => \N__21087\,
            lcout => \uu2.N_397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIR9TO_1_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__20790\,
            in1 => \N__25170\,
            in2 => \_gnd_net_\,
            in3 => \N__20758\,
            lcout => \uu2.bitmap_pmux_sn_N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNILMVP_180_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20674\,
            in1 => \N__21081\,
            in2 => \_gnd_net_\,
            in3 => \N__24900\,
            lcout => \uu2.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIBP86_0_2_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20675\,
            in2 => \_gnd_net_\,
            in3 => \N__20634\,
            lcout => \uu2.w_addr_displaying_fast_RNIBP86_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_314_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110101"
        )
    port map (
            in0 => \N__21421\,
            in1 => \N__21529\,
            in2 => \N__21578\,
            in3 => \N__21475\,
            lcout => \uu2.bitmapZ0Z_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__25776\
        );

    \uu2.bitmap_218_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000011101"
        )
    port map (
            in0 => \N__21474\,
            in1 => \N__21571\,
            in2 => \N__21531\,
            in3 => \N__21420\,
            lcout => \uu2.bitmapZ0Z_218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__25776\
        );

    \uu2.bitmap_90_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100001101"
        )
    port map (
            in0 => \N__21422\,
            in1 => \N__21530\,
            in2 => \N__21579\,
            in3 => \N__21476\,
            lcout => \uu2.bitmapZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_314C_net\,
            ce => 'H',
            sr => \N__25776\
        );

    \uu2.bitmap_RNIC7SJ_90_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21159\,
            in1 => \N__21153\,
            in2 => \_gnd_net_\,
            in3 => \N__21133\,
            lcout => \uu2.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNIE7RK_58_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__21080\,
            in1 => \N__24892\,
            in2 => \_gnd_net_\,
            in3 => \N__21384\,
            lcout => OPEN,
            ltout => \uu2.bitmap_RNIE7RKZ0Z_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_RNIOQVH1_7_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21134\,
            in1 => \_gnd_net_\,
            in2 => \N__21090\,
            in3 => \N__21063\,
            lcout => \uu2.w_addr_displaying_fast_RNIOQVH1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNI020Q_186_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21057\,
            in1 => \N__24891\,
            in2 => \_gnd_net_\,
            in3 => \N__21079\,
            lcout => \uu2.bitmap_RNI020QZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_87_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100101111111"
        )
    port map (
            in0 => \N__24621\,
            in1 => \N__24687\,
            in2 => \N__24730\,
            in3 => \N__24786\,
            lcout => \uu2.bitmapZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__25773\
        );

    \uu2.bitmap_308_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000011101"
        )
    port map (
            in0 => \N__24784\,
            in1 => \N__24718\,
            in2 => \N__24694\,
            in3 => \N__24619\,
            lcout => \uu2.bitmapZ0Z_308\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__25773\
        );

    \uu2.bitmap_186_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100111100"
        )
    port map (
            in0 => \N__21428\,
            in1 => \N__21470\,
            in2 => \N__21525\,
            in3 => \N__21569\,
            lcout => \uu2.bitmapZ0Z_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__25773\
        );

    \uu2.bitmap_58_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011011011101111"
        )
    port map (
            in0 => \N__21570\,
            in1 => \N__21517\,
            in2 => \N__21477\,
            in3 => \N__21429\,
            lcout => \uu2.bitmapZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__25773\
        );

    \uu2.bitmap_52_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001111011111101"
        )
    port map (
            in0 => \N__24785\,
            in1 => \N__24719\,
            in2 => \N__24695\,
            in3 => \N__24620\,
            lcout => \uu2.bitmapZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_87C_net\,
            ce => 'H',
            sr => \N__25773\
        );

    \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25554\,
            in1 => \N__25588\,
            in2 => \N__25226\,
            in3 => \N__25297\,
            lcout => \Lab_UT.didp.un24_ce_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_0_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__25260\,
            in1 => \N__21806\,
            in2 => \_gnd_net_\,
            in3 => \N__25555\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_0_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__25556\,
            in1 => \N__25330\,
            in2 => \N__21378\,
            in3 => \N__25362\,
            lcout => \Lab_UT.di_Stens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNIJI4L3_0_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21345\,
            in1 => \N__25553\,
            in2 => \_gnd_net_\,
            in3 => \N__21374\,
            lcout => \Lab_UT.sec1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce2.q_esr_RNILK4L3_1_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21221\,
            in1 => \N__21346\,
            in2 => \_gnd_net_\,
            in3 => \N__25296\,
            lcout => \Lab_UT.sec1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__21264\,
            in1 => \N__21220\,
            in2 => \N__25302\,
            in3 => \N__21194\,
            lcout => \Lab_UT.dispString.m49Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.regrce3.q_esr_1_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25524\,
            lcout => \Lab_UT.di_AMones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26171\,
            ce => \N__21828\,
            sr => \N__25816\
        );

    \Lab_UT.didp.regrce3.q_esr_2_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26739\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.di_AMones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26171\,
            ce => \N__21828\,
            sr => \N__25816\
        );

    \Lab_UT.didp.regrce3.q_esr_3_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26424\,
            lcout => \Lab_UT.di_AMones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26171\,
            ce => \N__21828\,
            sr => \N__25816\
        );

    \Lab_UT.didp.countrce3.q_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001001"
        )
    port map (
            in0 => \N__22320\,
            in1 => \N__21666\,
            in2 => \N__26259\,
            in3 => \N__26458\,
            lcout => \Lab_UT.di_Mones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26164\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_0_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__26457\,
            in1 => \N__21807\,
            in2 => \_gnd_net_\,
            in3 => \N__26531\,
            lcout => \Lab_UT.didp.countrce3.q_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI4EIS1_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22319\,
            in2 => \_gnd_net_\,
            in3 => \N__26455\,
            lcout => \Lab_UT.didp.un1_dicLdMones_0\,
            ltout => \Lab_UT.didp.un1_dicLdMones_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000000010"
        )
    port map (
            in0 => \N__21657\,
            in1 => \N__26256\,
            in2 => \N__21660\,
            in3 => \N__26566\,
            lcout => \Lab_UT.di_Mones_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26164\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_1_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__26530\,
            in1 => \N__26456\,
            in2 => \N__26573\,
            in3 => \N__25481\,
            lcout => \Lab_UT.didp.countrce3.q_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dispString.m49_2_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__21640\,
            in1 => \N__26562\,
            in2 => \N__21613\,
            in3 => \N__26482\,
            lcout => \Lab_UT.dispString.m49Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22147\,
            in1 => \_gnd_net_\,
            in2 => \N__22111\,
            in3 => \N__22302\,
            lcout => \Lab_UT.didp.resetZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.ce_3_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__25184\,
            in1 => \N__22095\,
            in2 => \N__22305\,
            in3 => \N__22148\,
            lcout => \Lab_UT.didp.ceZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.reset_2_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22149\,
            in1 => \N__25185\,
            in2 => \N__22112\,
            in3 => \N__22304\,
            lcout => \Lab_UT.didp.resetZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.ce_2_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22303\,
            in1 => \N__22094\,
            in2 => \_gnd_net_\,
            in3 => \N__22145\,
            lcout => \Lab_UT.didp.ceZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__22144\,
            in1 => \N__25183\,
            in2 => \N__22109\,
            in3 => \N__22298\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.ce_12_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.reset_3_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__21882\,
            in1 => \N__22280\,
            in2 => \N__22221\,
            in3 => \N__22218\,
            lcout => \Lab_UT.didp.resetZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.reset_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__22146\,
            in1 => \_gnd_net_\,
            in2 => \N__22110\,
            in3 => \_gnd_net_\,
            lcout => \Lab_UT.didp.resetZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26155\,
            ce => 'H',
            sr => \N__25811\
        );

    \Lab_UT.didp.reset_RNO_0_3_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__21972\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21918\,
            lcout => \Lab_UT.didp.reset_12_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.ce_RNI5U3I_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21876\,
            in2 => \_gnd_net_\,
            in3 => \N__21864\,
            lcout => \Lab_UT.didp.un1_dicLdStens_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_2_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__23132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23958\,
            lcout => \Lab_UT.dictrl.g2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24535\,
            in1 => \N__22765\,
            in2 => \N__23160\,
            in3 => \N__24308\,
            lcout => \Lab_UT.LdMones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__22854\,
            in1 => \N__22689\,
            in2 => \N__22674\,
            in3 => \N__22980\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_state_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__23204\,
            in1 => \N__22567\,
            in2 => \N__22662\,
            in3 => \N__22605\,
            lcout => \Lab_UT.LdSones_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26143\,
            ce => \N__22486\,
            sr => \N__25815\
        );

    \Lab_UT.dictrl.state_ret_6_esr_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23001\,
            in1 => \N__22604\,
            in2 => \N__22569\,
            in3 => \N__23203\,
            lcout => \Lab_UT.LdStens\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26143\,
            ce => \N__22486\,
            sr => \N__25815\
        );

    \Lab_UT.didp.ce_RNI51AM_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22659\,
            in2 => \_gnd_net_\,
            in3 => \N__22650\,
            lcout => \Lab_UT.didp.un1_dicLdSones_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__23172\,
            in1 => \N__22603\,
            in2 => \N__22568\,
            in3 => \N__23202\,
            lcout => \Lab_UT.LdSones\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26143\,
            ce => \N__22486\,
            sr => \N__25815\
        );

    \Lab_UT.dictrl.state_0_esr_RNIP2CG_0_1_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23133\,
            in2 => \_gnd_net_\,
            in3 => \N__23827\,
            lcout => \Lab_UT.dictrl.g2_5\,
            ltout => \Lab_UT.dictrl.g2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_2_ess_RNIRP7EL_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__22418\,
            in1 => \N__22967\,
            in2 => \N__22383\,
            in3 => \N__22370\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.next_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_12_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__23229\,
            in1 => \N__23220\,
            in2 => \N__23211\,
            in3 => \N__23208\,
            lcout => \Lab_UT.dictrl.un1_next_state66_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_2_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__23828\,
            in1 => \_gnd_net_\,
            in2 => \N__23161\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__23715\,
            in1 => \N__22966\,
            in2 => \N__23175\,
            in3 => \N__22833\,
            lcout => \Lab_UT.dictrl.next_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_2_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__23137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23829\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.g2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__23013\,
            in1 => \N__24351\,
            in2 => \N__23004\,
            in3 => \N__22973\,
            lcout => \Lab_UT.dictrl.next_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_3_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__24306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24545\,
            lcout => OPEN,
            ltout => \Lab_UT.dictrl.N_1105_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_1_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000000"
        )
    port map (
            in0 => \N__22992\,
            in1 => \N__24108\,
            in2 => \N__22983\,
            in3 => \N__22972\,
            lcout => \Lab_UT.dictrl.N_79_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_8_ess_RNO_1_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__24584\,
            in1 => \N__22866\,
            in2 => \N__24323\,
            in3 => \N__24543\,
            lcout => \Lab_UT.dictrl.g1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110000000"
        )
    port map (
            in0 => \N__22845\,
            in1 => \N__24309\,
            in2 => \N__24554\,
            in3 => \N__24582\,
            lcout => \Lab_UT.dictrl.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_6_esr_RNO_1_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__24583\,
            in1 => \N__24307\,
            in2 => \N__24553\,
            in3 => \N__24372\,
            lcout => \Lab_UT.dictrl.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_3_ess_RNO_4_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__24341\,
            in1 => \N__24305\,
            in2 => \N__24162\,
            in3 => \N__24147\,
            lcout => \Lab_UT.dictrl.N_1106_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_ret_4_esr_RNO_3_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001010"
        )
    port map (
            in0 => \N__24099\,
            in1 => \N__24087\,
            in2 => \N__24075\,
            in3 => \N__24056\,
            lcout => \Lab_UT.dictrl.N_1460_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.mem0.ram512X8_inst_RNO_7_LC_12_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__23704\,
            in1 => \N__23616\,
            in2 => \N__23544\,
            in3 => \N__25171\,
            lcout => \uu2.mem0.w_addr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_0_LC_12_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23327\,
            in2 => \_gnd_net_\,
            in3 => \N__25030\,
            lcout => \uu2.w_addr_displayingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__25780\
        );

    \uu2.w_addr_displaying_nesr_RNIA8E42_5_LC_12_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23486\,
            in1 => \N__23417\,
            in2 => \N__23342\,
            in3 => \N__23295\,
            lcout => \uu2.N_14_i\,
            ltout => \uu2.N_14_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_RNI6OAF2_6_LC_12_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23259\,
            in3 => \N__24936\,
            lcout => \uu2.N_15_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_fast_0_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__25031\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24824\,
            lcout => \uu2.w_addr_displaying_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__25780\
        );

    \uu2.w_addr_displaying_RNO_0_6_LC_12_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25172\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25103\,
            lcout => OPEN,
            ltout => \uu2.N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.w_addr_displaying_6_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101100111001100"
        )
    port map (
            in0 => \N__25032\,
            in1 => \N__24937\,
            in2 => \N__24966\,
            in3 => \N__24963\,
            lcout => \uu2.w_addr_displayingZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.w_addr_displaying_0C_net\,
            ce => 'H',
            sr => \N__25780\
        );

    \uu2.bitmap_212_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000101"
        )
    port map (
            in0 => \N__24632\,
            in1 => \N__24692\,
            in2 => \N__24795\,
            in3 => \N__24740\,
            lcout => \uu2.bitmapZ0Z_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_212C_net\,
            ce => 'H',
            sr => \N__25779\
        );

    \uu2.bitmap_180_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100111100"
        )
    port map (
            in0 => \N__24631\,
            in1 => \N__24691\,
            in2 => \N__24794\,
            in3 => \N__24739\,
            lcout => \uu2.bitmapZ0Z_180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_212C_net\,
            ce => 'H',
            sr => \N__25779\
        );

    \uu2.bitmap_RNIB3QK_52_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__24893\,
            in1 => \N__24855\,
            in2 => \_gnd_net_\,
            in3 => \N__24849\,
            lcout => \uu2.N_194\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_RNISLTD_84_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24837\,
            in1 => \N__24594\,
            in2 => \_gnd_net_\,
            in3 => \N__24820\,
            lcout => \uu2.N_197\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uu2.bitmap_84_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000011011"
        )
    port map (
            in0 => \N__24787\,
            in1 => \N__24723\,
            in2 => \N__24696\,
            in3 => \N__24622\,
            lcout => \uu2.bitmapZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuu2.bitmap_84C_net\,
            ce => 'H',
            sr => \N__25777\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_3_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__25298\,
            in1 => \N__25586\,
            in2 => \_gnd_net_\,
            in3 => \N__25557\,
            lcout => \Lab_UT.didp.countrce2.un20_qPone\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_1_2_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25558\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25299\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_2_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001011010"
        )
    port map (
            in0 => \N__25589\,
            in1 => \N__26738\,
            in2 => \N__25605\,
            in3 => \N__25264\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_2_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__25587\,
            in1 => \N__25331\,
            in2 => \N__25602\,
            in3 => \N__25364\,
            lcout => \Lab_UT.di_Stens_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_3_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000100"
        )
    port map (
            in0 => \N__25365\,
            in1 => \N__25191\,
            in2 => \N__25335\,
            in3 => \N__25221\,
            lcout => \Lab_UT.di_Stens_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_1_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__25559\,
            in1 => \N__25493\,
            in2 => \N__25266\,
            in3 => \N__25300\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce2.q_5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111000"
        )
    port map (
            in0 => \N__25301\,
            in1 => \N__25363\,
            in2 => \N__25338\,
            in3 => \N__25329\,
            lcout => \Lab_UT.di_Stens_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce2.q_RNO_0_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__25272\,
            in1 => \N__26423\,
            in2 => \N__25265\,
            in3 => \N__25220\,
            lcout => \Lab_UT.didp.countrce2.q_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__26570\,
            in1 => \N__26527\,
            in2 => \N__26497\,
            in3 => \N__26228\,
            lcout => \Lab_UT.didp.countrce3.ce_12_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_2_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__26528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26572\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un13_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_2_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__26492\,
            in1 => \N__26459\,
            in2 => \N__26742\,
            in3 => \N__26731\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_2_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__26257\,
            in1 => \N__26267\,
            in2 => \N__26580\,
            in3 => \N__26493\,
            lcout => \Lab_UT.di_Mones_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_1_3_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__26571\,
            in1 => \N__26529\,
            in2 => \N__26498\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.un20_qPone_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_RNO_0_3_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111000010010"
        )
    port map (
            in0 => \N__26229\,
            in1 => \N__26460\,
            in2 => \N__26427\,
            in3 => \N__26388\,
            lcout => OPEN,
            ltout => \Lab_UT.didp.countrce3.q_5_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.didp.countrce3.q_3_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__26268\,
            in1 => \N__26258\,
            in2 => \N__26238\,
            in3 => \N__26230\,
            lcout => \Lab_UT.di_Mones_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__26172\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Lab_UT.dictrl.state_0_1_rep2_esr_ctle_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25918\,
            in2 => \_gnd_net_\,
            in3 => \N__25875\,
            lcout => bu_rx_data_rdy_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
