// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 19 2019 07:46:31

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__18473;
    wire N__18472;
    wire N__18471;
    wire N__18464;
    wire N__18463;
    wire N__18462;
    wire N__18455;
    wire N__18454;
    wire N__18453;
    wire N__18446;
    wire N__18445;
    wire N__18444;
    wire N__18437;
    wire N__18436;
    wire N__18435;
    wire N__18428;
    wire N__18427;
    wire N__18426;
    wire N__18419;
    wire N__18418;
    wire N__18417;
    wire N__18410;
    wire N__18409;
    wire N__18408;
    wire N__18401;
    wire N__18400;
    wire N__18399;
    wire N__18392;
    wire N__18391;
    wire N__18390;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18363;
    wire N__18358;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18352;
    wire N__18349;
    wire N__18342;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18319;
    wire N__18318;
    wire N__18317;
    wire N__18316;
    wire N__18309;
    wire N__18306;
    wire N__18305;
    wire N__18304;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18290;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18261;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18253;
    wire N__18250;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18222;
    wire N__18219;
    wire N__18218;
    wire N__18217;
    wire N__18216;
    wire N__18215;
    wire N__18212;
    wire N__18207;
    wire N__18204;
    wire N__18199;
    wire N__18190;
    wire N__18189;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18182;
    wire N__18181;
    wire N__18180;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18162;
    wire N__18159;
    wire N__18148;
    wire N__18147;
    wire N__18146;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18134;
    wire N__18127;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18119;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18097;
    wire N__18096;
    wire N__18095;
    wire N__18094;
    wire N__18093;
    wire N__18092;
    wire N__18091;
    wire N__18090;
    wire N__18089;
    wire N__18088;
    wire N__18087;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18077;
    wire N__18076;
    wire N__18075;
    wire N__18074;
    wire N__18073;
    wire N__18072;
    wire N__18071;
    wire N__18070;
    wire N__18069;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18064;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18045;
    wire N__18044;
    wire N__18043;
    wire N__18042;
    wire N__18041;
    wire N__18040;
    wire N__18039;
    wire N__18038;
    wire N__18037;
    wire N__18036;
    wire N__18035;
    wire N__18034;
    wire N__18033;
    wire N__18032;
    wire N__18031;
    wire N__18030;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18025;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18021;
    wire N__18020;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17853;
    wire N__17852;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17833;
    wire N__17832;
    wire N__17831;
    wire N__17830;
    wire N__17829;
    wire N__17828;
    wire N__17827;
    wire N__17826;
    wire N__17825;
    wire N__17824;
    wire N__17823;
    wire N__17822;
    wire N__17821;
    wire N__17820;
    wire N__17819;
    wire N__17818;
    wire N__17817;
    wire N__17816;
    wire N__17815;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17810;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17789;
    wire N__17788;
    wire N__17787;
    wire N__17786;
    wire N__17785;
    wire N__17784;
    wire N__17783;
    wire N__17782;
    wire N__17781;
    wire N__17780;
    wire N__17779;
    wire N__17778;
    wire N__17777;
    wire N__17776;
    wire N__17773;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17646;
    wire N__17645;
    wire N__17644;
    wire N__17643;
    wire N__17642;
    wire N__17639;
    wire N__17638;
    wire N__17637;
    wire N__17632;
    wire N__17625;
    wire N__17622;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17603;
    wire N__17598;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17580;
    wire N__17579;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17559;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17551;
    wire N__17550;
    wire N__17549;
    wire N__17548;
    wire N__17547;
    wire N__17546;
    wire N__17545;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17528;
    wire N__17523;
    wire N__17520;
    wire N__17509;
    wire N__17494;
    wire N__17493;
    wire N__17492;
    wire N__17489;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17475;
    wire N__17474;
    wire N__17473;
    wire N__17472;
    wire N__17471;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17457;
    wire N__17454;
    wire N__17453;
    wire N__17452;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17434;
    wire N__17431;
    wire N__17426;
    wire N__17421;
    wire N__17416;
    wire N__17409;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17388;
    wire N__17387;
    wire N__17386;
    wire N__17385;
    wire N__17382;
    wire N__17377;
    wire N__17372;
    wire N__17365;
    wire N__17364;
    wire N__17363;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17351;
    wire N__17348;
    wire N__17341;
    wire N__17340;
    wire N__17337;
    wire N__17336;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17303;
    wire N__17296;
    wire N__17293;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17254;
    wire N__17253;
    wire N__17252;
    wire N__17251;
    wire N__17250;
    wire N__17249;
    wire N__17248;
    wire N__17243;
    wire N__17240;
    wire N__17231;
    wire N__17230;
    wire N__17227;
    wire N__17222;
    wire N__17221;
    wire N__17220;
    wire N__17219;
    wire N__17216;
    wire N__17215;
    wire N__17214;
    wire N__17209;
    wire N__17204;
    wire N__17203;
    wire N__17202;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17177;
    wire N__17164;
    wire N__17163;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17146;
    wire N__17145;
    wire N__17144;
    wire N__17143;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17127;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17080;
    wire N__17079;
    wire N__17078;
    wire N__17075;
    wire N__17074;
    wire N__17073;
    wire N__17072;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17053;
    wire N__17044;
    wire N__17043;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17020;
    wire N__17019;
    wire N__17018;
    wire N__17017;
    wire N__17016;
    wire N__17015;
    wire N__17010;
    wire N__17009;
    wire N__17008;
    wire N__17005;
    wire N__17004;
    wire N__17001;
    wire N__16996;
    wire N__16993;
    wire N__16984;
    wire N__16981;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16963;
    wire N__16962;
    wire N__16961;
    wire N__16958;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16942;
    wire N__16941;
    wire N__16940;
    wire N__16933;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16918;
    wire N__16915;
    wire N__16914;
    wire N__16913;
    wire N__16912;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16901;
    wire N__16898;
    wire N__16897;
    wire N__16896;
    wire N__16893;
    wire N__16888;
    wire N__16887;
    wire N__16886;
    wire N__16881;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16860;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16844;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16810;
    wire N__16807;
    wire N__16806;
    wire N__16805;
    wire N__16802;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16786;
    wire N__16785;
    wire N__16784;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16773;
    wire N__16772;
    wire N__16769;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16759;
    wire N__16756;
    wire N__16755;
    wire N__16752;
    wire N__16747;
    wire N__16740;
    wire N__16737;
    wire N__16734;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16710;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16698;
    wire N__16697;
    wire N__16696;
    wire N__16687;
    wire N__16684;
    wire N__16681;
    wire N__16680;
    wire N__16675;
    wire N__16672;
    wire N__16671;
    wire N__16668;
    wire N__16667;
    wire N__16664;
    wire N__16663;
    wire N__16658;
    wire N__16653;
    wire N__16648;
    wire N__16647;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16636;
    wire N__16633;
    wire N__16626;
    wire N__16619;
    wire N__16618;
    wire N__16617;
    wire N__16614;
    wire N__16613;
    wire N__16612;
    wire N__16611;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16597;
    wire N__16590;
    wire N__16587;
    wire N__16576;
    wire N__16575;
    wire N__16574;
    wire N__16573;
    wire N__16570;
    wire N__16569;
    wire N__16568;
    wire N__16567;
    wire N__16566;
    wire N__16559;
    wire N__16558;
    wire N__16555;
    wire N__16554;
    wire N__16553;
    wire N__16550;
    wire N__16549;
    wire N__16548;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16527;
    wire N__16520;
    wire N__16515;
    wire N__16504;
    wire N__16503;
    wire N__16502;
    wire N__16501;
    wire N__16500;
    wire N__16499;
    wire N__16496;
    wire N__16493;
    wire N__16490;
    wire N__16483;
    wire N__16482;
    wire N__16481;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16462;
    wire N__16461;
    wire N__16460;
    wire N__16459;
    wire N__16454;
    wire N__16451;
    wire N__16444;
    wire N__16441;
    wire N__16434;
    wire N__16431;
    wire N__16420;
    wire N__16419;
    wire N__16418;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16410;
    wire N__16409;
    wire N__16408;
    wire N__16407;
    wire N__16406;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16367;
    wire N__16362;
    wire N__16359;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16341;
    wire N__16340;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16328;
    wire N__16321;
    wire N__16320;
    wire N__16319;
    wire N__16314;
    wire N__16313;
    wire N__16312;
    wire N__16311;
    wire N__16310;
    wire N__16309;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16297;
    wire N__16296;
    wire N__16293;
    wire N__16292;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16280;
    wire N__16275;
    wire N__16262;
    wire N__16255;
    wire N__16252;
    wire N__16251;
    wire N__16250;
    wire N__16247;
    wire N__16244;
    wire N__16243;
    wire N__16240;
    wire N__16239;
    wire N__16236;
    wire N__16231;
    wire N__16230;
    wire N__16229;
    wire N__16226;
    wire N__16225;
    wire N__16224;
    wire N__16223;
    wire N__16222;
    wire N__16221;
    wire N__16220;
    wire N__16217;
    wire N__16212;
    wire N__16207;
    wire N__16204;
    wire N__16191;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16172;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16164;
    wire N__16163;
    wire N__16162;
    wire N__16161;
    wire N__16160;
    wire N__16157;
    wire N__16156;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16138;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16126;
    wire N__16121;
    wire N__16114;
    wire N__16103;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16071;
    wire N__16070;
    wire N__16069;
    wire N__16064;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16049;
    wire N__16048;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16032;
    wire N__16031;
    wire N__16028;
    wire N__16027;
    wire N__16026;
    wire N__16025;
    wire N__16022;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__15999;
    wire N__15996;
    wire N__15985;
    wire N__15984;
    wire N__15983;
    wire N__15982;
    wire N__15981;
    wire N__15980;
    wire N__15979;
    wire N__15978;
    wire N__15977;
    wire N__15974;
    wire N__15969;
    wire N__15968;
    wire N__15963;
    wire N__15954;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15946;
    wire N__15945;
    wire N__15944;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15916;
    wire N__15909;
    wire N__15898;
    wire N__15895;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15880;
    wire N__15879;
    wire N__15876;
    wire N__15875;
    wire N__15872;
    wire N__15867;
    wire N__15864;
    wire N__15859;
    wire N__15856;
    wire N__15855;
    wire N__15852;
    wire N__15851;
    wire N__15848;
    wire N__15847;
    wire N__15844;
    wire N__15837;
    wire N__15832;
    wire N__15829;
    wire N__15826;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15820;
    wire N__15819;
    wire N__15818;
    wire N__15815;
    wire N__15814;
    wire N__15813;
    wire N__15808;
    wire N__15803;
    wire N__15796;
    wire N__15795;
    wire N__15794;
    wire N__15791;
    wire N__15788;
    wire N__15785;
    wire N__15782;
    wire N__15779;
    wire N__15778;
    wire N__15775;
    wire N__15774;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15762;
    wire N__15753;
    wire N__15750;
    wire N__15739;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15731;
    wire N__15730;
    wire N__15729;
    wire N__15728;
    wire N__15727;
    wire N__15726;
    wire N__15721;
    wire N__15716;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15702;
    wire N__15701;
    wire N__15700;
    wire N__15699;
    wire N__15698;
    wire N__15693;
    wire N__15692;
    wire N__15689;
    wire N__15686;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15651;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15639;
    wire N__15638;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15623;
    wire N__15622;
    wire N__15619;
    wire N__15614;
    wire N__15611;
    wire N__15604;
    wire N__15601;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15584;
    wire N__15581;
    wire N__15574;
    wire N__15571;
    wire N__15570;
    wire N__15569;
    wire N__15566;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15548;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15526;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15512;
    wire N__15511;
    wire N__15508;
    wire N__15503;
    wire N__15498;
    wire N__15495;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15489;
    wire N__15488;
    wire N__15487;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15469;
    wire N__15466;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15450;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15402;
    wire N__15401;
    wire N__15394;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15382;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15376;
    wire N__15375;
    wire N__15374;
    wire N__15373;
    wire N__15372;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15362;
    wire N__15359;
    wire N__15348;
    wire N__15341;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15325;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15311;
    wire N__15308;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15290;
    wire N__15289;
    wire N__15286;
    wire N__15283;
    wire N__15278;
    wire N__15271;
    wire N__15270;
    wire N__15269;
    wire N__15268;
    wire N__15267;
    wire N__15266;
    wire N__15265;
    wire N__15262;
    wire N__15251;
    wire N__15248;
    wire N__15247;
    wire N__15246;
    wire N__15245;
    wire N__15244;
    wire N__15243;
    wire N__15242;
    wire N__15241;
    wire N__15236;
    wire N__15233;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15207;
    wire N__15206;
    wire N__15199;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15178;
    wire N__15175;
    wire N__15174;
    wire N__15173;
    wire N__15172;
    wire N__15171;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15147;
    wire N__15142;
    wire N__15131;
    wire N__15126;
    wire N__15123;
    wire N__15122;
    wire N__15121;
    wire N__15120;
    wire N__15117;
    wire N__15112;
    wire N__15109;
    wire N__15100;
    wire N__15091;
    wire N__15088;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15067;
    wire N__15064;
    wire N__15061;
    wire N__15058;
    wire N__15057;
    wire N__15056;
    wire N__15055;
    wire N__15052;
    wire N__15045;
    wire N__15040;
    wire N__15037;
    wire N__15034;
    wire N__15031;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15011;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14991;
    wire N__14988;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14977;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14962;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14943;
    wire N__14942;
    wire N__14941;
    wire N__14938;
    wire N__14937;
    wire N__14936;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14920;
    wire N__14919;
    wire N__14918;
    wire N__14917;
    wire N__14916;
    wire N__14915;
    wire N__14914;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14896;
    wire N__14893;
    wire N__14888;
    wire N__14883;
    wire N__14882;
    wire N__14879;
    wire N__14874;
    wire N__14867;
    wire N__14862;
    wire N__14859;
    wire N__14852;
    wire N__14845;
    wire N__14842;
    wire N__14839;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14831;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14815;
    wire N__14814;
    wire N__14809;
    wire N__14806;
    wire N__14803;
    wire N__14800;
    wire N__14797;
    wire N__14794;
    wire N__14791;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14752;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14734;
    wire N__14733;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14710;
    wire N__14707;
    wire N__14706;
    wire N__14701;
    wire N__14700;
    wire N__14699;
    wire N__14696;
    wire N__14691;
    wire N__14686;
    wire N__14685;
    wire N__14680;
    wire N__14677;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14659;
    wire N__14656;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14631;
    wire N__14630;
    wire N__14629;
    wire N__14628;
    wire N__14627;
    wire N__14624;
    wire N__14619;
    wire N__14612;
    wire N__14605;
    wire N__14604;
    wire N__14603;
    wire N__14602;
    wire N__14601;
    wire N__14598;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14588;
    wire N__14587;
    wire N__14584;
    wire N__14583;
    wire N__14582;
    wire N__14577;
    wire N__14574;
    wire N__14567;
    wire N__14564;
    wire N__14559;
    wire N__14548;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14542;
    wire N__14541;
    wire N__14538;
    wire N__14533;
    wire N__14530;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14500;
    wire N__14497;
    wire N__14496;
    wire N__14493;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14470;
    wire N__14469;
    wire N__14466;
    wire N__14465;
    wire N__14462;
    wire N__14457;
    wire N__14454;
    wire N__14449;
    wire N__14448;
    wire N__14447;
    wire N__14446;
    wire N__14445;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14422;
    wire N__14419;
    wire N__14418;
    wire N__14417;
    wire N__14416;
    wire N__14413;
    wire N__14408;
    wire N__14405;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14389;
    wire N__14388;
    wire N__14387;
    wire N__14384;
    wire N__14383;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14365;
    wire N__14362;
    wire N__14359;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14323;
    wire N__14320;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14310;
    wire N__14309;
    wire N__14308;
    wire N__14305;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14287;
    wire N__14286;
    wire N__14283;
    wire N__14282;
    wire N__14281;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14263;
    wire N__14262;
    wire N__14261;
    wire N__14260;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14242;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14238;
    wire N__14237;
    wire N__14236;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14231;
    wire N__14230;
    wire N__14229;
    wire N__14228;
    wire N__14227;
    wire N__14226;
    wire N__14225;
    wire N__14224;
    wire N__14223;
    wire N__14218;
    wire N__14217;
    wire N__14216;
    wire N__14215;
    wire N__14212;
    wire N__14211;
    wire N__14210;
    wire N__14209;
    wire N__14208;
    wire N__14207;
    wire N__14204;
    wire N__14199;
    wire N__14192;
    wire N__14187;
    wire N__14180;
    wire N__14173;
    wire N__14166;
    wire N__14163;
    wire N__14156;
    wire N__14153;
    wire N__14146;
    wire N__14141;
    wire N__14138;
    wire N__14129;
    wire N__14126;
    wire N__14125;
    wire N__14124;
    wire N__14115;
    wire N__14104;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14086;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14074;
    wire N__14073;
    wire N__14072;
    wire N__14069;
    wire N__14064;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14040;
    wire N__14035;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14007;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13997;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13983;
    wire N__13982;
    wire N__13981;
    wire N__13980;
    wire N__13979;
    wire N__13978;
    wire N__13975;
    wire N__13970;
    wire N__13961;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13947;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13939;
    wire N__13938;
    wire N__13937;
    wire N__13934;
    wire N__13931;
    wire N__13920;
    wire N__13917;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13903;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13839;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13831;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13825;
    wire N__13824;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13804;
    wire N__13803;
    wire N__13802;
    wire N__13801;
    wire N__13800;
    wire N__13797;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13771;
    wire N__13764;
    wire N__13753;
    wire N__13752;
    wire N__13751;
    wire N__13748;
    wire N__13747;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13739;
    wire N__13738;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13712;
    wire N__13711;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13707;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13680;
    wire N__13671;
    wire N__13664;
    wire N__13655;
    wire N__13650;
    wire N__13641;
    wire N__13630;
    wire N__13629;
    wire N__13628;
    wire N__13627;
    wire N__13626;
    wire N__13625;
    wire N__13624;
    wire N__13623;
    wire N__13620;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13610;
    wire N__13609;
    wire N__13606;
    wire N__13595;
    wire N__13594;
    wire N__13593;
    wire N__13588;
    wire N__13585;
    wire N__13580;
    wire N__13579;
    wire N__13578;
    wire N__13577;
    wire N__13574;
    wire N__13569;
    wire N__13564;
    wire N__13561;
    wire N__13554;
    wire N__13551;
    wire N__13546;
    wire N__13541;
    wire N__13534;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13507;
    wire N__13506;
    wire N__13505;
    wire N__13504;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13500;
    wire N__13499;
    wire N__13498;
    wire N__13495;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13464;
    wire N__13459;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13429;
    wire N__13422;
    wire N__13411;
    wire N__13410;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13402;
    wire N__13399;
    wire N__13398;
    wire N__13397;
    wire N__13396;
    wire N__13395;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13384;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13353;
    wire N__13350;
    wire N__13343;
    wire N__13340;
    wire N__13335;
    wire N__13318;
    wire N__13317;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13304;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13290;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13260;
    wire N__13253;
    wire N__13248;
    wire N__13231;
    wire N__13230;
    wire N__13229;
    wire N__13226;
    wire N__13225;
    wire N__13220;
    wire N__13217;
    wire N__13216;
    wire N__13215;
    wire N__13214;
    wire N__13213;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13205;
    wire N__13204;
    wire N__13203;
    wire N__13202;
    wire N__13201;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13168;
    wire N__13163;
    wire N__13154;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13132;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13106;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13071;
    wire N__13070;
    wire N__13069;
    wire N__13066;
    wire N__13065;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13043;
    wire N__13038;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13029;
    wire N__13028;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13008;
    wire N__13003;
    wire N__12994;
    wire N__12979;
    wire N__12978;
    wire N__12975;
    wire N__12974;
    wire N__12973;
    wire N__12972;
    wire N__12971;
    wire N__12970;
    wire N__12969;
    wire N__12966;
    wire N__12959;
    wire N__12956;
    wire N__12955;
    wire N__12954;
    wire N__12949;
    wire N__12948;
    wire N__12947;
    wire N__12946;
    wire N__12945;
    wire N__12942;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12918;
    wire N__12915;
    wire N__12910;
    wire N__12895;
    wire N__12894;
    wire N__12893;
    wire N__12892;
    wire N__12889;
    wire N__12888;
    wire N__12885;
    wire N__12884;
    wire N__12883;
    wire N__12882;
    wire N__12881;
    wire N__12880;
    wire N__12879;
    wire N__12878;
    wire N__12877;
    wire N__12876;
    wire N__12875;
    wire N__12874;
    wire N__12869;
    wire N__12868;
    wire N__12867;
    wire N__12866;
    wire N__12865;
    wire N__12864;
    wire N__12861;
    wire N__12860;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12841;
    wire N__12840;
    wire N__12839;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12799;
    wire N__12794;
    wire N__12791;
    wire N__12784;
    wire N__12779;
    wire N__12754;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12742;
    wire N__12741;
    wire N__12740;
    wire N__12739;
    wire N__12738;
    wire N__12735;
    wire N__12734;
    wire N__12733;
    wire N__12730;
    wire N__12727;
    wire N__12720;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12700;
    wire N__12697;
    wire N__12696;
    wire N__12689;
    wire N__12686;
    wire N__12677;
    wire N__12670;
    wire N__12661;
    wire N__12660;
    wire N__12659;
    wire N__12654;
    wire N__12653;
    wire N__12650;
    wire N__12649;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12634;
    wire N__12631;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12597;
    wire N__12596;
    wire N__12589;
    wire N__12588;
    wire N__12587;
    wire N__12586;
    wire N__12583;
    wire N__12582;
    wire N__12581;
    wire N__12580;
    wire N__12573;
    wire N__12570;
    wire N__12563;
    wire N__12560;
    wire N__12553;
    wire N__12552;
    wire N__12549;
    wire N__12548;
    wire N__12545;
    wire N__12544;
    wire N__12541;
    wire N__12540;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12510;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12478;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12446;
    wire N__12439;
    wire N__12436;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12412;
    wire N__12411;
    wire N__12410;
    wire N__12409;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12395;
    wire N__12392;
    wire N__12387;
    wire N__12382;
    wire N__12379;
    wire N__12378;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12366;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12349;
    wire N__12348;
    wire N__12345;
    wire N__12344;
    wire N__12343;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12332;
    wire N__12329;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12280;
    wire N__12277;
    wire N__12270;
    wire N__12267;
    wire N__12262;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12246;
    wire N__12243;
    wire N__12240;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12220;
    wire N__12219;
    wire N__12216;
    wire N__12215;
    wire N__12212;
    wire N__12211;
    wire N__12210;
    wire N__12207;
    wire N__12206;
    wire N__12201;
    wire N__12198;
    wire N__12197;
    wire N__12196;
    wire N__12195;
    wire N__12194;
    wire N__12181;
    wire N__12176;
    wire N__12167;
    wire N__12164;
    wire N__12163;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12130;
    wire N__12125;
    wire N__12120;
    wire N__12115;
    wire N__12114;
    wire N__12109;
    wire N__12106;
    wire N__12105;
    wire N__12102;
    wire N__12097;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12085;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12070;
    wire N__12063;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12045;
    wire N__12042;
    wire N__12033;
    wire N__12028;
    wire N__12027;
    wire N__12026;
    wire N__12019;
    wire N__12018;
    wire N__12017;
    wire N__12016;
    wire N__12013;
    wire N__12006;
    wire N__12005;
    wire N__12004;
    wire N__12003;
    wire N__12002;
    wire N__12001;
    wire N__12000;
    wire N__11999;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11991;
    wire N__11976;
    wire N__11971;
    wire N__11968;
    wire N__11959;
    wire N__11958;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11933;
    wire N__11932;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11914;
    wire N__11913;
    wire N__11912;
    wire N__11911;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11884;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11878;
    wire N__11875;
    wire N__11874;
    wire N__11867;
    wire N__11864;
    wire N__11861;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11826;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11809;
    wire N__11806;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11779;
    wire N__11776;
    wire N__11775;
    wire N__11774;
    wire N__11773;
    wire N__11772;
    wire N__11763;
    wire N__11760;
    wire N__11755;
    wire N__11752;
    wire N__11749;
    wire N__11746;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11740;
    wire N__11739;
    wire N__11738;
    wire N__11735;
    wire N__11730;
    wire N__11727;
    wire N__11722;
    wire N__11713;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11705;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11680;
    wire N__11677;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11647;
    wire N__11644;
    wire N__11641;
    wire N__11638;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11614;
    wire N__11611;
    wire N__11608;
    wire N__11605;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11532;
    wire N__11531;
    wire N__11530;
    wire N__11525;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11510;
    wire N__11505;
    wire N__11500;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11474;
    wire N__11467;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11445;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11423;
    wire N__11420;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11408;
    wire N__11401;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11387;
    wire N__11386;
    wire N__11383;
    wire N__11374;
    wire N__11369;
    wire N__11362;
    wire N__11361;
    wire N__11358;
    wire N__11357;
    wire N__11352;
    wire N__11351;
    wire N__11348;
    wire N__11347;
    wire N__11344;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11234;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11205;
    wire N__11202;
    wire N__11201;
    wire N__11200;
    wire N__11199;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11182;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11110;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11095;
    wire N__11090;
    wire N__11087;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11063;
    wire N__11060;
    wire N__11059;
    wire N__11058;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11032;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11007;
    wire N__11006;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10956;
    wire N__10955;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10912;
    wire N__10909;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10885;
    wire N__10884;
    wire N__10881;
    wire N__10880;
    wire N__10877;
    wire N__10872;
    wire N__10869;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10822;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10806;
    wire N__10805;
    wire N__10804;
    wire N__10803;
    wire N__10800;
    wire N__10799;
    wire N__10796;
    wire N__10791;
    wire N__10788;
    wire N__10783;
    wire N__10776;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10760;
    wire N__10759;
    wire N__10758;
    wire N__10753;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10737;
    wire N__10734;
    wire N__10723;
    wire N__10720;
    wire N__10719;
    wire N__10718;
    wire N__10717;
    wire N__10716;
    wire N__10715;
    wire N__10714;
    wire N__10711;
    wire N__10704;
    wire N__10701;
    wire N__10696;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10581;
    wire N__10580;
    wire N__10579;
    wire N__10578;
    wire N__10577;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10561;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10528;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10504;
    wire N__10497;
    wire N__10494;
    wire N__10489;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10483;
    wire N__10482;
    wire N__10481;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10465;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10421;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10383;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10369;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10359;
    wire N__10358;
    wire N__10357;
    wire N__10356;
    wire N__10355;
    wire N__10352;
    wire N__10347;
    wire N__10344;
    wire N__10339;
    wire N__10336;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10226;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10177;
    wire N__10176;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10143;
    wire N__10142;
    wire N__10141;
    wire N__10138;
    wire N__10133;
    wire N__10130;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10078;
    wire N__10077;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10022;
    wire N__10019;
    wire N__10014;
    wire N__10009;
    wire N__10008;
    wire N__10007;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9961;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9879;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9864;
    wire N__9861;
    wire N__9856;
    wire N__9855;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9810;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9798;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9784;
    wire N__9781;
    wire N__9780;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9732;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9711;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9666;
    wire N__9661;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9649;
    wire N__9646;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9598;
    wire N__9595;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9516;
    wire N__9511;
    wire N__9506;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9435;
    wire N__9434;
    wire N__9431;
    wire N__9430;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9405;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9387;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9375;
    wire N__9372;
    wire N__9371;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9347;
    wire N__9340;
    wire N__9339;
    wire N__9336;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9313;
    wire N__9310;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9294;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9268;
    wire N__9267;
    wire N__9264;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9256;
    wire N__9255;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9238;
    wire N__9235;
    wire N__9226;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9216;
    wire N__9211;
    wire N__9206;
    wire N__9199;
    wire N__9196;
    wire N__9195;
    wire N__9194;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9182;
    wire N__9179;
    wire N__9172;
    wire N__9169;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9158;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9146;
    wire N__9143;
    wire N__9136;
    wire N__9133;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9101;
    wire N__9100;
    wire N__9099;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8802;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8790;
    wire N__8789;
    wire N__8788;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8776;
    wire N__8771;
    wire N__8766;
    wire N__8763;
    wire N__8758;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8750;
    wire N__8745;
    wire N__8742;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8647;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8634;
    wire N__8633;
    wire N__8626;
    wire N__8623;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8599;
    wire N__8598;
    wire N__8597;
    wire N__8596;
    wire N__8595;
    wire N__8594;
    wire N__8593;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8589;
    wire N__8588;
    wire N__8585;
    wire N__8578;
    wire N__8569;
    wire N__8566;
    wire N__8559;
    wire N__8556;
    wire N__8551;
    wire N__8542;
    wire N__8541;
    wire N__8540;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8528;
    wire N__8523;
    wire N__8518;
    wire N__8517;
    wire N__8516;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8501;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8487;
    wire N__8486;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8458;
    wire N__8457;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8442;
    wire N__8437;
    wire N__8436;
    wire N__8435;
    wire N__8432;
    wire N__8427;
    wire N__8422;
    wire N__8421;
    wire N__8420;
    wire N__8417;
    wire N__8416;
    wire N__8413;
    wire N__8408;
    wire N__8407;
    wire N__8406;
    wire N__8405;
    wire N__8404;
    wire N__8401;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8383;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8361;
    wire N__8358;
    wire N__8347;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8341;
    wire N__8338;
    wire N__8333;
    wire N__8330;
    wire N__8323;
    wire N__8322;
    wire N__8319;
    wire N__8318;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8302;
    wire N__8301;
    wire N__8300;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8275;
    wire N__8272;
    wire N__8269;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8257;
    wire N__8256;
    wire N__8255;
    wire N__8254;
    wire N__8247;
    wire N__8244;
    wire N__8239;
    wire N__8238;
    wire N__8237;
    wire N__8232;
    wire N__8229;
    wire N__8224;
    wire N__8221;
    wire N__8220;
    wire N__8219;
    wire N__8214;
    wire N__8211;
    wire N__8206;
    wire N__8205;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8176;
    wire N__8173;
    wire N__8172;
    wire N__8171;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8163;
    wire N__8154;
    wire N__8151;
    wire N__8146;
    wire N__8145;
    wire N__8144;
    wire N__8139;
    wire N__8136;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8112;
    wire N__8107;
    wire N__8100;
    wire N__8095;
    wire N__8094;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8074;
    wire N__8073;
    wire N__8072;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7993;
    wire N__7990;
    wire N__7989;
    wire N__7988;
    wire N__7987;
    wire N__7986;
    wire N__7985;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7974;
    wire N__7973;
    wire N__7972;
    wire N__7971;
    wire N__7958;
    wire N__7953;
    wire N__7942;
    wire N__7939;
    wire N__7938;
    wire N__7937;
    wire N__7930;
    wire N__7927;
    wire N__7922;
    wire N__7919;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7888;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7861;
    wire N__7858;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7815;
    wire N__7814;
    wire N__7809;
    wire N__7806;
    wire N__7801;
    wire N__7798;
    wire N__7797;
    wire N__7796;
    wire N__7793;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7777;
    wire N__7776;
    wire N__7775;
    wire N__7772;
    wire N__7767;
    wire N__7762;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7758;
    wire N__7753;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7732;
    wire N__7731;
    wire N__7730;
    wire N__7727;
    wire N__7724;
    wire N__7717;
    wire N__7714;
    wire N__7713;
    wire N__7712;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7700;
    wire N__7695;
    wire N__7690;
    wire N__7689;
    wire N__7688;
    wire N__7687;
    wire N__7680;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7668;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7660;
    wire N__7659;
    wire N__7654;
    wire N__7647;
    wire N__7642;
    wire N__7639;
    wire N__7638;
    wire N__7633;
    wire N__7630;
    wire N__7629;
    wire N__7628;
    wire N__7627;
    wire N__7624;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7572;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7564;
    wire N__7557;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7534;
    wire N__7533;
    wire N__7532;
    wire N__7531;
    wire N__7530;
    wire N__7521;
    wire N__7518;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7506;
    wire N__7503;
    wire N__7502;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7482;
    wire N__7479;
    wire N__7474;
    wire N__7471;
    wire N__7470;
    wire N__7465;
    wire N__7462;
    wire N__7461;
    wire N__7456;
    wire N__7453;
    wire N__7452;
    wire N__7449;
    wire N__7446;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7434;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7415;
    wire N__7412;
    wire N__7407;
    wire N__7402;
    wire N__7401;
    wire N__7400;
    wire N__7399;
    wire N__7394;
    wire N__7389;
    wire N__7384;
    wire N__7381;
    wire N__7380;
    wire N__7379;
    wire N__7378;
    wire N__7371;
    wire N__7368;
    wire N__7363;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7357;
    wire N__7354;
    wire N__7347;
    wire N__7342;
    wire N__7341;
    wire N__7340;
    wire N__7339;
    wire N__7334;
    wire N__7329;
    wire N__7324;
    wire N__7323;
    wire N__7322;
    wire N__7319;
    wire N__7314;
    wire N__7311;
    wire N__7306;
    wire N__7303;
    wire N__7302;
    wire N__7301;
    wire N__7300;
    wire N__7297;
    wire N__7292;
    wire N__7287;
    wire N__7282;
    wire N__7281;
    wire N__7280;
    wire N__7279;
    wire N__7278;
    wire N__7269;
    wire N__7266;
    wire N__7263;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7242;
    wire N__7241;
    wire N__7240;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7221;
    wire N__7220;
    wire N__7219;
    wire N__7218;
    wire N__7217;
    wire N__7204;
    wire N__7201;
    wire N__7198;
    wire N__7195;
    wire N__7192;
    wire N__7189;
    wire N__7188;
    wire N__7185;
    wire N__7182;
    wire N__7177;
    wire N__7176;
    wire N__7175;
    wire N__7168;
    wire N__7165;
    wire N__7164;
    wire N__7163;
    wire N__7160;
    wire N__7155;
    wire N__7150;
    wire N__7147;
    wire N__7146;
    wire N__7145;
    wire N__7144;
    wire N__7143;
    wire N__7140;
    wire N__7139;
    wire N__7126;
    wire N__7123;
    wire N__7122;
    wire N__7121;
    wire N__7120;
    wire N__7119;
    wire N__7110;
    wire N__7107;
    wire N__7102;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7094;
    wire N__7093;
    wire N__7086;
    wire N__7083;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7065;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7048;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7030;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7020;
    wire N__7017;
    wire N__7014;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__7000;
    wire N__6997;
    wire N__6994;
    wire N__6993;
    wire N__6992;
    wire N__6991;
    wire N__6988;
    wire N__6981;
    wire N__6978;
    wire N__6973;
    wire N__6970;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6895;
    wire N__6892;
    wire N__6889;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire \uu2.un284_ci_cascade_ ;
    wire \uu2.un306_ci_cascade_ ;
    wire \uu2.un350_ci_cascade_ ;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.un4_l_count_16_cascade_ ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.un11_l_count_i ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un55_ci_cascade_ ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.un143_ci_0 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.un165_ci_0 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_0_8_cascade_ ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire bfn_2_3_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.un1_bitcount_c3 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \uu2.un350_ci ;
    wire \uu2.un1_l_count_2_2_cascade_ ;
    wire \uu2.un284_ci ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.un1_l_count_1_2_0_cascade_ ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.un306_ci ;
    wire \uu2.r_data_wire_0 ;
    wire vbuf_tx_data_0;
    wire \uu2.r_data_wire_1 ;
    wire vbuf_tx_data_1;
    wire \uu2.r_data_wire_2 ;
    wire vbuf_tx_data_2;
    wire \uu2.r_data_wire_3 ;
    wire vbuf_tx_data_3;
    wire \uu2.r_data_wire_4 ;
    wire vbuf_tx_data_4;
    wire \uu2.r_data_wire_5 ;
    wire vbuf_tx_data_5;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu0.sec_clkDZ0 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu0.un88_ci_3_cascade_ ;
    wire vbuf_tx_data_rdy;
    wire \resetGen.escKeyZ0_cascade_ ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_count_2_0_4 ;
    wire \resetGen.escKeyZ0 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un88_ci_3 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un66_ci ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.un110_ci ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.trig_rd_is_det_cascade_ ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.mem0.N_77_i ;
    wire \uu2.mem0.w_data_i_a3_1_0_cascade_ ;
    wire \uu2.mem0.N_79_i_0 ;
    wire clk;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.N_75_i ;
    wire \uu2.N_361 ;
    wire \uu2.N_361_cascade_ ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.mem0.N_69_i ;
    wire \uu2.mem0.w_data_0_a3_0_4 ;
    wire \uu2.N_61_cascade_ ;
    wire \uu2.mem0.un51_w_data_displaying_cascade_ ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.mem0.N_71_i ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.N_76_i_0 ;
    wire \uu2.mem0.N_2166_0_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_0_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_42 ;
    wire \uu2.mem0.bitmap_pmux_sn_i7_mux_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_43 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_ ;
    wire \uu2.bitmap_RNIMQ601Z0Z_58_cascade_ ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_ ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \INVuu2.bitmap_186C_net ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.bitmap_RNI8LB51Z0Z_186 ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ;
    wire \Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_ ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmapZ0Z_218 ;
    wire o_One_Sec_Pulse;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu0.l_precountZ0Z_0 ;
    wire uart_RXD;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.mem0.N_70_i ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.un404_ci ;
    wire \uu2.bitmap_pmux_20_ns_1_cascade_ ;
    wire \Lab_UT.bcd2segment4.segment_0Z0Z_2 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_ ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \Lab_UT.bcd2segment4.N_217 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \Lab_UT.bcd2segment4.segment_i_1Z0Z_5 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \INVuu2.bitmap_197C_net ;
    wire \uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_ ;
    wire \uu2.mem0.g1_2_0 ;
    wire \uu2.N_40_0 ;
    wire \uu2.N_48_i_0 ;
    wire \uu2.N_404 ;
    wire \uu2.mem0.g1_1_1_0 ;
    wire \uu2.N_404_cascade_ ;
    wire \uu2.mem0.bitmap_pmux_1_0_0 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_42_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_46 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_ ;
    wire \uu2.g2_0_0 ;
    wire \uu2.mem0.g1_6_cascade_ ;
    wire \uu2.mem0.N_1201_0_0_0 ;
    wire \uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0 ;
    wire \uu2.bitmap_pmux_sn_N_20_0 ;
    wire \uu2.bitmap_pmux_19_i_m2_ns_1 ;
    wire \uu2.N_55_0 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_20_1_0_1 ;
    wire \uu2.mem0.N_2166_1_0_1 ;
    wire \uu2.mem0.N_247_0_cascade_ ;
    wire \uu2.mem0.N_2171_1_0_1_cascade_ ;
    wire \uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7 ;
    wire \uu2.mem0.N_397_1_0_1 ;
    wire \uu2.mem0.g1_3_0 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.N_247_cascade_ ;
    wire \uu2.N_2171_0 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_44 ;
    wire \Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_ ;
    wire \Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_ ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.N_383 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ;
    wire \Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_ ;
    wire \INVuu2.bitmap_296C_net ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmap_pmux_15_i_m2_ns_1 ;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.bitmap_pmux_sn_N_54_mux_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_15 ;
    wire \uu2.N_395_cascade_ ;
    wire \uu2.N_56 ;
    wire \uu2.N_401 ;
    wire \buart.Z_rx.idle_1_cascade_ ;
    wire \buart.Z_rx.valid_1_cascade_ ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire bfn_6_3_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \uu2.N_150_cascade_ ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \INVuu2.w_addr_user_nesr_6C_net ;
    wire \uu2.mem0.N_78_i_0 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.N_93 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \Lab_UT.bcd2segment1.segment_0Z0Z_2 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \INVuu2.w_addr_displaying_4C_net ;
    wire \uu2.mem0.g0_7_3_cascade_ ;
    wire \uu2.bitmap_pmux_27_ns_1_0 ;
    wire \uu2.mem0.g0_6_4 ;
    wire \uu2.mem0.g0_6_5_cascade_ ;
    wire \uu2.un426_ci ;
    wire \INVuu2.w_addr_displaying_2_rep1C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \uu2.N_46_cascade_ ;
    wire \INVuu2.w_addr_displaying_fast_nesr_8C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_ ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_ ;
    wire \uu2.N_4_cascade_ ;
    wire \uu2.g0_17_1 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.N_5 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \INVuu2.bitmap_200C_net ;
    wire \Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_ ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.bitmap_RNISSSNZ0Z_162 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_ ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \INVuu2.bitmap_168C_net ;
    wire \Lab_UT.bcd2segment3.segment_i_0Z0Z_1 ;
    wire \Lab_UT.bcd2segment3.segment_i_0Z0Z_2 ;
    wire \resetGen.escKeyZ0Z_3 ;
    wire CONSTANT_ONE_NET;
    wire \buart.Z_rx.N_27_0_i_cascade_ ;
    wire \buart.Z_rx.bitcount_lm_0_cascade_ ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_lm_1_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_lm_2_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \buart.Z_rx.bitcount_lm_4 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \buart.Z_rx.bitcount_lm_3_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \uu2.N_153 ;
    wire \uu2.N_90_cascade_ ;
    wire \uu2.N_105 ;
    wire \uu2.N_90 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.mem0.N_111 ;
    wire \uu2.un28_w_addr_user_i_0_0 ;
    wire \uu2.mem0.N_73_i ;
    wire \uu2.un31_w_data_displaying_0_a2_1_cascade_ ;
    wire \uu2.un31_w_data_displaying ;
    wire \uu2.un15_w_data_displaying_6 ;
    wire \uu2.un15_w_data_displaying_6_cascade_ ;
    wire \uu2.un49_w_data_displaying_1 ;
    wire \uu2.un49_w_data_displaying ;
    wire \uu2.un15_w_data_displaying_i_i_o2_0 ;
    wire \uu2.un15_w_data_displaying_i_i_o2_0_cascade_ ;
    wire \INVuu2.w_addr_displaying_nesr_8C_net ;
    wire \uu2.mem0.un49_w_data_displaying_0 ;
    wire \uu2.mem0.g0_5_5 ;
    wire \uu2.mem0.un31_w_data_displaying_0 ;
    wire \uu2.mem0.g1_1_1 ;
    wire \uu2.w_addr_displaying_7_repZ0Z1 ;
    wire \uu2.w_addr_displaying_8_repZ0Z1 ;
    wire \uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_45 ;
    wire \uu2.w_addr_displaying_2_repZ0Z1 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.bitmap_pmux_sn_N_31_0 ;
    wire \uu2.bitmap_pmux_sn_N_31_0_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_48 ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_ ;
    wire \uu2.mem0.ram512X8_inst_RNOZ0Z_47 ;
    wire \uu2.mem0.bitmap_pmux_u_ns_1 ;
    wire \uu2.mem0.g0_5_3_cascade_ ;
    wire \uu2.mem0.g0_5_6 ;
    wire \Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_ ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.N_7_cascade_ ;
    wire \uu2.N_10 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.N_8 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \INVuu2.bitmap_215C_net ;
    wire \Lab_UT.didp.countrce2.N_178 ;
    wire \Lab_UT.didp.countrce2.N_175 ;
    wire \Lab_UT.didp.countrce2.N_170 ;
    wire \Lab_UT.didp.countrce2.N_183 ;
    wire \Lab_UT.didp.countrce2.N_180 ;
    wire \Lab_UT.didp.countrce4.N_80_i_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_RNO_0Z0Z_3 ;
    wire \Lab_UT.bcd2segment4.segment_i_0Z0Z_6 ;
    wire \Lab_UT.dictrl.next_alarmstate4_1Z0Z_0 ;
    wire \Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_ ;
    wire resetGen_escKey_4_cascade_;
    wire bu_rx_data_5;
    wire bu_rx_data_2;
    wire \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_ ;
    wire bu_rx_data_4;
    wire \Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ;
    wire resetGen_escKey_2_0;
    wire bu_rx_data_6;
    wire bu_rx_data_3;
    wire bu_rx_data_7;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa_2 ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa_1 ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa_cascade_ ;
    wire \Lab_UT.m37_ns_cascade_ ;
    wire \Lab_UT.dictrl.next_state_out_2 ;
    wire \Lab_UT.m45 ;
    wire \Lab_UT.m40_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2 ;
    wire \Lab_UT.dictrl.next_state_out_0 ;
    wire \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.dicRun_2_reti ;
    wire \buart.Z_rx.idle ;
    wire bu_rx_data_rdy;
    wire \buart.Z_rx.bitcountlde_0 ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.ser_clk_2_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.sample ;
    wire bfn_8_3_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.ser_clk_2 ;
    wire \buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ;
    wire \buart.Z_rx.ser_clk_3 ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \Lab_UT.didp.countrce4.q_RNO_0Z0Z_2 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.w_addr_user_3_i_a2_2_6 ;
    wire \uu2.mem0.N_72_i ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.mem0.N_74_i ;
    wire \Lab_UT.dispString.dOutP_0_iv_3_0 ;
    wire \uu2.N_84_cascade_ ;
    wire \uu2.N_97 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.N_97_cascade_ ;
    wire \uu2.N_159 ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire L3_tx_data_0;
    wire \uu2.N_86 ;
    wire L3_tx_data_rdy;
    wire \uu2.N_86_cascade_ ;
    wire \uu2.N_84 ;
    wire \uu2.w_addr_i_0_tzZ0Z_0 ;
    wire \uu2.w_addr_i_0_tzZ0Z_0_cascade_ ;
    wire \uu2.N_61 ;
    wire \uu2.un21_w_addr_displaying_i ;
    wire \uu2.N_49 ;
    wire \uu2.mem0.g0_7_5_0_cascade_ ;
    wire \uu2.mem0.un31_w_data_displaying_1_0_0_cascade_ ;
    wire \uu2.mem0.g1_0_1 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.mem0.g1_0_1_1 ;
    wire \uu2.mem0.g1_5_5 ;
    wire \uu2.w_addr_displaying_3_repZ0Z2 ;
    wire \uu2.mem0.g0_7_4_0 ;
    wire \uu2.N_46 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \INVuu2.w_addr_displaying_nesr_5C_net ;
    wire \uu2.un21_w_addr_displaying_i_0 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.mem0.g0_16_1 ;
    wire \Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_ ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \Lab_UT.nine_cascade_ ;
    wire \Lab_UT.bcd2segment2.segment_i_0Z0Z_1 ;
    wire \Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_ ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \INVuu2.bitmap_93C_net ;
    wire \Lab_UT.three_2_cascade_ ;
    wire \Lab_UT.didp.countrce1.un20_qPone ;
    wire \Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_sqmuxa ;
    wire \Lab_UT.didp.m34_nsZ0Z_1 ;
    wire \Lab_UT.dictrl.next_state16Z0Z_4 ;
    wire \Lab_UT.m34_ns_cascade_ ;
    wire resetGen_escKey_4;
    wire bu_rx_data_1;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \Lab_UT.dictrl.next_state_out_3 ;
    wire \Lab_UT.m34_ns ;
    wire \Lab_UT.didp.N_164_cascade_ ;
    wire \Lab_UT.m42 ;
    wire \Lab_UT.didp.countrce4.N_88_i ;
    wire \Lab_UT.N_68_0 ;
    wire \Lab_UT.didp.un31_reset_i_a4_1 ;
    wire \Lab_UT.dictrl.next_state_set_1 ;
    wire \Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2 ;
    wire \Lab_UT.m37_ns ;
    wire \Lab_UT.Run ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3 ;
    wire \Lab_UT.dictrl.un1_state_12_cascade_ ;
    wire \Lab_UT.didp.m37_nsZ0Z_1 ;
    wire \Lab_UT.state_i_3_1 ;
    wire \Lab_UT.state_2 ;
    wire \Lab_UT.state_3 ;
    wire \Lab_UT.dictrl.un1_state_24_ns_1_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ;
    wire \Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1 ;
    wire \Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ;
    wire \Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_set_0 ;
    wire \Lab_UT.dictrl.next_state_out_1 ;
    wire \Lab_UT.dictrl.un1_state_21_reti_i ;
    wire \Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1 ;
    wire L3_tx_data_5;
    wire \Lab_UT.dispString.dOutP_0_iv_3_2_cascade_ ;
    wire L3_tx_data_2;
    wire L3_tx_data_6;
    wire L3_tx_data_4;
    wire \Lab_UT.dispString.dOutP_0_iv_0_0_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_0 ;
    wire \Lab_UT.un29_dOutP ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_1 ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_1_cascade_ ;
    wire L3_tx_data_1;
    wire \Lab_UT.dispString.dOutP_0_iv_3_1 ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0 ;
    wire \Lab_UT.m24 ;
    wire \Lab_UT.dispString.un22_dOutP ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_3 ;
    wire \Lab_UT.dispString.dOutP_0_iv_3_3_cascade_ ;
    wire L3_tx_data_3;
    wire \Lab_UT.alarmcharZ0Z_0 ;
    wire \Lab_UT.alarmchar9_cascade_ ;
    wire \Lab_UT.alarmcharZ0Z_1 ;
    wire \Lab_UT.zero ;
    wire \Lab_UT.didp.countrce3.qPone_3_cascade_ ;
    wire \Lab_UT.didp.countrce3.N_79_i_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_3 ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.N_207_cascade_ ;
    wire \Lab_UT.didp.q_RNIIKFH3_3 ;
    wire \Lab_UT.m40 ;
    wire \Lab_UT.dictrl.next_state_RNI970UZ0Z_3 ;
    wire \Lab_UT.dictrl.next_state_set_2 ;
    wire \Lab_UT.alarmcharZ0Z_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_2_cascade_ ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_2 ;
    wire \Lab_UT.un3_dOutP ;
    wire \Lab_UT.cnt_3 ;
    wire \Lab_UT.cnt_0 ;
    wire \Lab_UT.cnt_1 ;
    wire \Lab_UT.cnt_2 ;
    wire \Lab_UT.N_204 ;
    wire \Lab_UT.N_204_cascade_ ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.nine ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.di_Stens_0 ;
    wire \Lab_UT.didp.countrce2.three_2 ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.didp.countrce2.three_2_cascade_ ;
    wire \Lab_UT.didp.countrce2.un20_qPone ;
    wire \Lab_UT.di_Mones_3 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.N_207 ;
    wire \Lab_UT.didp.q_RNI84NN1_3 ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.bcd2segment4.G_64_a0Z0Z_1 ;
    wire bu_rx_data_0;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_ ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.dictrl.dicRun_2 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire oneSecStrb_i;
    wire \Lab_UT.state_1 ;
    wire \Lab_UT.dictrl.state_i_3Z0Z_2 ;
    wire \Lab_UT.state_i_3_3 ;
    wire \Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ;
    wire \Lab_UT.dictrl.state_ret_3_RNIDH8UZ0 ;
    wire \Lab_UT.dictrl.state_retZ0Z_4 ;
    wire \Lab_UT.dictrl.next_state_set ;
    wire \Lab_UT.state_0 ;
    wire \Lab_UT.alarmcharZ0Z_4 ;
    wire \Lab_UT.alarmchar_2_1_1_cascade_ ;
    wire \Lab_UT.alarmcharZ0Z_6 ;
    wire \Lab_UT.dictrl.next_alarmstate_1_cascade_ ;
    wire rst;
    wire \Lab_UT.G_3_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ;
    wire \Lab_UT.dictrl.next_alarmstateZ0Z_0 ;
    wire \Lab_UT.alarmMatch ;
    wire \Lab_UT.dictrl.idle ;
    wire \Lab_UT.alarmchar10 ;
    wire \Lab_UT.dictrl.next_alarmstate_1 ;
    wire \Lab_UT.next_alarmstate4 ;
    wire \Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ;
    wire \Lab_UT.alarmstate_1 ;
    wire \Lab_UT.alarmchar10_i_2 ;
    wire \Lab_UT.alarmcharZ0Z_5 ;
    wire \Lab_UT.alarmstate_0 ;
    wire \Lab_UT.bcd2segment4.GZ0Z_1 ;
    wire \Lab_UT.dictrl.next_alarmstate_0_0 ;
    wire \Lab_UT.un1_next_alarmstate21_0 ;
    wire \Lab_UT.dictrl.next_alarmstate_1_0 ;
    wire \Lab_UT.dictrl.alarmstate_i_3_0 ;
    wire _gnd_net_;
    wire clk_g;
    wire rst_g;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__6901),
            .RESETB(N__10413),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__9037,N__9412,N__9442,N__9499,N__9532,N__9301,N__9375,N__9339,N__9267}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__9457,N__8941,N__11848,N__10600,N__12622,N__8890,N__8926,N__8734,N__10060}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__8836,dangling_wire_31,N__8842,dangling_wire_32,N__8869,dangling_wire_33,N__8908,dangling_wire_34,N__8863,dangling_wire_35,N__8932,dangling_wire_36,N__8722}),
            .RCLKE(),
            .RCLK(N__18081),
            .RE(N__10414),
            .WCLKE(N__8679),
            .WCLK(N__18080),
            .WE(N__8689));
    IO_PAD led_obuft_3_iopad (
            .OE(N__18473),
            .DIN(N__18472),
            .DOUT(N__18471),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__18473),
            .PADOUT(N__18472),
            .PADIN(N__18471),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__18464),
            .DIN(N__18463),
            .DOUT(N__18462),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__18464),
            .PADOUT(N__18463),
            .PADIN(N__18462),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__18455),
            .DIN(N__18454),
            .DOUT(N__18453),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__18455),
            .PADOUT(N__18454),
            .PADIN(N__18453),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__18446),
            .DIN(N__18445),
            .DOUT(N__18444),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__18446),
            .PADOUT(N__18445),
            .PADIN(N__18444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__18437),
            .DIN(N__18436),
            .DOUT(N__18435),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__18437),
            .PADOUT(N__18436),
            .PADIN(N__18435),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__18076),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__18428),
            .DIN(N__18427),
            .DOUT(N__18426),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__18428),
            .PADOUT(N__18427),
            .PADIN(N__18426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__18419),
            .DIN(N__18418),
            .DOUT(N__18417),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__18419),
            .PADOUT(N__18418),
            .PADIN(N__18417),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__18410),
            .DIN(N__18409),
            .DOUT(N__18408),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__18410),
            .PADOUT(N__18409),
            .PADIN(N__18408),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__18401),
            .DIN(N__18400),
            .DOUT(N__18399),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__18401),
            .PADOUT(N__18400),
            .PADIN(N__18399),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__18392),
            .DIN(N__18391),
            .DOUT(N__18390),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__18392),
            .PADOUT(N__18391),
            .PADIN(N__18390),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6913),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__4412 (
            .O(N__18373),
            .I(N__18370));
    LocalMux I__4411 (
            .O(N__18370),
            .I(N__18367));
    Odrv4 I__4410 (
            .O(N__18367),
            .I(\Lab_UT.alarmchar10 ));
    InMux I__4409 (
            .O(N__18364),
            .I(N__18358));
    InMux I__4408 (
            .O(N__18363),
            .I(N__18358));
    LocalMux I__4407 (
            .O(N__18358),
            .I(\Lab_UT.dictrl.next_alarmstate_1 ));
    InMux I__4406 (
            .O(N__18355),
            .I(N__18349));
    InMux I__4405 (
            .O(N__18354),
            .I(N__18342));
    InMux I__4404 (
            .O(N__18353),
            .I(N__18342));
    InMux I__4403 (
            .O(N__18352),
            .I(N__18342));
    LocalMux I__4402 (
            .O(N__18349),
            .I(N__18337));
    LocalMux I__4401 (
            .O(N__18342),
            .I(N__18337));
    Span12Mux_s10_v I__4400 (
            .O(N__18337),
            .I(N__18334));
    Odrv12 I__4399 (
            .O(N__18334),
            .I(\Lab_UT.next_alarmstate4 ));
    InMux I__4398 (
            .O(N__18331),
            .I(N__18327));
    InMux I__4397 (
            .O(N__18330),
            .I(N__18324));
    LocalMux I__4396 (
            .O(N__18327),
            .I(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ));
    LocalMux I__4395 (
            .O(N__18324),
            .I(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ));
    InMux I__4394 (
            .O(N__18319),
            .I(N__18309));
    InMux I__4393 (
            .O(N__18318),
            .I(N__18309));
    InMux I__4392 (
            .O(N__18317),
            .I(N__18309));
    InMux I__4391 (
            .O(N__18316),
            .I(N__18306));
    LocalMux I__4390 (
            .O(N__18309),
            .I(N__18300));
    LocalMux I__4389 (
            .O(N__18306),
            .I(N__18297));
    InMux I__4388 (
            .O(N__18305),
            .I(N__18290));
    InMux I__4387 (
            .O(N__18304),
            .I(N__18290));
    InMux I__4386 (
            .O(N__18303),
            .I(N__18290));
    Odrv4 I__4385 (
            .O(N__18300),
            .I(\Lab_UT.alarmstate_1 ));
    Odrv4 I__4384 (
            .O(N__18297),
            .I(\Lab_UT.alarmstate_1 ));
    LocalMux I__4383 (
            .O(N__18290),
            .I(\Lab_UT.alarmstate_1 ));
    InMux I__4382 (
            .O(N__18283),
            .I(N__18280));
    LocalMux I__4381 (
            .O(N__18280),
            .I(\Lab_UT.alarmchar10_i_2 ));
    CascadeMux I__4380 (
            .O(N__18277),
            .I(N__18274));
    InMux I__4379 (
            .O(N__18274),
            .I(N__18271));
    LocalMux I__4378 (
            .O(N__18271),
            .I(N__18268));
    Span4Mux_v I__4377 (
            .O(N__18268),
            .I(N__18265));
    Odrv4 I__4376 (
            .O(N__18265),
            .I(\Lab_UT.alarmcharZ0Z_5 ));
    InMux I__4375 (
            .O(N__18262),
            .I(N__18257));
    InMux I__4374 (
            .O(N__18261),
            .I(N__18254));
    CascadeMux I__4373 (
            .O(N__18260),
            .I(N__18250));
    LocalMux I__4372 (
            .O(N__18257),
            .I(N__18245));
    LocalMux I__4371 (
            .O(N__18254),
            .I(N__18245));
    InMux I__4370 (
            .O(N__18253),
            .I(N__18242));
    InMux I__4369 (
            .O(N__18250),
            .I(N__18239));
    Odrv4 I__4368 (
            .O(N__18245),
            .I(\Lab_UT.alarmstate_0 ));
    LocalMux I__4367 (
            .O(N__18242),
            .I(\Lab_UT.alarmstate_0 ));
    LocalMux I__4366 (
            .O(N__18239),
            .I(\Lab_UT.alarmstate_0 ));
    CascadeMux I__4365 (
            .O(N__18232),
            .I(N__18229));
    InMux I__4364 (
            .O(N__18229),
            .I(N__18226));
    LocalMux I__4363 (
            .O(N__18226),
            .I(\Lab_UT.bcd2segment4.GZ0Z_1 ));
    CascadeMux I__4362 (
            .O(N__18223),
            .I(N__18219));
    InMux I__4361 (
            .O(N__18222),
            .I(N__18212));
    InMux I__4360 (
            .O(N__18219),
            .I(N__18207));
    InMux I__4359 (
            .O(N__18218),
            .I(N__18207));
    InMux I__4358 (
            .O(N__18217),
            .I(N__18204));
    InMux I__4357 (
            .O(N__18216),
            .I(N__18199));
    InMux I__4356 (
            .O(N__18215),
            .I(N__18199));
    LocalMux I__4355 (
            .O(N__18212),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    LocalMux I__4354 (
            .O(N__18207),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    LocalMux I__4353 (
            .O(N__18204),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    LocalMux I__4352 (
            .O(N__18199),
            .I(\Lab_UT.dictrl.next_alarmstate_0_0 ));
    CascadeMux I__4351 (
            .O(N__18190),
            .I(N__18182));
    InMux I__4350 (
            .O(N__18189),
            .I(N__18173));
    InMux I__4349 (
            .O(N__18188),
            .I(N__18173));
    InMux I__4348 (
            .O(N__18187),
            .I(N__18173));
    InMux I__4347 (
            .O(N__18186),
            .I(N__18170));
    InMux I__4346 (
            .O(N__18185),
            .I(N__18167));
    InMux I__4345 (
            .O(N__18182),
            .I(N__18162));
    InMux I__4344 (
            .O(N__18181),
            .I(N__18162));
    InMux I__4343 (
            .O(N__18180),
            .I(N__18159));
    LocalMux I__4342 (
            .O(N__18173),
            .I(\Lab_UT.un1_next_alarmstate21_0 ));
    LocalMux I__4341 (
            .O(N__18170),
            .I(\Lab_UT.un1_next_alarmstate21_0 ));
    LocalMux I__4340 (
            .O(N__18167),
            .I(\Lab_UT.un1_next_alarmstate21_0 ));
    LocalMux I__4339 (
            .O(N__18162),
            .I(\Lab_UT.un1_next_alarmstate21_0 ));
    LocalMux I__4338 (
            .O(N__18159),
            .I(\Lab_UT.un1_next_alarmstate21_0 ));
    InMux I__4337 (
            .O(N__18148),
            .I(N__18142));
    InMux I__4336 (
            .O(N__18147),
            .I(N__18139));
    InMux I__4335 (
            .O(N__18146),
            .I(N__18134));
    InMux I__4334 (
            .O(N__18145),
            .I(N__18134));
    LocalMux I__4333 (
            .O(N__18142),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    LocalMux I__4332 (
            .O(N__18139),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    LocalMux I__4331 (
            .O(N__18134),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0 ));
    InMux I__4330 (
            .O(N__18127),
            .I(N__18123));
    InMux I__4329 (
            .O(N__18126),
            .I(N__18120));
    LocalMux I__4328 (
            .O(N__18123),
            .I(N__18115));
    LocalMux I__4327 (
            .O(N__18120),
            .I(N__18112));
    InMux I__4326 (
            .O(N__18119),
            .I(N__18109));
    InMux I__4325 (
            .O(N__18118),
            .I(N__18106));
    Odrv4 I__4324 (
            .O(N__18115),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    Odrv4 I__4323 (
            .O(N__18112),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__4322 (
            .O(N__18109),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    LocalMux I__4321 (
            .O(N__18106),
            .I(\Lab_UT.dictrl.alarmstate_i_3_0 ));
    ClkMux I__4320 (
            .O(N__18097),
            .I(N__17863));
    ClkMux I__4319 (
            .O(N__18096),
            .I(N__17863));
    ClkMux I__4318 (
            .O(N__18095),
            .I(N__17863));
    ClkMux I__4317 (
            .O(N__18094),
            .I(N__17863));
    ClkMux I__4316 (
            .O(N__18093),
            .I(N__17863));
    ClkMux I__4315 (
            .O(N__18092),
            .I(N__17863));
    ClkMux I__4314 (
            .O(N__18091),
            .I(N__17863));
    ClkMux I__4313 (
            .O(N__18090),
            .I(N__17863));
    ClkMux I__4312 (
            .O(N__18089),
            .I(N__17863));
    ClkMux I__4311 (
            .O(N__18088),
            .I(N__17863));
    ClkMux I__4310 (
            .O(N__18087),
            .I(N__17863));
    ClkMux I__4309 (
            .O(N__18086),
            .I(N__17863));
    ClkMux I__4308 (
            .O(N__18085),
            .I(N__17863));
    ClkMux I__4307 (
            .O(N__18084),
            .I(N__17863));
    ClkMux I__4306 (
            .O(N__18083),
            .I(N__17863));
    ClkMux I__4305 (
            .O(N__18082),
            .I(N__17863));
    ClkMux I__4304 (
            .O(N__18081),
            .I(N__17863));
    ClkMux I__4303 (
            .O(N__18080),
            .I(N__17863));
    ClkMux I__4302 (
            .O(N__18079),
            .I(N__17863));
    ClkMux I__4301 (
            .O(N__18078),
            .I(N__17863));
    ClkMux I__4300 (
            .O(N__18077),
            .I(N__17863));
    ClkMux I__4299 (
            .O(N__18076),
            .I(N__17863));
    ClkMux I__4298 (
            .O(N__18075),
            .I(N__17863));
    ClkMux I__4297 (
            .O(N__18074),
            .I(N__17863));
    ClkMux I__4296 (
            .O(N__18073),
            .I(N__17863));
    ClkMux I__4295 (
            .O(N__18072),
            .I(N__17863));
    ClkMux I__4294 (
            .O(N__18071),
            .I(N__17863));
    ClkMux I__4293 (
            .O(N__18070),
            .I(N__17863));
    ClkMux I__4292 (
            .O(N__18069),
            .I(N__17863));
    ClkMux I__4291 (
            .O(N__18068),
            .I(N__17863));
    ClkMux I__4290 (
            .O(N__18067),
            .I(N__17863));
    ClkMux I__4289 (
            .O(N__18066),
            .I(N__17863));
    ClkMux I__4288 (
            .O(N__18065),
            .I(N__17863));
    ClkMux I__4287 (
            .O(N__18064),
            .I(N__17863));
    ClkMux I__4286 (
            .O(N__18063),
            .I(N__17863));
    ClkMux I__4285 (
            .O(N__18062),
            .I(N__17863));
    ClkMux I__4284 (
            .O(N__18061),
            .I(N__17863));
    ClkMux I__4283 (
            .O(N__18060),
            .I(N__17863));
    ClkMux I__4282 (
            .O(N__18059),
            .I(N__17863));
    ClkMux I__4281 (
            .O(N__18058),
            .I(N__17863));
    ClkMux I__4280 (
            .O(N__18057),
            .I(N__17863));
    ClkMux I__4279 (
            .O(N__18056),
            .I(N__17863));
    ClkMux I__4278 (
            .O(N__18055),
            .I(N__17863));
    ClkMux I__4277 (
            .O(N__18054),
            .I(N__17863));
    ClkMux I__4276 (
            .O(N__18053),
            .I(N__17863));
    ClkMux I__4275 (
            .O(N__18052),
            .I(N__17863));
    ClkMux I__4274 (
            .O(N__18051),
            .I(N__17863));
    ClkMux I__4273 (
            .O(N__18050),
            .I(N__17863));
    ClkMux I__4272 (
            .O(N__18049),
            .I(N__17863));
    ClkMux I__4271 (
            .O(N__18048),
            .I(N__17863));
    ClkMux I__4270 (
            .O(N__18047),
            .I(N__17863));
    ClkMux I__4269 (
            .O(N__18046),
            .I(N__17863));
    ClkMux I__4268 (
            .O(N__18045),
            .I(N__17863));
    ClkMux I__4267 (
            .O(N__18044),
            .I(N__17863));
    ClkMux I__4266 (
            .O(N__18043),
            .I(N__17863));
    ClkMux I__4265 (
            .O(N__18042),
            .I(N__17863));
    ClkMux I__4264 (
            .O(N__18041),
            .I(N__17863));
    ClkMux I__4263 (
            .O(N__18040),
            .I(N__17863));
    ClkMux I__4262 (
            .O(N__18039),
            .I(N__17863));
    ClkMux I__4261 (
            .O(N__18038),
            .I(N__17863));
    ClkMux I__4260 (
            .O(N__18037),
            .I(N__17863));
    ClkMux I__4259 (
            .O(N__18036),
            .I(N__17863));
    ClkMux I__4258 (
            .O(N__18035),
            .I(N__17863));
    ClkMux I__4257 (
            .O(N__18034),
            .I(N__17863));
    ClkMux I__4256 (
            .O(N__18033),
            .I(N__17863));
    ClkMux I__4255 (
            .O(N__18032),
            .I(N__17863));
    ClkMux I__4254 (
            .O(N__18031),
            .I(N__17863));
    ClkMux I__4253 (
            .O(N__18030),
            .I(N__17863));
    ClkMux I__4252 (
            .O(N__18029),
            .I(N__17863));
    ClkMux I__4251 (
            .O(N__18028),
            .I(N__17863));
    ClkMux I__4250 (
            .O(N__18027),
            .I(N__17863));
    ClkMux I__4249 (
            .O(N__18026),
            .I(N__17863));
    ClkMux I__4248 (
            .O(N__18025),
            .I(N__17863));
    ClkMux I__4247 (
            .O(N__18024),
            .I(N__17863));
    ClkMux I__4246 (
            .O(N__18023),
            .I(N__17863));
    ClkMux I__4245 (
            .O(N__18022),
            .I(N__17863));
    ClkMux I__4244 (
            .O(N__18021),
            .I(N__17863));
    ClkMux I__4243 (
            .O(N__18020),
            .I(N__17863));
    GlobalMux I__4242 (
            .O(N__17863),
            .I(N__17860));
    gio2CtrlBuf I__4241 (
            .O(N__17860),
            .I(clk_g));
    InMux I__4240 (
            .O(N__17857),
            .I(N__17847));
    InMux I__4239 (
            .O(N__17856),
            .I(N__17847));
    InMux I__4238 (
            .O(N__17855),
            .I(N__17844));
    InMux I__4237 (
            .O(N__17854),
            .I(N__17841));
    InMux I__4236 (
            .O(N__17853),
            .I(N__17838));
    InMux I__4235 (
            .O(N__17852),
            .I(N__17835));
    LocalMux I__4234 (
            .O(N__17847),
            .I(N__17802));
    LocalMux I__4233 (
            .O(N__17844),
            .I(N__17799));
    LocalMux I__4232 (
            .O(N__17841),
            .I(N__17796));
    LocalMux I__4231 (
            .O(N__17838),
            .I(N__17793));
    LocalMux I__4230 (
            .O(N__17835),
            .I(N__17773));
    SRMux I__4229 (
            .O(N__17834),
            .I(N__17668));
    SRMux I__4228 (
            .O(N__17833),
            .I(N__17668));
    SRMux I__4227 (
            .O(N__17832),
            .I(N__17668));
    SRMux I__4226 (
            .O(N__17831),
            .I(N__17668));
    SRMux I__4225 (
            .O(N__17830),
            .I(N__17668));
    SRMux I__4224 (
            .O(N__17829),
            .I(N__17668));
    SRMux I__4223 (
            .O(N__17828),
            .I(N__17668));
    SRMux I__4222 (
            .O(N__17827),
            .I(N__17668));
    SRMux I__4221 (
            .O(N__17826),
            .I(N__17668));
    SRMux I__4220 (
            .O(N__17825),
            .I(N__17668));
    SRMux I__4219 (
            .O(N__17824),
            .I(N__17668));
    SRMux I__4218 (
            .O(N__17823),
            .I(N__17668));
    SRMux I__4217 (
            .O(N__17822),
            .I(N__17668));
    SRMux I__4216 (
            .O(N__17821),
            .I(N__17668));
    SRMux I__4215 (
            .O(N__17820),
            .I(N__17668));
    SRMux I__4214 (
            .O(N__17819),
            .I(N__17668));
    SRMux I__4213 (
            .O(N__17818),
            .I(N__17668));
    SRMux I__4212 (
            .O(N__17817),
            .I(N__17668));
    SRMux I__4211 (
            .O(N__17816),
            .I(N__17668));
    SRMux I__4210 (
            .O(N__17815),
            .I(N__17668));
    SRMux I__4209 (
            .O(N__17814),
            .I(N__17668));
    SRMux I__4208 (
            .O(N__17813),
            .I(N__17668));
    SRMux I__4207 (
            .O(N__17812),
            .I(N__17668));
    SRMux I__4206 (
            .O(N__17811),
            .I(N__17668));
    SRMux I__4205 (
            .O(N__17810),
            .I(N__17668));
    SRMux I__4204 (
            .O(N__17809),
            .I(N__17668));
    SRMux I__4203 (
            .O(N__17808),
            .I(N__17668));
    SRMux I__4202 (
            .O(N__17807),
            .I(N__17668));
    SRMux I__4201 (
            .O(N__17806),
            .I(N__17668));
    SRMux I__4200 (
            .O(N__17805),
            .I(N__17668));
    Glb2LocalMux I__4199 (
            .O(N__17802),
            .I(N__17668));
    Glb2LocalMux I__4198 (
            .O(N__17799),
            .I(N__17668));
    Glb2LocalMux I__4197 (
            .O(N__17796),
            .I(N__17668));
    Glb2LocalMux I__4196 (
            .O(N__17793),
            .I(N__17668));
    SRMux I__4195 (
            .O(N__17792),
            .I(N__17668));
    SRMux I__4194 (
            .O(N__17791),
            .I(N__17668));
    SRMux I__4193 (
            .O(N__17790),
            .I(N__17668));
    SRMux I__4192 (
            .O(N__17789),
            .I(N__17668));
    SRMux I__4191 (
            .O(N__17788),
            .I(N__17668));
    SRMux I__4190 (
            .O(N__17787),
            .I(N__17668));
    SRMux I__4189 (
            .O(N__17786),
            .I(N__17668));
    SRMux I__4188 (
            .O(N__17785),
            .I(N__17668));
    SRMux I__4187 (
            .O(N__17784),
            .I(N__17668));
    SRMux I__4186 (
            .O(N__17783),
            .I(N__17668));
    SRMux I__4185 (
            .O(N__17782),
            .I(N__17668));
    SRMux I__4184 (
            .O(N__17781),
            .I(N__17668));
    SRMux I__4183 (
            .O(N__17780),
            .I(N__17668));
    SRMux I__4182 (
            .O(N__17779),
            .I(N__17668));
    SRMux I__4181 (
            .O(N__17778),
            .I(N__17668));
    SRMux I__4180 (
            .O(N__17777),
            .I(N__17668));
    SRMux I__4179 (
            .O(N__17776),
            .I(N__17668));
    Glb2LocalMux I__4178 (
            .O(N__17773),
            .I(N__17668));
    GlobalMux I__4177 (
            .O(N__17668),
            .I(N__17665));
    gio2CtrlBuf I__4176 (
            .O(N__17665),
            .I(rst_g));
    CascadeMux I__4175 (
            .O(N__17662),
            .I(\Lab_UT.alarmchar_2_1_1_cascade_ ));
    InMux I__4174 (
            .O(N__17659),
            .I(N__17656));
    LocalMux I__4173 (
            .O(N__17656),
            .I(N__17653));
    Odrv4 I__4172 (
            .O(N__17653),
            .I(\Lab_UT.alarmcharZ0Z_6 ));
    CascadeMux I__4171 (
            .O(N__17650),
            .I(\Lab_UT.dictrl.next_alarmstate_1_cascade_ ));
    IoInMux I__4170 (
            .O(N__17647),
            .I(N__17639));
    InMux I__4169 (
            .O(N__17646),
            .I(N__17632));
    InMux I__4168 (
            .O(N__17645),
            .I(N__17632));
    InMux I__4167 (
            .O(N__17644),
            .I(N__17625));
    InMux I__4166 (
            .O(N__17643),
            .I(N__17625));
    InMux I__4165 (
            .O(N__17642),
            .I(N__17625));
    LocalMux I__4164 (
            .O(N__17639),
            .I(N__17622));
    InMux I__4163 (
            .O(N__17638),
            .I(N__17617));
    InMux I__4162 (
            .O(N__17637),
            .I(N__17617));
    LocalMux I__4161 (
            .O(N__17632),
            .I(N__17614));
    LocalMux I__4160 (
            .O(N__17625),
            .I(N__17611));
    Span4Mux_s3_h I__4159 (
            .O(N__17622),
            .I(N__17608));
    LocalMux I__4158 (
            .O(N__17617),
            .I(N__17603));
    Span12Mux_s4_h I__4157 (
            .O(N__17614),
            .I(N__17603));
    Span4Mux_v I__4156 (
            .O(N__17611),
            .I(N__17598));
    Span4Mux_h I__4155 (
            .O(N__17608),
            .I(N__17598));
    Odrv12 I__4154 (
            .O(N__17603),
            .I(rst));
    Odrv4 I__4153 (
            .O(N__17598),
            .I(rst));
    CascadeMux I__4152 (
            .O(N__17593),
            .I(\Lab_UT.G_3_cascade_ ));
    CascadeMux I__4151 (
            .O(N__17590),
            .I(\Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ));
    InMux I__4150 (
            .O(N__17587),
            .I(N__17584));
    LocalMux I__4149 (
            .O(N__17584),
            .I(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ));
    InMux I__4148 (
            .O(N__17581),
            .I(N__17572));
    InMux I__4147 (
            .O(N__17580),
            .I(N__17572));
    InMux I__4146 (
            .O(N__17579),
            .I(N__17572));
    LocalMux I__4145 (
            .O(N__17572),
            .I(N__17569));
    Odrv4 I__4144 (
            .O(N__17569),
            .I(\Lab_UT.alarmMatch ));
    InMux I__4143 (
            .O(N__17566),
            .I(N__17563));
    LocalMux I__4142 (
            .O(N__17563),
            .I(\Lab_UT.dictrl.idle ));
    CascadeMux I__4141 (
            .O(N__17560),
            .I(N__17555));
    InMux I__4140 (
            .O(N__17559),
            .I(N__17552));
    InMux I__4139 (
            .O(N__17558),
            .I(N__17539));
    InMux I__4138 (
            .O(N__17555),
            .I(N__17536));
    LocalMux I__4137 (
            .O(N__17552),
            .I(N__17533));
    InMux I__4136 (
            .O(N__17551),
            .I(N__17528));
    InMux I__4135 (
            .O(N__17550),
            .I(N__17528));
    InMux I__4134 (
            .O(N__17549),
            .I(N__17523));
    InMux I__4133 (
            .O(N__17548),
            .I(N__17523));
    InMux I__4132 (
            .O(N__17547),
            .I(N__17520));
    InMux I__4131 (
            .O(N__17546),
            .I(N__17509));
    InMux I__4130 (
            .O(N__17545),
            .I(N__17509));
    InMux I__4129 (
            .O(N__17544),
            .I(N__17509));
    InMux I__4128 (
            .O(N__17543),
            .I(N__17509));
    InMux I__4127 (
            .O(N__17542),
            .I(N__17509));
    LocalMux I__4126 (
            .O(N__17539),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4125 (
            .O(N__17536),
            .I(\Lab_UT.di_Stens_3 ));
    Odrv4 I__4124 (
            .O(N__17533),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4123 (
            .O(N__17528),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4122 (
            .O(N__17523),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4121 (
            .O(N__17520),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__4120 (
            .O(N__17509),
            .I(\Lab_UT.di_Stens_3 ));
    CascadeMux I__4119 (
            .O(N__17494),
            .I(N__17489));
    InMux I__4118 (
            .O(N__17493),
            .I(N__17483));
    InMux I__4117 (
            .O(N__17492),
            .I(N__17480));
    InMux I__4116 (
            .O(N__17489),
            .I(N__17475));
    InMux I__4115 (
            .O(N__17488),
            .I(N__17475));
    InMux I__4114 (
            .O(N__17487),
            .I(N__17466));
    InMux I__4113 (
            .O(N__17486),
            .I(N__17466));
    LocalMux I__4112 (
            .O(N__17483),
            .I(N__17463));
    LocalMux I__4111 (
            .O(N__17480),
            .I(N__17460));
    LocalMux I__4110 (
            .O(N__17475),
            .I(N__17457));
    InMux I__4109 (
            .O(N__17474),
            .I(N__17454));
    InMux I__4108 (
            .O(N__17473),
            .I(N__17447));
    InMux I__4107 (
            .O(N__17472),
            .I(N__17447));
    InMux I__4106 (
            .O(N__17471),
            .I(N__17444));
    LocalMux I__4105 (
            .O(N__17466),
            .I(N__17441));
    Span4Mux_h I__4104 (
            .O(N__17463),
            .I(N__17434));
    Span4Mux_v I__4103 (
            .O(N__17460),
            .I(N__17434));
    Span4Mux_h I__4102 (
            .O(N__17457),
            .I(N__17434));
    LocalMux I__4101 (
            .O(N__17454),
            .I(N__17431));
    InMux I__4100 (
            .O(N__17453),
            .I(N__17426));
    InMux I__4099 (
            .O(N__17452),
            .I(N__17426));
    LocalMux I__4098 (
            .O(N__17447),
            .I(N__17421));
    LocalMux I__4097 (
            .O(N__17444),
            .I(N__17421));
    Span4Mux_h I__4096 (
            .O(N__17441),
            .I(N__17416));
    Span4Mux_v I__4095 (
            .O(N__17434),
            .I(N__17416));
    Span4Mux_h I__4094 (
            .O(N__17431),
            .I(N__17409));
    LocalMux I__4093 (
            .O(N__17426),
            .I(N__17409));
    Span4Mux_h I__4092 (
            .O(N__17421),
            .I(N__17409));
    Odrv4 I__4091 (
            .O(N__17416),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__4090 (
            .O(N__17409),
            .I(\Lab_UT.di_Mtens_3 ));
    InMux I__4089 (
            .O(N__17404),
            .I(N__17401));
    LocalMux I__4088 (
            .O(N__17401),
            .I(N__17398));
    Odrv12 I__4087 (
            .O(N__17398),
            .I(\Lab_UT.bcd2segment4.G_64_a0Z0Z_1 ));
    InMux I__4086 (
            .O(N__17395),
            .I(N__17392));
    LocalMux I__4085 (
            .O(N__17392),
            .I(N__17389));
    Span4Mux_h I__4084 (
            .O(N__17389),
            .I(N__17382));
    InMux I__4083 (
            .O(N__17388),
            .I(N__17377));
    InMux I__4082 (
            .O(N__17387),
            .I(N__17377));
    InMux I__4081 (
            .O(N__17386),
            .I(N__17372));
    InMux I__4080 (
            .O(N__17385),
            .I(N__17372));
    Odrv4 I__4079 (
            .O(N__17382),
            .I(bu_rx_data_0));
    LocalMux I__4078 (
            .O(N__17377),
            .I(bu_rx_data_0));
    LocalMux I__4077 (
            .O(N__17372),
            .I(bu_rx_data_0));
    CascadeMux I__4076 (
            .O(N__17365),
            .I(N__17359));
    InMux I__4075 (
            .O(N__17364),
            .I(N__17356));
    InMux I__4074 (
            .O(N__17363),
            .I(N__17351));
    InMux I__4073 (
            .O(N__17362),
            .I(N__17351));
    InMux I__4072 (
            .O(N__17359),
            .I(N__17348));
    LocalMux I__4071 (
            .O(N__17356),
            .I(\Lab_UT.LdMtens ));
    LocalMux I__4070 (
            .O(N__17351),
            .I(\Lab_UT.LdMtens ));
    LocalMux I__4069 (
            .O(N__17348),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__4068 (
            .O(N__17341),
            .I(N__17337));
    InMux I__4067 (
            .O(N__17340),
            .I(N__17332));
    InMux I__4066 (
            .O(N__17337),
            .I(N__17329));
    CascadeMux I__4065 (
            .O(N__17336),
            .I(N__17326));
    InMux I__4064 (
            .O(N__17335),
            .I(N__17323));
    LocalMux I__4063 (
            .O(N__17332),
            .I(N__17320));
    LocalMux I__4062 (
            .O(N__17329),
            .I(N__17317));
    InMux I__4061 (
            .O(N__17326),
            .I(N__17314));
    LocalMux I__4060 (
            .O(N__17323),
            .I(N__17311));
    Span4Mux_v I__4059 (
            .O(N__17320),
            .I(N__17308));
    Span4Mux_v I__4058 (
            .O(N__17317),
            .I(N__17303));
    LocalMux I__4057 (
            .O(N__17314),
            .I(N__17303));
    Odrv12 I__4056 (
            .O(N__17311),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    Odrv4 I__4055 (
            .O(N__17308),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    Odrv4 I__4054 (
            .O(N__17303),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    CascadeMux I__4053 (
            .O(N__17296),
            .I(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_ ));
    InMux I__4052 (
            .O(N__17293),
            .I(N__17289));
    InMux I__4051 (
            .O(N__17292),
            .I(N__17286));
    LocalMux I__4050 (
            .O(N__17289),
            .I(N__17282));
    LocalMux I__4049 (
            .O(N__17286),
            .I(N__17279));
    InMux I__4048 (
            .O(N__17285),
            .I(N__17276));
    Span4Mux_v I__4047 (
            .O(N__17282),
            .I(N__17272));
    Span4Mux_v I__4046 (
            .O(N__17279),
            .I(N__17269));
    LocalMux I__4045 (
            .O(N__17276),
            .I(N__17266));
    InMux I__4044 (
            .O(N__17275),
            .I(N__17263));
    Odrv4 I__4043 (
            .O(N__17272),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv4 I__4042 (
            .O(N__17269),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv4 I__4041 (
            .O(N__17266),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    LocalMux I__4040 (
            .O(N__17263),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    InMux I__4039 (
            .O(N__17254),
            .I(N__17243));
    InMux I__4038 (
            .O(N__17253),
            .I(N__17243));
    InMux I__4037 (
            .O(N__17252),
            .I(N__17240));
    InMux I__4036 (
            .O(N__17251),
            .I(N__17231));
    InMux I__4035 (
            .O(N__17250),
            .I(N__17231));
    InMux I__4034 (
            .O(N__17249),
            .I(N__17231));
    InMux I__4033 (
            .O(N__17248),
            .I(N__17231));
    LocalMux I__4032 (
            .O(N__17243),
            .I(N__17227));
    LocalMux I__4031 (
            .O(N__17240),
            .I(N__17222));
    LocalMux I__4030 (
            .O(N__17231),
            .I(N__17222));
    InMux I__4029 (
            .O(N__17230),
            .I(N__17216));
    Span4Mux_v I__4028 (
            .O(N__17227),
            .I(N__17209));
    Span4Mux_v I__4027 (
            .O(N__17222),
            .I(N__17209));
    InMux I__4026 (
            .O(N__17221),
            .I(N__17204));
    InMux I__4025 (
            .O(N__17220),
            .I(N__17204));
    InMux I__4024 (
            .O(N__17219),
            .I(N__17198));
    LocalMux I__4023 (
            .O(N__17216),
            .I(N__17195));
    InMux I__4022 (
            .O(N__17215),
            .I(N__17190));
    InMux I__4021 (
            .O(N__17214),
            .I(N__17190));
    Span4Mux_h I__4020 (
            .O(N__17209),
            .I(N__17187));
    LocalMux I__4019 (
            .O(N__17204),
            .I(N__17184));
    InMux I__4018 (
            .O(N__17203),
            .I(N__17177));
    InMux I__4017 (
            .O(N__17202),
            .I(N__17177));
    InMux I__4016 (
            .O(N__17201),
            .I(N__17177));
    LocalMux I__4015 (
            .O(N__17198),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv12 I__4014 (
            .O(N__17195),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4013 (
            .O(N__17190),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__4012 (
            .O(N__17187),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv12 I__4011 (
            .O(N__17184),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__4010 (
            .O(N__17177),
            .I(\Lab_UT.di_Mtens_0 ));
    InMux I__4009 (
            .O(N__17164),
            .I(N__17159));
    InMux I__4008 (
            .O(N__17163),
            .I(N__17156));
    InMux I__4007 (
            .O(N__17162),
            .I(N__17153));
    LocalMux I__4006 (
            .O(N__17159),
            .I(\Lab_UT.dictrl.dicRun_2 ));
    LocalMux I__4005 (
            .O(N__17156),
            .I(\Lab_UT.dictrl.dicRun_2 ));
    LocalMux I__4004 (
            .O(N__17153),
            .I(\Lab_UT.dictrl.dicRun_2 ));
    InMux I__4003 (
            .O(N__17146),
            .I(N__17134));
    InMux I__4002 (
            .O(N__17145),
            .I(N__17134));
    InMux I__4001 (
            .O(N__17144),
            .I(N__17134));
    InMux I__4000 (
            .O(N__17143),
            .I(N__17134));
    LocalMux I__3999 (
            .O(N__17134),
            .I(N__17131));
    Odrv4 I__3998 (
            .O(N__17131),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    SRMux I__3997 (
            .O(N__17128),
            .I(N__17123));
    SRMux I__3996 (
            .O(N__17127),
            .I(N__17120));
    SRMux I__3995 (
            .O(N__17126),
            .I(N__17117));
    LocalMux I__3994 (
            .O(N__17123),
            .I(N__17114));
    LocalMux I__3993 (
            .O(N__17120),
            .I(N__17111));
    LocalMux I__3992 (
            .O(N__17117),
            .I(N__17108));
    Span4Mux_h I__3991 (
            .O(N__17114),
            .I(N__17105));
    Span4Mux_h I__3990 (
            .O(N__17111),
            .I(N__17102));
    Span4Mux_h I__3989 (
            .O(N__17108),
            .I(N__17099));
    Span4Mux_h I__3988 (
            .O(N__17105),
            .I(N__17096));
    Span4Mux_h I__3987 (
            .O(N__17102),
            .I(N__17093));
    Span4Mux_h I__3986 (
            .O(N__17099),
            .I(N__17090));
    Span4Mux_v I__3985 (
            .O(N__17096),
            .I(N__17087));
    Odrv4 I__3984 (
            .O(N__17093),
            .I(oneSecStrb_i));
    Odrv4 I__3983 (
            .O(N__17090),
            .I(oneSecStrb_i));
    Odrv4 I__3982 (
            .O(N__17087),
            .I(oneSecStrb_i));
    InMux I__3981 (
            .O(N__17080),
            .I(N__17075));
    InMux I__3980 (
            .O(N__17079),
            .I(N__17068));
    InMux I__3979 (
            .O(N__17078),
            .I(N__17065));
    LocalMux I__3978 (
            .O(N__17075),
            .I(N__17062));
    InMux I__3977 (
            .O(N__17074),
            .I(N__17053));
    InMux I__3976 (
            .O(N__17073),
            .I(N__17053));
    InMux I__3975 (
            .O(N__17072),
            .I(N__17053));
    InMux I__3974 (
            .O(N__17071),
            .I(N__17053));
    LocalMux I__3973 (
            .O(N__17068),
            .I(\Lab_UT.state_1 ));
    LocalMux I__3972 (
            .O(N__17065),
            .I(\Lab_UT.state_1 ));
    Odrv12 I__3971 (
            .O(N__17062),
            .I(\Lab_UT.state_1 ));
    LocalMux I__3970 (
            .O(N__17053),
            .I(\Lab_UT.state_1 ));
    InMux I__3969 (
            .O(N__17044),
            .I(N__17038));
    InMux I__3968 (
            .O(N__17043),
            .I(N__17035));
    InMux I__3967 (
            .O(N__17042),
            .I(N__17032));
    InMux I__3966 (
            .O(N__17041),
            .I(N__17029));
    LocalMux I__3965 (
            .O(N__17038),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_2 ));
    LocalMux I__3964 (
            .O(N__17035),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_2 ));
    LocalMux I__3963 (
            .O(N__17032),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_2 ));
    LocalMux I__3962 (
            .O(N__17029),
            .I(\Lab_UT.dictrl.state_i_3Z0Z_2 ));
    InMux I__3961 (
            .O(N__17020),
            .I(N__17010));
    InMux I__3960 (
            .O(N__17019),
            .I(N__17010));
    CascadeMux I__3959 (
            .O(N__17018),
            .I(N__17005));
    CascadeMux I__3958 (
            .O(N__17017),
            .I(N__17001));
    InMux I__3957 (
            .O(N__17016),
            .I(N__16996));
    InMux I__3956 (
            .O(N__17015),
            .I(N__16996));
    LocalMux I__3955 (
            .O(N__17010),
            .I(N__16993));
    InMux I__3954 (
            .O(N__17009),
            .I(N__16984));
    InMux I__3953 (
            .O(N__17008),
            .I(N__16984));
    InMux I__3952 (
            .O(N__17005),
            .I(N__16984));
    InMux I__3951 (
            .O(N__17004),
            .I(N__16984));
    InMux I__3950 (
            .O(N__17001),
            .I(N__16981));
    LocalMux I__3949 (
            .O(N__16996),
            .I(N__16974));
    Span4Mux_s3_v I__3948 (
            .O(N__16993),
            .I(N__16974));
    LocalMux I__3947 (
            .O(N__16984),
            .I(N__16974));
    LocalMux I__3946 (
            .O(N__16981),
            .I(N__16971));
    Span4Mux_v I__3945 (
            .O(N__16974),
            .I(N__16968));
    Odrv12 I__3944 (
            .O(N__16971),
            .I(\Lab_UT.state_i_3_3 ));
    Odrv4 I__3943 (
            .O(N__16968),
            .I(\Lab_UT.state_i_3_3 ));
    InMux I__3942 (
            .O(N__16963),
            .I(N__16958));
    InMux I__3941 (
            .O(N__16962),
            .I(N__16953));
    InMux I__3940 (
            .O(N__16961),
            .I(N__16953));
    LocalMux I__3939 (
            .O(N__16958),
            .I(N__16950));
    LocalMux I__3938 (
            .O(N__16953),
            .I(N__16947));
    Odrv4 I__3937 (
            .O(N__16950),
            .I(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ));
    Odrv4 I__3936 (
            .O(N__16947),
            .I(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ));
    InMux I__3935 (
            .O(N__16942),
            .I(N__16933));
    InMux I__3934 (
            .O(N__16941),
            .I(N__16933));
    InMux I__3933 (
            .O(N__16940),
            .I(N__16933));
    LocalMux I__3932 (
            .O(N__16933),
            .I(N__16929));
    InMux I__3931 (
            .O(N__16932),
            .I(N__16926));
    Span4Mux_h I__3930 (
            .O(N__16929),
            .I(N__16923));
    LocalMux I__3929 (
            .O(N__16926),
            .I(\Lab_UT.dictrl.state_ret_3_RNIDH8UZ0 ));
    Odrv4 I__3928 (
            .O(N__16923),
            .I(\Lab_UT.dictrl.state_ret_3_RNIDH8UZ0 ));
    CascadeMux I__3927 (
            .O(N__16918),
            .I(N__16915));
    InMux I__3926 (
            .O(N__16915),
            .I(N__16908));
    InMux I__3925 (
            .O(N__16914),
            .I(N__16905));
    CascadeMux I__3924 (
            .O(N__16913),
            .I(N__16902));
    CascadeMux I__3923 (
            .O(N__16912),
            .I(N__16898));
    CascadeMux I__3922 (
            .O(N__16911),
            .I(N__16893));
    LocalMux I__3921 (
            .O(N__16908),
            .I(N__16888));
    LocalMux I__3920 (
            .O(N__16905),
            .I(N__16888));
    InMux I__3919 (
            .O(N__16902),
            .I(N__16881));
    InMux I__3918 (
            .O(N__16901),
            .I(N__16881));
    InMux I__3917 (
            .O(N__16898),
            .I(N__16874));
    InMux I__3916 (
            .O(N__16897),
            .I(N__16874));
    InMux I__3915 (
            .O(N__16896),
            .I(N__16874));
    InMux I__3914 (
            .O(N__16893),
            .I(N__16871));
    Span4Mux_h I__3913 (
            .O(N__16888),
            .I(N__16868));
    CascadeMux I__3912 (
            .O(N__16887),
            .I(N__16864));
    InMux I__3911 (
            .O(N__16886),
            .I(N__16860));
    LocalMux I__3910 (
            .O(N__16881),
            .I(N__16855));
    LocalMux I__3909 (
            .O(N__16874),
            .I(N__16855));
    LocalMux I__3908 (
            .O(N__16871),
            .I(N__16852));
    Span4Mux_s2_v I__3907 (
            .O(N__16868),
            .I(N__16849));
    InMux I__3906 (
            .O(N__16867),
            .I(N__16844));
    InMux I__3905 (
            .O(N__16864),
            .I(N__16844));
    InMux I__3904 (
            .O(N__16863),
            .I(N__16841));
    LocalMux I__3903 (
            .O(N__16860),
            .I(N__16838));
    Span4Mux_v I__3902 (
            .O(N__16855),
            .I(N__16835));
    Sp12to4 I__3901 (
            .O(N__16852),
            .I(N__16826));
    Sp12to4 I__3900 (
            .O(N__16849),
            .I(N__16826));
    LocalMux I__3899 (
            .O(N__16844),
            .I(N__16826));
    LocalMux I__3898 (
            .O(N__16841),
            .I(N__16826));
    Span4Mux_v I__3897 (
            .O(N__16838),
            .I(N__16823));
    Span4Mux_v I__3896 (
            .O(N__16835),
            .I(N__16820));
    Span12Mux_s10_v I__3895 (
            .O(N__16826),
            .I(N__16817));
    Odrv4 I__3894 (
            .O(N__16823),
            .I(\Lab_UT.dictrl.state_retZ0Z_4 ));
    Odrv4 I__3893 (
            .O(N__16820),
            .I(\Lab_UT.dictrl.state_retZ0Z_4 ));
    Odrv12 I__3892 (
            .O(N__16817),
            .I(\Lab_UT.dictrl.state_retZ0Z_4 ));
    InMux I__3891 (
            .O(N__16810),
            .I(N__16807));
    LocalMux I__3890 (
            .O(N__16807),
            .I(N__16802));
    InMux I__3889 (
            .O(N__16806),
            .I(N__16797));
    InMux I__3888 (
            .O(N__16805),
            .I(N__16797));
    Span4Mux_v I__3887 (
            .O(N__16802),
            .I(N__16794));
    LocalMux I__3886 (
            .O(N__16797),
            .I(N__16791));
    Odrv4 I__3885 (
            .O(N__16794),
            .I(\Lab_UT.dictrl.next_state_set ));
    Odrv4 I__3884 (
            .O(N__16791),
            .I(\Lab_UT.dictrl.next_state_set ));
    InMux I__3883 (
            .O(N__16786),
            .I(N__16773));
    InMux I__3882 (
            .O(N__16785),
            .I(N__16773));
    InMux I__3881 (
            .O(N__16784),
            .I(N__16773));
    InMux I__3880 (
            .O(N__16783),
            .I(N__16769));
    InMux I__3879 (
            .O(N__16782),
            .I(N__16762));
    InMux I__3878 (
            .O(N__16781),
            .I(N__16762));
    InMux I__3877 (
            .O(N__16780),
            .I(N__16762));
    LocalMux I__3876 (
            .O(N__16773),
            .I(N__16756));
    InMux I__3875 (
            .O(N__16772),
            .I(N__16752));
    LocalMux I__3874 (
            .O(N__16769),
            .I(N__16747));
    LocalMux I__3873 (
            .O(N__16762),
            .I(N__16747));
    InMux I__3872 (
            .O(N__16761),
            .I(N__16740));
    InMux I__3871 (
            .O(N__16760),
            .I(N__16740));
    InMux I__3870 (
            .O(N__16759),
            .I(N__16740));
    Span4Mux_h I__3869 (
            .O(N__16756),
            .I(N__16737));
    InMux I__3868 (
            .O(N__16755),
            .I(N__16734));
    LocalMux I__3867 (
            .O(N__16752),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__3866 (
            .O(N__16747),
            .I(\Lab_UT.state_0 ));
    LocalMux I__3865 (
            .O(N__16740),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__3864 (
            .O(N__16737),
            .I(\Lab_UT.state_0 ));
    LocalMux I__3863 (
            .O(N__16734),
            .I(\Lab_UT.state_0 ));
    CascadeMux I__3862 (
            .O(N__16723),
            .I(N__16720));
    InMux I__3861 (
            .O(N__16720),
            .I(N__16717));
    LocalMux I__3860 (
            .O(N__16717),
            .I(N__16714));
    Odrv4 I__3859 (
            .O(N__16714),
            .I(\Lab_UT.alarmcharZ0Z_4 ));
    InMux I__3858 (
            .O(N__16711),
            .I(N__16705));
    InMux I__3857 (
            .O(N__16710),
            .I(N__16705));
    LocalMux I__3856 (
            .O(N__16705),
            .I(\Lab_UT.N_204 ));
    CascadeMux I__3855 (
            .O(N__16702),
            .I(\Lab_UT.N_204_cascade_ ));
    InMux I__3854 (
            .O(N__16699),
            .I(N__16687));
    InMux I__3853 (
            .O(N__16698),
            .I(N__16687));
    InMux I__3852 (
            .O(N__16697),
            .I(N__16687));
    InMux I__3851 (
            .O(N__16696),
            .I(N__16687));
    LocalMux I__3850 (
            .O(N__16687),
            .I(N__16684));
    Odrv4 I__3849 (
            .O(N__16684),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__3848 (
            .O(N__16681),
            .I(N__16675));
    InMux I__3847 (
            .O(N__16680),
            .I(N__16675));
    LocalMux I__3846 (
            .O(N__16675),
            .I(\Lab_UT.nine ));
    CascadeMux I__3845 (
            .O(N__16672),
            .I(N__16668));
    CascadeMux I__3844 (
            .O(N__16671),
            .I(N__16664));
    InMux I__3843 (
            .O(N__16668),
            .I(N__16658));
    InMux I__3842 (
            .O(N__16667),
            .I(N__16658));
    InMux I__3841 (
            .O(N__16664),
            .I(N__16653));
    InMux I__3840 (
            .O(N__16663),
            .I(N__16653));
    LocalMux I__3839 (
            .O(N__16658),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    LocalMux I__3838 (
            .O(N__16653),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    CascadeMux I__3837 (
            .O(N__16648),
            .I(N__16640));
    CascadeMux I__3836 (
            .O(N__16647),
            .I(N__16637));
    InMux I__3835 (
            .O(N__16646),
            .I(N__16633));
    InMux I__3834 (
            .O(N__16645),
            .I(N__16626));
    InMux I__3833 (
            .O(N__16644),
            .I(N__16626));
    InMux I__3832 (
            .O(N__16643),
            .I(N__16626));
    InMux I__3831 (
            .O(N__16640),
            .I(N__16619));
    InMux I__3830 (
            .O(N__16637),
            .I(N__16619));
    InMux I__3829 (
            .O(N__16636),
            .I(N__16619));
    LocalMux I__3828 (
            .O(N__16633),
            .I(N__16614));
    LocalMux I__3827 (
            .O(N__16626),
            .I(N__16606));
    LocalMux I__3826 (
            .O(N__16619),
            .I(N__16606));
    InMux I__3825 (
            .O(N__16618),
            .I(N__16603));
    InMux I__3824 (
            .O(N__16617),
            .I(N__16600));
    Span4Mux_v I__3823 (
            .O(N__16614),
            .I(N__16597));
    InMux I__3822 (
            .O(N__16613),
            .I(N__16590));
    InMux I__3821 (
            .O(N__16612),
            .I(N__16590));
    InMux I__3820 (
            .O(N__16611),
            .I(N__16590));
    Span4Mux_v I__3819 (
            .O(N__16606),
            .I(N__16587));
    LocalMux I__3818 (
            .O(N__16603),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3817 (
            .O(N__16600),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__3816 (
            .O(N__16597),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3815 (
            .O(N__16590),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__3814 (
            .O(N__16587),
            .I(\Lab_UT.di_Sones_2 ));
    InMux I__3813 (
            .O(N__16576),
            .I(N__16570));
    InMux I__3812 (
            .O(N__16575),
            .I(N__16559));
    InMux I__3811 (
            .O(N__16574),
            .I(N__16559));
    InMux I__3810 (
            .O(N__16573),
            .I(N__16559));
    LocalMux I__3809 (
            .O(N__16570),
            .I(N__16555));
    CascadeMux I__3808 (
            .O(N__16569),
            .I(N__16550));
    InMux I__3807 (
            .O(N__16568),
            .I(N__16541));
    InMux I__3806 (
            .O(N__16567),
            .I(N__16541));
    InMux I__3805 (
            .O(N__16566),
            .I(N__16541));
    LocalMux I__3804 (
            .O(N__16559),
            .I(N__16538));
    InMux I__3803 (
            .O(N__16558),
            .I(N__16535));
    Span4Mux_s3_h I__3802 (
            .O(N__16555),
            .I(N__16532));
    InMux I__3801 (
            .O(N__16554),
            .I(N__16527));
    InMux I__3800 (
            .O(N__16553),
            .I(N__16527));
    InMux I__3799 (
            .O(N__16550),
            .I(N__16520));
    InMux I__3798 (
            .O(N__16549),
            .I(N__16520));
    InMux I__3797 (
            .O(N__16548),
            .I(N__16520));
    LocalMux I__3796 (
            .O(N__16541),
            .I(N__16515));
    Span12Mux_s9_v I__3795 (
            .O(N__16538),
            .I(N__16515));
    LocalMux I__3794 (
            .O(N__16535),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3793 (
            .O(N__16532),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3792 (
            .O(N__16527),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3791 (
            .O(N__16520),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv12 I__3790 (
            .O(N__16515),
            .I(\Lab_UT.di_Sones_1 ));
    CascadeMux I__3789 (
            .O(N__16504),
            .I(N__16496));
    CascadeMux I__3788 (
            .O(N__16503),
            .I(N__16493));
    CascadeMux I__3787 (
            .O(N__16502),
            .I(N__16490));
    InMux I__3786 (
            .O(N__16501),
            .I(N__16483));
    InMux I__3785 (
            .O(N__16500),
            .I(N__16483));
    InMux I__3784 (
            .O(N__16499),
            .I(N__16483));
    InMux I__3783 (
            .O(N__16496),
            .I(N__16474));
    InMux I__3782 (
            .O(N__16493),
            .I(N__16474));
    InMux I__3781 (
            .O(N__16490),
            .I(N__16474));
    LocalMux I__3780 (
            .O(N__16483),
            .I(N__16471));
    CascadeMux I__3779 (
            .O(N__16482),
            .I(N__16468));
    InMux I__3778 (
            .O(N__16481),
            .I(N__16462));
    LocalMux I__3777 (
            .O(N__16474),
            .I(N__16454));
    Span4Mux_v I__3776 (
            .O(N__16471),
            .I(N__16454));
    InMux I__3775 (
            .O(N__16468),
            .I(N__16451));
    InMux I__3774 (
            .O(N__16467),
            .I(N__16444));
    InMux I__3773 (
            .O(N__16466),
            .I(N__16444));
    InMux I__3772 (
            .O(N__16465),
            .I(N__16444));
    LocalMux I__3771 (
            .O(N__16462),
            .I(N__16441));
    InMux I__3770 (
            .O(N__16461),
            .I(N__16434));
    InMux I__3769 (
            .O(N__16460),
            .I(N__16434));
    InMux I__3768 (
            .O(N__16459),
            .I(N__16434));
    Span4Mux_h I__3767 (
            .O(N__16454),
            .I(N__16431));
    LocalMux I__3766 (
            .O(N__16451),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3765 (
            .O(N__16444),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv12 I__3764 (
            .O(N__16441),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__3763 (
            .O(N__16434),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__3762 (
            .O(N__16431),
            .I(\Lab_UT.di_Sones_0 ));
    CascadeMux I__3761 (
            .O(N__16420),
            .I(N__16414));
    InMux I__3760 (
            .O(N__16419),
            .I(N__16411));
    InMux I__3759 (
            .O(N__16418),
            .I(N__16399));
    InMux I__3758 (
            .O(N__16417),
            .I(N__16399));
    InMux I__3757 (
            .O(N__16414),
            .I(N__16399));
    LocalMux I__3756 (
            .O(N__16411),
            .I(N__16394));
    InMux I__3755 (
            .O(N__16410),
            .I(N__16387));
    InMux I__3754 (
            .O(N__16409),
            .I(N__16387));
    InMux I__3753 (
            .O(N__16408),
            .I(N__16387));
    CascadeMux I__3752 (
            .O(N__16407),
            .I(N__16384));
    CascadeMux I__3751 (
            .O(N__16406),
            .I(N__16381));
    LocalMux I__3750 (
            .O(N__16399),
            .I(N__16378));
    InMux I__3749 (
            .O(N__16398),
            .I(N__16375));
    InMux I__3748 (
            .O(N__16397),
            .I(N__16372));
    Span12Mux_s9_v I__3747 (
            .O(N__16394),
            .I(N__16367));
    LocalMux I__3746 (
            .O(N__16387),
            .I(N__16367));
    InMux I__3745 (
            .O(N__16384),
            .I(N__16362));
    InMux I__3744 (
            .O(N__16381),
            .I(N__16362));
    Span4Mux_h I__3743 (
            .O(N__16378),
            .I(N__16359));
    LocalMux I__3742 (
            .O(N__16375),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3741 (
            .O(N__16372),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv12 I__3740 (
            .O(N__16367),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__3739 (
            .O(N__16362),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv4 I__3738 (
            .O(N__16359),
            .I(\Lab_UT.di_Sones_3 ));
    InMux I__3737 (
            .O(N__16348),
            .I(N__16345));
    LocalMux I__3736 (
            .O(N__16345),
            .I(N__16342));
    Span4Mux_h I__3735 (
            .O(N__16342),
            .I(N__16336));
    InMux I__3734 (
            .O(N__16341),
            .I(N__16333));
    InMux I__3733 (
            .O(N__16340),
            .I(N__16328));
    InMux I__3732 (
            .O(N__16339),
            .I(N__16328));
    Odrv4 I__3731 (
            .O(N__16336),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    LocalMux I__3730 (
            .O(N__16333),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    LocalMux I__3729 (
            .O(N__16328),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__3728 (
            .O(N__16321),
            .I(N__16314));
    InMux I__3727 (
            .O(N__16320),
            .I(N__16314));
    CascadeMux I__3726 (
            .O(N__16319),
            .I(N__16305));
    LocalMux I__3725 (
            .O(N__16314),
            .I(N__16302));
    InMux I__3724 (
            .O(N__16313),
            .I(N__16297));
    InMux I__3723 (
            .O(N__16312),
            .I(N__16297));
    CascadeMux I__3722 (
            .O(N__16311),
            .I(N__16293));
    CascadeMux I__3721 (
            .O(N__16310),
            .I(N__16288));
    CascadeMux I__3720 (
            .O(N__16309),
            .I(N__16285));
    InMux I__3719 (
            .O(N__16308),
            .I(N__16280));
    InMux I__3718 (
            .O(N__16305),
            .I(N__16280));
    Span4Mux_v I__3717 (
            .O(N__16302),
            .I(N__16275));
    LocalMux I__3716 (
            .O(N__16297),
            .I(N__16275));
    InMux I__3715 (
            .O(N__16296),
            .I(N__16262));
    InMux I__3714 (
            .O(N__16293),
            .I(N__16262));
    InMux I__3713 (
            .O(N__16292),
            .I(N__16262));
    InMux I__3712 (
            .O(N__16291),
            .I(N__16262));
    InMux I__3711 (
            .O(N__16288),
            .I(N__16262));
    InMux I__3710 (
            .O(N__16285),
            .I(N__16262));
    LocalMux I__3709 (
            .O(N__16280),
            .I(\Lab_UT.di_Stens_1 ));
    Odrv4 I__3708 (
            .O(N__16275),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__3707 (
            .O(N__16262),
            .I(\Lab_UT.di_Stens_1 ));
    CascadeMux I__3706 (
            .O(N__16255),
            .I(N__16252));
    InMux I__3705 (
            .O(N__16252),
            .I(N__16247));
    CascadeMux I__3704 (
            .O(N__16251),
            .I(N__16244));
    InMux I__3703 (
            .O(N__16250),
            .I(N__16240));
    LocalMux I__3702 (
            .O(N__16247),
            .I(N__16236));
    InMux I__3701 (
            .O(N__16244),
            .I(N__16231));
    InMux I__3700 (
            .O(N__16243),
            .I(N__16231));
    LocalMux I__3699 (
            .O(N__16240),
            .I(N__16226));
    InMux I__3698 (
            .O(N__16239),
            .I(N__16217));
    Span4Mux_v I__3697 (
            .O(N__16236),
            .I(N__16212));
    LocalMux I__3696 (
            .O(N__16231),
            .I(N__16212));
    InMux I__3695 (
            .O(N__16230),
            .I(N__16207));
    InMux I__3694 (
            .O(N__16229),
            .I(N__16207));
    Span4Mux_s3_h I__3693 (
            .O(N__16226),
            .I(N__16204));
    InMux I__3692 (
            .O(N__16225),
            .I(N__16191));
    InMux I__3691 (
            .O(N__16224),
            .I(N__16191));
    InMux I__3690 (
            .O(N__16223),
            .I(N__16191));
    InMux I__3689 (
            .O(N__16222),
            .I(N__16191));
    InMux I__3688 (
            .O(N__16221),
            .I(N__16191));
    InMux I__3687 (
            .O(N__16220),
            .I(N__16191));
    LocalMux I__3686 (
            .O(N__16217),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv4 I__3685 (
            .O(N__16212),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__3684 (
            .O(N__16207),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv4 I__3683 (
            .O(N__16204),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__3682 (
            .O(N__16191),
            .I(\Lab_UT.di_Stens_0 ));
    InMux I__3681 (
            .O(N__16180),
            .I(N__16177));
    LocalMux I__3680 (
            .O(N__16177),
            .I(\Lab_UT.didp.countrce2.three_2 ));
    InMux I__3679 (
            .O(N__16174),
            .I(N__16168));
    CascadeMux I__3678 (
            .O(N__16173),
            .I(N__16165));
    CascadeMux I__3677 (
            .O(N__16172),
            .I(N__16157));
    InMux I__3676 (
            .O(N__16171),
            .I(N__16152));
    LocalMux I__3675 (
            .O(N__16168),
            .I(N__16149));
    InMux I__3674 (
            .O(N__16165),
            .I(N__16146));
    CascadeMux I__3673 (
            .O(N__16164),
            .I(N__16142));
    CascadeMux I__3672 (
            .O(N__16163),
            .I(N__16139));
    InMux I__3671 (
            .O(N__16162),
            .I(N__16134));
    InMux I__3670 (
            .O(N__16161),
            .I(N__16131));
    InMux I__3669 (
            .O(N__16160),
            .I(N__16126));
    InMux I__3668 (
            .O(N__16157),
            .I(N__16126));
    InMux I__3667 (
            .O(N__16156),
            .I(N__16121));
    InMux I__3666 (
            .O(N__16155),
            .I(N__16121));
    LocalMux I__3665 (
            .O(N__16152),
            .I(N__16114));
    Span4Mux_v I__3664 (
            .O(N__16149),
            .I(N__16114));
    LocalMux I__3663 (
            .O(N__16146),
            .I(N__16114));
    InMux I__3662 (
            .O(N__16145),
            .I(N__16103));
    InMux I__3661 (
            .O(N__16142),
            .I(N__16103));
    InMux I__3660 (
            .O(N__16139),
            .I(N__16103));
    InMux I__3659 (
            .O(N__16138),
            .I(N__16103));
    InMux I__3658 (
            .O(N__16137),
            .I(N__16103));
    LocalMux I__3657 (
            .O(N__16134),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__3656 (
            .O(N__16131),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__3655 (
            .O(N__16126),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__3654 (
            .O(N__16121),
            .I(\Lab_UT.di_Stens_2 ));
    Odrv4 I__3653 (
            .O(N__16114),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__3652 (
            .O(N__16103),
            .I(\Lab_UT.di_Stens_2 ));
    CascadeMux I__3651 (
            .O(N__16090),
            .I(\Lab_UT.didp.countrce2.three_2_cascade_ ));
    InMux I__3650 (
            .O(N__16087),
            .I(N__16084));
    LocalMux I__3649 (
            .O(N__16084),
            .I(\Lab_UT.didp.countrce2.un20_qPone ));
    CascadeMux I__3648 (
            .O(N__16081),
            .I(N__16075));
    CascadeMux I__3647 (
            .O(N__16080),
            .I(N__16072));
    InMux I__3646 (
            .O(N__16079),
            .I(N__16064));
    InMux I__3645 (
            .O(N__16078),
            .I(N__16064));
    InMux I__3644 (
            .O(N__16075),
            .I(N__16059));
    InMux I__3643 (
            .O(N__16072),
            .I(N__16059));
    CascadeMux I__3642 (
            .O(N__16071),
            .I(N__16056));
    CascadeMux I__3641 (
            .O(N__16070),
            .I(N__16053));
    CascadeMux I__3640 (
            .O(N__16069),
            .I(N__16050));
    LocalMux I__3639 (
            .O(N__16064),
            .I(N__16044));
    LocalMux I__3638 (
            .O(N__16059),
            .I(N__16041));
    InMux I__3637 (
            .O(N__16056),
            .I(N__16032));
    InMux I__3636 (
            .O(N__16053),
            .I(N__16032));
    InMux I__3635 (
            .O(N__16050),
            .I(N__16032));
    InMux I__3634 (
            .O(N__16049),
            .I(N__16032));
    InMux I__3633 (
            .O(N__16048),
            .I(N__16028));
    CascadeMux I__3632 (
            .O(N__16047),
            .I(N__16022));
    Span4Mux_v I__3631 (
            .O(N__16044),
            .I(N__16015));
    Span4Mux_h I__3630 (
            .O(N__16041),
            .I(N__16015));
    LocalMux I__3629 (
            .O(N__16032),
            .I(N__16015));
    InMux I__3628 (
            .O(N__16031),
            .I(N__16012));
    LocalMux I__3627 (
            .O(N__16028),
            .I(N__16009));
    InMux I__3626 (
            .O(N__16027),
            .I(N__16006));
    InMux I__3625 (
            .O(N__16026),
            .I(N__15999));
    InMux I__3624 (
            .O(N__16025),
            .I(N__15999));
    InMux I__3623 (
            .O(N__16022),
            .I(N__15999));
    Span4Mux_h I__3622 (
            .O(N__16015),
            .I(N__15996));
    LocalMux I__3621 (
            .O(N__16012),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__3620 (
            .O(N__16009),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3619 (
            .O(N__16006),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3618 (
            .O(N__15999),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv4 I__3617 (
            .O(N__15996),
            .I(\Lab_UT.di_Mones_3 ));
    CascadeMux I__3616 (
            .O(N__15985),
            .I(N__15974));
    InMux I__3615 (
            .O(N__15984),
            .I(N__15969));
    InMux I__3614 (
            .O(N__15983),
            .I(N__15969));
    InMux I__3613 (
            .O(N__15982),
            .I(N__15963));
    InMux I__3612 (
            .O(N__15981),
            .I(N__15963));
    InMux I__3611 (
            .O(N__15980),
            .I(N__15954));
    InMux I__3610 (
            .O(N__15979),
            .I(N__15954));
    InMux I__3609 (
            .O(N__15978),
            .I(N__15954));
    InMux I__3608 (
            .O(N__15977),
            .I(N__15954));
    InMux I__3607 (
            .O(N__15974),
            .I(N__15950));
    LocalMux I__3606 (
            .O(N__15969),
            .I(N__15947));
    InMux I__3605 (
            .O(N__15968),
            .I(N__15940));
    LocalMux I__3604 (
            .O(N__15963),
            .I(N__15937));
    LocalMux I__3603 (
            .O(N__15954),
            .I(N__15934));
    InMux I__3602 (
            .O(N__15953),
            .I(N__15931));
    LocalMux I__3601 (
            .O(N__15950),
            .I(N__15928));
    Span4Mux_v I__3600 (
            .O(N__15947),
            .I(N__15925));
    InMux I__3599 (
            .O(N__15946),
            .I(N__15916));
    InMux I__3598 (
            .O(N__15945),
            .I(N__15916));
    InMux I__3597 (
            .O(N__15944),
            .I(N__15916));
    InMux I__3596 (
            .O(N__15943),
            .I(N__15916));
    LocalMux I__3595 (
            .O(N__15940),
            .I(N__15909));
    Span4Mux_h I__3594 (
            .O(N__15937),
            .I(N__15909));
    Span4Mux_h I__3593 (
            .O(N__15934),
            .I(N__15909));
    LocalMux I__3592 (
            .O(N__15931),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv12 I__3591 (
            .O(N__15928),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3590 (
            .O(N__15925),
            .I(\Lab_UT.di_Mones_2 ));
    LocalMux I__3589 (
            .O(N__15916),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3588 (
            .O(N__15909),
            .I(\Lab_UT.di_Mones_2 ));
    InMux I__3587 (
            .O(N__15898),
            .I(N__15895));
    LocalMux I__3586 (
            .O(N__15895),
            .I(N__15891));
    InMux I__3585 (
            .O(N__15894),
            .I(N__15888));
    Span4Mux_h I__3584 (
            .O(N__15891),
            .I(N__15885));
    LocalMux I__3583 (
            .O(N__15888),
            .I(\Lab_UT.N_207 ));
    Odrv4 I__3582 (
            .O(N__15885),
            .I(\Lab_UT.N_207 ));
    CascadeMux I__3581 (
            .O(N__15880),
            .I(N__15876));
    InMux I__3580 (
            .O(N__15879),
            .I(N__15872));
    InMux I__3579 (
            .O(N__15876),
            .I(N__15867));
    InMux I__3578 (
            .O(N__15875),
            .I(N__15867));
    LocalMux I__3577 (
            .O(N__15872),
            .I(N__15864));
    LocalMux I__3576 (
            .O(N__15867),
            .I(\Lab_UT.didp.q_RNI84NN1_3 ));
    Odrv4 I__3575 (
            .O(N__15864),
            .I(\Lab_UT.didp.q_RNI84NN1_3 ));
    CascadeMux I__3574 (
            .O(N__15859),
            .I(N__15856));
    InMux I__3573 (
            .O(N__15856),
            .I(N__15852));
    CascadeMux I__3572 (
            .O(N__15855),
            .I(N__15848));
    LocalMux I__3571 (
            .O(N__15852),
            .I(N__15844));
    InMux I__3570 (
            .O(N__15851),
            .I(N__15837));
    InMux I__3569 (
            .O(N__15848),
            .I(N__15837));
    InMux I__3568 (
            .O(N__15847),
            .I(N__15837));
    Odrv4 I__3567 (
            .O(N__15844),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    LocalMux I__3566 (
            .O(N__15837),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    InMux I__3565 (
            .O(N__15832),
            .I(N__15829));
    LocalMux I__3564 (
            .O(N__15829),
            .I(N__15826));
    Odrv4 I__3563 (
            .O(N__15826),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_3 ));
    CascadeMux I__3562 (
            .O(N__15823),
            .I(N__15815));
    InMux I__3561 (
            .O(N__15822),
            .I(N__15808));
    InMux I__3560 (
            .O(N__15821),
            .I(N__15808));
    InMux I__3559 (
            .O(N__15820),
            .I(N__15803));
    InMux I__3558 (
            .O(N__15819),
            .I(N__15803));
    InMux I__3557 (
            .O(N__15818),
            .I(N__15796));
    InMux I__3556 (
            .O(N__15815),
            .I(N__15796));
    InMux I__3555 (
            .O(N__15814),
            .I(N__15796));
    InMux I__3554 (
            .O(N__15813),
            .I(N__15791));
    LocalMux I__3553 (
            .O(N__15808),
            .I(N__15788));
    LocalMux I__3552 (
            .O(N__15803),
            .I(N__15785));
    LocalMux I__3551 (
            .O(N__15796),
            .I(N__15782));
    CascadeMux I__3550 (
            .O(N__15795),
            .I(N__15779));
    CascadeMux I__3549 (
            .O(N__15794),
            .I(N__15775));
    LocalMux I__3548 (
            .O(N__15791),
            .I(N__15770));
    Span4Mux_v I__3547 (
            .O(N__15788),
            .I(N__15767));
    Span4Mux_h I__3546 (
            .O(N__15785),
            .I(N__15762));
    Span4Mux_h I__3545 (
            .O(N__15782),
            .I(N__15762));
    InMux I__3544 (
            .O(N__15779),
            .I(N__15753));
    InMux I__3543 (
            .O(N__15778),
            .I(N__15753));
    InMux I__3542 (
            .O(N__15775),
            .I(N__15753));
    InMux I__3541 (
            .O(N__15774),
            .I(N__15753));
    InMux I__3540 (
            .O(N__15773),
            .I(N__15750));
    Odrv4 I__3539 (
            .O(N__15770),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv4 I__3538 (
            .O(N__15767),
            .I(\Lab_UT.di_Mones_1 ));
    Odrv4 I__3537 (
            .O(N__15762),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3536 (
            .O(N__15753),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3535 (
            .O(N__15750),
            .I(\Lab_UT.di_Mones_1 ));
    CascadeMux I__3534 (
            .O(N__15739),
            .I(N__15735));
    CascadeMux I__3533 (
            .O(N__15738),
            .I(N__15732));
    InMux I__3532 (
            .O(N__15735),
            .I(N__15721));
    InMux I__3531 (
            .O(N__15732),
            .I(N__15721));
    InMux I__3530 (
            .O(N__15731),
            .I(N__15716));
    InMux I__3529 (
            .O(N__15730),
            .I(N__15716));
    InMux I__3528 (
            .O(N__15729),
            .I(N__15709));
    InMux I__3527 (
            .O(N__15728),
            .I(N__15709));
    InMux I__3526 (
            .O(N__15727),
            .I(N__15709));
    InMux I__3525 (
            .O(N__15726),
            .I(N__15706));
    LocalMux I__3524 (
            .O(N__15721),
            .I(N__15703));
    LocalMux I__3523 (
            .O(N__15716),
            .I(N__15693));
    LocalMux I__3522 (
            .O(N__15709),
            .I(N__15693));
    LocalMux I__3521 (
            .O(N__15706),
            .I(N__15689));
    Span4Mux_h I__3520 (
            .O(N__15703),
            .I(N__15686));
    InMux I__3519 (
            .O(N__15702),
            .I(N__15675));
    InMux I__3518 (
            .O(N__15701),
            .I(N__15675));
    InMux I__3517 (
            .O(N__15700),
            .I(N__15675));
    InMux I__3516 (
            .O(N__15699),
            .I(N__15675));
    InMux I__3515 (
            .O(N__15698),
            .I(N__15675));
    Span4Mux_h I__3514 (
            .O(N__15693),
            .I(N__15672));
    InMux I__3513 (
            .O(N__15692),
            .I(N__15669));
    Odrv4 I__3512 (
            .O(N__15689),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__3511 (
            .O(N__15686),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__3510 (
            .O(N__15675),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__3509 (
            .O(N__15672),
            .I(\Lab_UT.di_Mones_0 ));
    LocalMux I__3508 (
            .O(N__15669),
            .I(\Lab_UT.di_Mones_0 ));
    CascadeMux I__3507 (
            .O(N__15658),
            .I(\Lab_UT.N_207_cascade_ ));
    CascadeMux I__3506 (
            .O(N__15655),
            .I(N__15652));
    InMux I__3505 (
            .O(N__15652),
            .I(N__15646));
    InMux I__3504 (
            .O(N__15651),
            .I(N__15646));
    LocalMux I__3503 (
            .O(N__15646),
            .I(N__15643));
    Odrv4 I__3502 (
            .O(N__15643),
            .I(\Lab_UT.didp.q_RNIIKFH3_3 ));
    CascadeMux I__3501 (
            .O(N__15640),
            .I(N__15635));
    InMux I__3500 (
            .O(N__15639),
            .I(N__15632));
    InMux I__3499 (
            .O(N__15638),
            .I(N__15629));
    InMux I__3498 (
            .O(N__15635),
            .I(N__15626));
    LocalMux I__3497 (
            .O(N__15632),
            .I(N__15623));
    LocalMux I__3496 (
            .O(N__15629),
            .I(N__15619));
    LocalMux I__3495 (
            .O(N__15626),
            .I(N__15614));
    Span4Mux_h I__3494 (
            .O(N__15623),
            .I(N__15614));
    InMux I__3493 (
            .O(N__15622),
            .I(N__15611));
    Odrv4 I__3492 (
            .O(N__15619),
            .I(\Lab_UT.m40 ));
    Odrv4 I__3491 (
            .O(N__15614),
            .I(\Lab_UT.m40 ));
    LocalMux I__3490 (
            .O(N__15611),
            .I(\Lab_UT.m40 ));
    CascadeMux I__3489 (
            .O(N__15604),
            .I(N__15601));
    InMux I__3488 (
            .O(N__15601),
            .I(N__15597));
    CascadeMux I__3487 (
            .O(N__15600),
            .I(N__15594));
    LocalMux I__3486 (
            .O(N__15597),
            .I(N__15590));
    InMux I__3485 (
            .O(N__15594),
            .I(N__15587));
    InMux I__3484 (
            .O(N__15593),
            .I(N__15584));
    Span4Mux_h I__3483 (
            .O(N__15590),
            .I(N__15581));
    LocalMux I__3482 (
            .O(N__15587),
            .I(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3 ));
    LocalMux I__3481 (
            .O(N__15584),
            .I(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3 ));
    Odrv4 I__3480 (
            .O(N__15581),
            .I(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3 ));
    InMux I__3479 (
            .O(N__15574),
            .I(N__15571));
    LocalMux I__3478 (
            .O(N__15571),
            .I(N__15566));
    InMux I__3477 (
            .O(N__15570),
            .I(N__15562));
    InMux I__3476 (
            .O(N__15569),
            .I(N__15559));
    Span4Mux_h I__3475 (
            .O(N__15566),
            .I(N__15556));
    InMux I__3474 (
            .O(N__15565),
            .I(N__15553));
    LocalMux I__3473 (
            .O(N__15562),
            .I(N__15548));
    LocalMux I__3472 (
            .O(N__15559),
            .I(N__15548));
    Odrv4 I__3471 (
            .O(N__15556),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    LocalMux I__3470 (
            .O(N__15553),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    Odrv4 I__3469 (
            .O(N__15548),
            .I(\Lab_UT.dictrl.next_state_set_2 ));
    InMux I__3468 (
            .O(N__15541),
            .I(N__15538));
    LocalMux I__3467 (
            .O(N__15538),
            .I(N__15535));
    Odrv4 I__3466 (
            .O(N__15535),
            .I(\Lab_UT.alarmcharZ0Z_2 ));
    CascadeMux I__3465 (
            .O(N__15532),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_2_cascade_ ));
    CascadeMux I__3464 (
            .O(N__15529),
            .I(N__15522));
    CascadeMux I__3463 (
            .O(N__15528),
            .I(N__15519));
    CascadeMux I__3462 (
            .O(N__15527),
            .I(N__15516));
    CascadeMux I__3461 (
            .O(N__15526),
            .I(N__15513));
    InMux I__3460 (
            .O(N__15525),
            .I(N__15508));
    InMux I__3459 (
            .O(N__15522),
            .I(N__15503));
    InMux I__3458 (
            .O(N__15519),
            .I(N__15503));
    InMux I__3457 (
            .O(N__15516),
            .I(N__15498));
    InMux I__3456 (
            .O(N__15513),
            .I(N__15498));
    InMux I__3455 (
            .O(N__15512),
            .I(N__15495));
    CascadeMux I__3454 (
            .O(N__15511),
            .I(N__15491));
    LocalMux I__3453 (
            .O(N__15508),
            .I(N__15483));
    LocalMux I__3452 (
            .O(N__15503),
            .I(N__15480));
    LocalMux I__3451 (
            .O(N__15498),
            .I(N__15477));
    LocalMux I__3450 (
            .O(N__15495),
            .I(N__15474));
    InMux I__3449 (
            .O(N__15494),
            .I(N__15469));
    InMux I__3448 (
            .O(N__15491),
            .I(N__15469));
    CascadeMux I__3447 (
            .O(N__15490),
            .I(N__15466));
    InMux I__3446 (
            .O(N__15489),
            .I(N__15461));
    InMux I__3445 (
            .O(N__15488),
            .I(N__15461));
    CascadeMux I__3444 (
            .O(N__15487),
            .I(N__15458));
    InMux I__3443 (
            .O(N__15486),
            .I(N__15455));
    Span4Mux_h I__3442 (
            .O(N__15483),
            .I(N__15450));
    Span4Mux_v I__3441 (
            .O(N__15480),
            .I(N__15450));
    Span4Mux_v I__3440 (
            .O(N__15477),
            .I(N__15443));
    Span4Mux_v I__3439 (
            .O(N__15474),
            .I(N__15443));
    LocalMux I__3438 (
            .O(N__15469),
            .I(N__15443));
    InMux I__3437 (
            .O(N__15466),
            .I(N__15440));
    LocalMux I__3436 (
            .O(N__15461),
            .I(N__15437));
    InMux I__3435 (
            .O(N__15458),
            .I(N__15434));
    LocalMux I__3434 (
            .O(N__15455),
            .I(N__15429));
    Span4Mux_v I__3433 (
            .O(N__15450),
            .I(N__15429));
    Span4Mux_h I__3432 (
            .O(N__15443),
            .I(N__15426));
    LocalMux I__3431 (
            .O(N__15440),
            .I(N__15423));
    Odrv12 I__3430 (
            .O(N__15437),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3429 (
            .O(N__15434),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__3428 (
            .O(N__15429),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__3427 (
            .O(N__15426),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv12 I__3426 (
            .O(N__15423),
            .I(\Lab_UT.di_Mtens_2 ));
    InMux I__3425 (
            .O(N__15412),
            .I(N__15409));
    LocalMux I__3424 (
            .O(N__15409),
            .I(N__15406));
    Odrv12 I__3423 (
            .O(N__15406),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_2 ));
    InMux I__3422 (
            .O(N__15403),
            .I(N__15394));
    InMux I__3421 (
            .O(N__15402),
            .I(N__15394));
    InMux I__3420 (
            .O(N__15401),
            .I(N__15394));
    LocalMux I__3419 (
            .O(N__15394),
            .I(N__15390));
    InMux I__3418 (
            .O(N__15393),
            .I(N__15387));
    Odrv4 I__3417 (
            .O(N__15390),
            .I(\Lab_UT.un3_dOutP ));
    LocalMux I__3416 (
            .O(N__15387),
            .I(\Lab_UT.un3_dOutP ));
    InMux I__3415 (
            .O(N__15382),
            .I(N__15378));
    InMux I__3414 (
            .O(N__15381),
            .I(N__15368));
    LocalMux I__3413 (
            .O(N__15378),
            .I(N__15365));
    InMux I__3412 (
            .O(N__15377),
            .I(N__15362));
    CascadeMux I__3411 (
            .O(N__15376),
            .I(N__15359));
    InMux I__3410 (
            .O(N__15375),
            .I(N__15348));
    InMux I__3409 (
            .O(N__15374),
            .I(N__15348));
    InMux I__3408 (
            .O(N__15373),
            .I(N__15348));
    InMux I__3407 (
            .O(N__15372),
            .I(N__15348));
    InMux I__3406 (
            .O(N__15371),
            .I(N__15348));
    LocalMux I__3405 (
            .O(N__15368),
            .I(N__15341));
    Span4Mux_h I__3404 (
            .O(N__15365),
            .I(N__15341));
    LocalMux I__3403 (
            .O(N__15362),
            .I(N__15341));
    InMux I__3402 (
            .O(N__15359),
            .I(N__15336));
    LocalMux I__3401 (
            .O(N__15348),
            .I(N__15333));
    Span4Mux_v I__3400 (
            .O(N__15341),
            .I(N__15330));
    InMux I__3399 (
            .O(N__15340),
            .I(N__15325));
    InMux I__3398 (
            .O(N__15339),
            .I(N__15325));
    LocalMux I__3397 (
            .O(N__15336),
            .I(\Lab_UT.cnt_3 ));
    Odrv12 I__3396 (
            .O(N__15333),
            .I(\Lab_UT.cnt_3 ));
    Odrv4 I__3395 (
            .O(N__15330),
            .I(\Lab_UT.cnt_3 ));
    LocalMux I__3394 (
            .O(N__15325),
            .I(\Lab_UT.cnt_3 ));
    InMux I__3393 (
            .O(N__15316),
            .I(N__15313));
    LocalMux I__3392 (
            .O(N__15313),
            .I(N__15308));
    InMux I__3391 (
            .O(N__15312),
            .I(N__15303));
    InMux I__3390 (
            .O(N__15311),
            .I(N__15303));
    Span4Mux_v I__3389 (
            .O(N__15308),
            .I(N__15300));
    LocalMux I__3388 (
            .O(N__15303),
            .I(N__15297));
    Sp12to4 I__3387 (
            .O(N__15300),
            .I(N__15294));
    Span4Mux_h I__3386 (
            .O(N__15297),
            .I(N__15291));
    Span12Mux_s6_h I__3385 (
            .O(N__15294),
            .I(N__15286));
    Span4Mux_h I__3384 (
            .O(N__15291),
            .I(N__15283));
    InMux I__3383 (
            .O(N__15290),
            .I(N__15278));
    InMux I__3382 (
            .O(N__15289),
            .I(N__15278));
    Odrv12 I__3381 (
            .O(N__15286),
            .I(\Lab_UT.cnt_0 ));
    Odrv4 I__3380 (
            .O(N__15283),
            .I(\Lab_UT.cnt_0 ));
    LocalMux I__3379 (
            .O(N__15278),
            .I(\Lab_UT.cnt_0 ));
    InMux I__3378 (
            .O(N__15271),
            .I(N__15262));
    InMux I__3377 (
            .O(N__15270),
            .I(N__15251));
    InMux I__3376 (
            .O(N__15269),
            .I(N__15251));
    InMux I__3375 (
            .O(N__15268),
            .I(N__15251));
    InMux I__3374 (
            .O(N__15267),
            .I(N__15251));
    InMux I__3373 (
            .O(N__15266),
            .I(N__15251));
    InMux I__3372 (
            .O(N__15265),
            .I(N__15248));
    LocalMux I__3371 (
            .O(N__15262),
            .I(N__15236));
    LocalMux I__3370 (
            .O(N__15251),
            .I(N__15236));
    LocalMux I__3369 (
            .O(N__15248),
            .I(N__15233));
    InMux I__3368 (
            .O(N__15247),
            .I(N__15224));
    InMux I__3367 (
            .O(N__15246),
            .I(N__15224));
    InMux I__3366 (
            .O(N__15245),
            .I(N__15224));
    InMux I__3365 (
            .O(N__15244),
            .I(N__15224));
    InMux I__3364 (
            .O(N__15243),
            .I(N__15221));
    InMux I__3363 (
            .O(N__15242),
            .I(N__15218));
    InMux I__3362 (
            .O(N__15241),
            .I(N__15215));
    Span4Mux_h I__3361 (
            .O(N__15236),
            .I(N__15212));
    Span4Mux_v I__3360 (
            .O(N__15233),
            .I(N__15207));
    LocalMux I__3359 (
            .O(N__15224),
            .I(N__15207));
    LocalMux I__3358 (
            .O(N__15221),
            .I(N__15199));
    LocalMux I__3357 (
            .O(N__15218),
            .I(N__15199));
    LocalMux I__3356 (
            .O(N__15215),
            .I(N__15199));
    Span4Mux_v I__3355 (
            .O(N__15212),
            .I(N__15194));
    Span4Mux_h I__3354 (
            .O(N__15207),
            .I(N__15194));
    InMux I__3353 (
            .O(N__15206),
            .I(N__15191));
    Span12Mux_s11_h I__3352 (
            .O(N__15199),
            .I(N__15188));
    Span4Mux_h I__3351 (
            .O(N__15194),
            .I(N__15185));
    LocalMux I__3350 (
            .O(N__15191),
            .I(\Lab_UT.cnt_1 ));
    Odrv12 I__3349 (
            .O(N__15188),
            .I(\Lab_UT.cnt_1 ));
    Odrv4 I__3348 (
            .O(N__15185),
            .I(\Lab_UT.cnt_1 ));
    CascadeMux I__3347 (
            .O(N__15178),
            .I(N__15175));
    InMux I__3346 (
            .O(N__15175),
            .I(N__15167));
    InMux I__3345 (
            .O(N__15174),
            .I(N__15164));
    CascadeMux I__3344 (
            .O(N__15173),
            .I(N__15159));
    CascadeMux I__3343 (
            .O(N__15172),
            .I(N__15156));
    InMux I__3342 (
            .O(N__15171),
            .I(N__15152));
    InMux I__3341 (
            .O(N__15170),
            .I(N__15149));
    LocalMux I__3340 (
            .O(N__15167),
            .I(N__15142));
    LocalMux I__3339 (
            .O(N__15164),
            .I(N__15142));
    InMux I__3338 (
            .O(N__15163),
            .I(N__15131));
    InMux I__3337 (
            .O(N__15162),
            .I(N__15131));
    InMux I__3336 (
            .O(N__15159),
            .I(N__15131));
    InMux I__3335 (
            .O(N__15156),
            .I(N__15131));
    InMux I__3334 (
            .O(N__15155),
            .I(N__15131));
    LocalMux I__3333 (
            .O(N__15152),
            .I(N__15126));
    LocalMux I__3332 (
            .O(N__15149),
            .I(N__15126));
    CascadeMux I__3331 (
            .O(N__15148),
            .I(N__15123));
    InMux I__3330 (
            .O(N__15147),
            .I(N__15117));
    Sp12to4 I__3329 (
            .O(N__15142),
            .I(N__15112));
    LocalMux I__3328 (
            .O(N__15131),
            .I(N__15112));
    Span4Mux_h I__3327 (
            .O(N__15126),
            .I(N__15109));
    InMux I__3326 (
            .O(N__15123),
            .I(N__15100));
    InMux I__3325 (
            .O(N__15122),
            .I(N__15100));
    InMux I__3324 (
            .O(N__15121),
            .I(N__15100));
    InMux I__3323 (
            .O(N__15120),
            .I(N__15100));
    LocalMux I__3322 (
            .O(N__15117),
            .I(\Lab_UT.cnt_2 ));
    Odrv12 I__3321 (
            .O(N__15112),
            .I(\Lab_UT.cnt_2 ));
    Odrv4 I__3320 (
            .O(N__15109),
            .I(\Lab_UT.cnt_2 ));
    LocalMux I__3319 (
            .O(N__15100),
            .I(\Lab_UT.cnt_2 ));
    CascadeMux I__3318 (
            .O(N__15091),
            .I(\Lab_UT.alarmchar9_cascade_ ));
    CascadeMux I__3317 (
            .O(N__15088),
            .I(N__15084));
    CascadeMux I__3316 (
            .O(N__15087),
            .I(N__15081));
    InMux I__3315 (
            .O(N__15084),
            .I(N__15076));
    InMux I__3314 (
            .O(N__15081),
            .I(N__15076));
    LocalMux I__3313 (
            .O(N__15076),
            .I(\Lab_UT.alarmcharZ0Z_1 ));
    InMux I__3312 (
            .O(N__15073),
            .I(N__15070));
    LocalMux I__3311 (
            .O(N__15070),
            .I(N__15067));
    Odrv4 I__3310 (
            .O(N__15067),
            .I(\Lab_UT.zero ));
    CascadeMux I__3309 (
            .O(N__15064),
            .I(\Lab_UT.didp.countrce3.qPone_3_cascade_ ));
    CascadeMux I__3308 (
            .O(N__15061),
            .I(\Lab_UT.didp.countrce3.N_79_i_cascade_ ));
    InMux I__3307 (
            .O(N__15058),
            .I(N__15052));
    InMux I__3306 (
            .O(N__15057),
            .I(N__15045));
    InMux I__3305 (
            .O(N__15056),
            .I(N__15045));
    InMux I__3304 (
            .O(N__15055),
            .I(N__15045));
    LocalMux I__3303 (
            .O(N__15052),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    LocalMux I__3302 (
            .O(N__15045),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    CascadeMux I__3301 (
            .O(N__15040),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_0_cascade_ ));
    InMux I__3300 (
            .O(N__15037),
            .I(N__15034));
    LocalMux I__3299 (
            .O(N__15034),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_0 ));
    CascadeMux I__3298 (
            .O(N__15031),
            .I(N__15025));
    CascadeMux I__3297 (
            .O(N__15030),
            .I(N__15022));
    InMux I__3296 (
            .O(N__15029),
            .I(N__15019));
    InMux I__3295 (
            .O(N__15028),
            .I(N__15016));
    InMux I__3294 (
            .O(N__15025),
            .I(N__15011));
    InMux I__3293 (
            .O(N__15022),
            .I(N__15011));
    LocalMux I__3292 (
            .O(N__15019),
            .I(\Lab_UT.un29_dOutP ));
    LocalMux I__3291 (
            .O(N__15016),
            .I(\Lab_UT.un29_dOutP ));
    LocalMux I__3290 (
            .O(N__15011),
            .I(\Lab_UT.un29_dOutP ));
    InMux I__3289 (
            .O(N__15004),
            .I(N__15001));
    LocalMux I__3288 (
            .O(N__15001),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_1 ));
    CascadeMux I__3287 (
            .O(N__14998),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_1_cascade_ ));
    InMux I__3286 (
            .O(N__14995),
            .I(N__14992));
    LocalMux I__3285 (
            .O(N__14992),
            .I(N__14988));
    InMux I__3284 (
            .O(N__14991),
            .I(N__14984));
    Span4Mux_h I__3283 (
            .O(N__14988),
            .I(N__14981));
    InMux I__3282 (
            .O(N__14987),
            .I(N__14978));
    LocalMux I__3281 (
            .O(N__14984),
            .I(N__14973));
    Span4Mux_h I__3280 (
            .O(N__14981),
            .I(N__14970));
    LocalMux I__3279 (
            .O(N__14978),
            .I(N__14967));
    InMux I__3278 (
            .O(N__14977),
            .I(N__14962));
    InMux I__3277 (
            .O(N__14976),
            .I(N__14962));
    Odrv12 I__3276 (
            .O(N__14973),
            .I(L3_tx_data_1));
    Odrv4 I__3275 (
            .O(N__14970),
            .I(L3_tx_data_1));
    Odrv4 I__3274 (
            .O(N__14967),
            .I(L3_tx_data_1));
    LocalMux I__3273 (
            .O(N__14962),
            .I(L3_tx_data_1));
    InMux I__3272 (
            .O(N__14953),
            .I(N__14950));
    LocalMux I__3271 (
            .O(N__14950),
            .I(N__14947));
    Odrv4 I__3270 (
            .O(N__14947),
            .I(\Lab_UT.dispString.dOutP_0_iv_3_1 ));
    InMux I__3269 (
            .O(N__14944),
            .I(N__14938));
    InMux I__3268 (
            .O(N__14943),
            .I(N__14932));
    InMux I__3267 (
            .O(N__14942),
            .I(N__14929));
    InMux I__3266 (
            .O(N__14941),
            .I(N__14926));
    LocalMux I__3265 (
            .O(N__14938),
            .I(N__14923));
    InMux I__3264 (
            .O(N__14937),
            .I(N__14920));
    InMux I__3263 (
            .O(N__14936),
            .I(N__14909));
    InMux I__3262 (
            .O(N__14935),
            .I(N__14909));
    LocalMux I__3261 (
            .O(N__14932),
            .I(N__14906));
    LocalMux I__3260 (
            .O(N__14929),
            .I(N__14903));
    LocalMux I__3259 (
            .O(N__14926),
            .I(N__14896));
    Span4Mux_v I__3258 (
            .O(N__14923),
            .I(N__14896));
    LocalMux I__3257 (
            .O(N__14920),
            .I(N__14896));
    InMux I__3256 (
            .O(N__14919),
            .I(N__14893));
    InMux I__3255 (
            .O(N__14918),
            .I(N__14888));
    InMux I__3254 (
            .O(N__14917),
            .I(N__14888));
    InMux I__3253 (
            .O(N__14916),
            .I(N__14883));
    InMux I__3252 (
            .O(N__14915),
            .I(N__14883));
    InMux I__3251 (
            .O(N__14914),
            .I(N__14879));
    LocalMux I__3250 (
            .O(N__14909),
            .I(N__14874));
    Span4Mux_v I__3249 (
            .O(N__14906),
            .I(N__14874));
    Span4Mux_s3_h I__3248 (
            .O(N__14903),
            .I(N__14867));
    Span4Mux_h I__3247 (
            .O(N__14896),
            .I(N__14867));
    LocalMux I__3246 (
            .O(N__14893),
            .I(N__14867));
    LocalMux I__3245 (
            .O(N__14888),
            .I(N__14862));
    LocalMux I__3244 (
            .O(N__14883),
            .I(N__14862));
    InMux I__3243 (
            .O(N__14882),
            .I(N__14859));
    LocalMux I__3242 (
            .O(N__14879),
            .I(N__14852));
    Span4Mux_h I__3241 (
            .O(N__14874),
            .I(N__14852));
    Span4Mux_v I__3240 (
            .O(N__14867),
            .I(N__14852));
    Odrv4 I__3239 (
            .O(N__14862),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__3238 (
            .O(N__14859),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__3237 (
            .O(N__14852),
            .I(\Lab_UT.di_Mtens_1 ));
    InMux I__3236 (
            .O(N__14845),
            .I(N__14842));
    LocalMux I__3235 (
            .O(N__14842),
            .I(\Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0 ));
    InMux I__3234 (
            .O(N__14839),
            .I(N__14835));
    InMux I__3233 (
            .O(N__14838),
            .I(N__14832));
    LocalMux I__3232 (
            .O(N__14835),
            .I(N__14826));
    LocalMux I__3231 (
            .O(N__14832),
            .I(N__14826));
    InMux I__3230 (
            .O(N__14831),
            .I(N__14823));
    Span4Mux_h I__3229 (
            .O(N__14826),
            .I(N__14820));
    LocalMux I__3228 (
            .O(N__14823),
            .I(\Lab_UT.m24 ));
    Odrv4 I__3227 (
            .O(N__14820),
            .I(\Lab_UT.m24 ));
    InMux I__3226 (
            .O(N__14815),
            .I(N__14809));
    InMux I__3225 (
            .O(N__14814),
            .I(N__14809));
    LocalMux I__3224 (
            .O(N__14809),
            .I(\Lab_UT.dispString.un22_dOutP ));
    InMux I__3223 (
            .O(N__14806),
            .I(N__14803));
    LocalMux I__3222 (
            .O(N__14803),
            .I(N__14800));
    Odrv4 I__3221 (
            .O(N__14800),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_3 ));
    CascadeMux I__3220 (
            .O(N__14797),
            .I(\Lab_UT.dispString.dOutP_0_iv_3_3_cascade_ ));
    InMux I__3219 (
            .O(N__14794),
            .I(N__14791));
    LocalMux I__3218 (
            .O(N__14791),
            .I(N__14787));
    InMux I__3217 (
            .O(N__14790),
            .I(N__14784));
    Span4Mux_h I__3216 (
            .O(N__14787),
            .I(N__14781));
    LocalMux I__3215 (
            .O(N__14784),
            .I(N__14778));
    Span4Mux_h I__3214 (
            .O(N__14781),
            .I(N__14774));
    Span12Mux_s8_h I__3213 (
            .O(N__14778),
            .I(N__14771));
    InMux I__3212 (
            .O(N__14777),
            .I(N__14768));
    Odrv4 I__3211 (
            .O(N__14774),
            .I(L3_tx_data_3));
    Odrv12 I__3210 (
            .O(N__14771),
            .I(L3_tx_data_3));
    LocalMux I__3209 (
            .O(N__14768),
            .I(L3_tx_data_3));
    InMux I__3208 (
            .O(N__14761),
            .I(N__14758));
    LocalMux I__3207 (
            .O(N__14758),
            .I(\Lab_UT.alarmcharZ0Z_0 ));
    SRMux I__3206 (
            .O(N__14755),
            .I(N__14752));
    LocalMux I__3205 (
            .O(N__14752),
            .I(N__14748));
    InMux I__3204 (
            .O(N__14751),
            .I(N__14745));
    Span4Mux_h I__3203 (
            .O(N__14748),
            .I(N__14742));
    LocalMux I__3202 (
            .O(N__14745),
            .I(N__14739));
    Odrv4 I__3201 (
            .O(N__14742),
            .I(\Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1 ));
    Odrv12 I__3200 (
            .O(N__14739),
            .I(\Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1 ));
    InMux I__3199 (
            .O(N__14734),
            .I(N__14728));
    InMux I__3198 (
            .O(N__14733),
            .I(N__14728));
    LocalMux I__3197 (
            .O(N__14728),
            .I(N__14725));
    Span4Mux_h I__3196 (
            .O(N__14725),
            .I(N__14722));
    Span4Mux_h I__3195 (
            .O(N__14722),
            .I(N__14718));
    InMux I__3194 (
            .O(N__14721),
            .I(N__14715));
    Odrv4 I__3193 (
            .O(N__14718),
            .I(L3_tx_data_5));
    LocalMux I__3192 (
            .O(N__14715),
            .I(L3_tx_data_5));
    CascadeMux I__3191 (
            .O(N__14710),
            .I(\Lab_UT.dispString.dOutP_0_iv_3_2_cascade_ ));
    InMux I__3190 (
            .O(N__14707),
            .I(N__14701));
    InMux I__3189 (
            .O(N__14706),
            .I(N__14701));
    LocalMux I__3188 (
            .O(N__14701),
            .I(N__14696));
    InMux I__3187 (
            .O(N__14700),
            .I(N__14691));
    InMux I__3186 (
            .O(N__14699),
            .I(N__14691));
    Odrv12 I__3185 (
            .O(N__14696),
            .I(L3_tx_data_2));
    LocalMux I__3184 (
            .O(N__14691),
            .I(L3_tx_data_2));
    InMux I__3183 (
            .O(N__14686),
            .I(N__14680));
    InMux I__3182 (
            .O(N__14685),
            .I(N__14680));
    LocalMux I__3181 (
            .O(N__14680),
            .I(N__14677));
    Span4Mux_v I__3180 (
            .O(N__14677),
            .I(N__14673));
    CascadeMux I__3179 (
            .O(N__14676),
            .I(N__14670));
    Span4Mux_h I__3178 (
            .O(N__14673),
            .I(N__14667));
    InMux I__3177 (
            .O(N__14670),
            .I(N__14664));
    Odrv4 I__3176 (
            .O(N__14667),
            .I(L3_tx_data_6));
    LocalMux I__3175 (
            .O(N__14664),
            .I(L3_tx_data_6));
    InMux I__3174 (
            .O(N__14659),
            .I(N__14656));
    LocalMux I__3173 (
            .O(N__14656),
            .I(N__14652));
    InMux I__3172 (
            .O(N__14655),
            .I(N__14649));
    Odrv12 I__3171 (
            .O(N__14652),
            .I(L3_tx_data_4));
    LocalMux I__3170 (
            .O(N__14649),
            .I(L3_tx_data_4));
    CascadeMux I__3169 (
            .O(N__14644),
            .I(\Lab_UT.dictrl.un1_state_12_cascade_ ));
    InMux I__3168 (
            .O(N__14641),
            .I(N__14638));
    LocalMux I__3167 (
            .O(N__14638),
            .I(\Lab_UT.didp.m37_nsZ0Z_1 ));
    InMux I__3166 (
            .O(N__14635),
            .I(N__14632));
    LocalMux I__3165 (
            .O(N__14632),
            .I(N__14624));
    InMux I__3164 (
            .O(N__14631),
            .I(N__14619));
    InMux I__3163 (
            .O(N__14630),
            .I(N__14619));
    InMux I__3162 (
            .O(N__14629),
            .I(N__14612));
    InMux I__3161 (
            .O(N__14628),
            .I(N__14612));
    InMux I__3160 (
            .O(N__14627),
            .I(N__14612));
    Odrv4 I__3159 (
            .O(N__14624),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__3158 (
            .O(N__14619),
            .I(\Lab_UT.state_i_3_1 ));
    LocalMux I__3157 (
            .O(N__14612),
            .I(\Lab_UT.state_i_3_1 ));
    CascadeMux I__3156 (
            .O(N__14605),
            .I(N__14598));
    InMux I__3155 (
            .O(N__14604),
            .I(N__14594));
    CascadeMux I__3154 (
            .O(N__14603),
            .I(N__14591));
    CascadeMux I__3153 (
            .O(N__14602),
            .I(N__14588));
    InMux I__3152 (
            .O(N__14601),
            .I(N__14584));
    InMux I__3151 (
            .O(N__14598),
            .I(N__14577));
    InMux I__3150 (
            .O(N__14597),
            .I(N__14577));
    LocalMux I__3149 (
            .O(N__14594),
            .I(N__14574));
    InMux I__3148 (
            .O(N__14591),
            .I(N__14567));
    InMux I__3147 (
            .O(N__14588),
            .I(N__14567));
    InMux I__3146 (
            .O(N__14587),
            .I(N__14567));
    LocalMux I__3145 (
            .O(N__14584),
            .I(N__14564));
    InMux I__3144 (
            .O(N__14583),
            .I(N__14559));
    InMux I__3143 (
            .O(N__14582),
            .I(N__14559));
    LocalMux I__3142 (
            .O(N__14577),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__3141 (
            .O(N__14574),
            .I(\Lab_UT.state_2 ));
    LocalMux I__3140 (
            .O(N__14567),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__3139 (
            .O(N__14564),
            .I(\Lab_UT.state_2 ));
    LocalMux I__3138 (
            .O(N__14559),
            .I(\Lab_UT.state_2 ));
    CascadeMux I__3137 (
            .O(N__14548),
            .I(N__14543));
    InMux I__3136 (
            .O(N__14547),
            .I(N__14538));
    InMux I__3135 (
            .O(N__14546),
            .I(N__14533));
    InMux I__3134 (
            .O(N__14543),
            .I(N__14533));
    CascadeMux I__3133 (
            .O(N__14542),
            .I(N__14530));
    CascadeMux I__3132 (
            .O(N__14541),
            .I(N__14526));
    LocalMux I__3131 (
            .O(N__14538),
            .I(N__14523));
    LocalMux I__3130 (
            .O(N__14533),
            .I(N__14520));
    InMux I__3129 (
            .O(N__14530),
            .I(N__14517));
    InMux I__3128 (
            .O(N__14529),
            .I(N__14514));
    InMux I__3127 (
            .O(N__14526),
            .I(N__14511));
    Odrv12 I__3126 (
            .O(N__14523),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__3125 (
            .O(N__14520),
            .I(\Lab_UT.state_3 ));
    LocalMux I__3124 (
            .O(N__14517),
            .I(\Lab_UT.state_3 ));
    LocalMux I__3123 (
            .O(N__14514),
            .I(\Lab_UT.state_3 ));
    LocalMux I__3122 (
            .O(N__14511),
            .I(\Lab_UT.state_3 ));
    CascadeMux I__3121 (
            .O(N__14500),
            .I(\Lab_UT.dictrl.un1_state_24_ns_1_cascade_ ));
    CascadeMux I__3120 (
            .O(N__14497),
            .I(N__14493));
    InMux I__3119 (
            .O(N__14496),
            .I(N__14489));
    InMux I__3118 (
            .O(N__14493),
            .I(N__14486));
    InMux I__3117 (
            .O(N__14492),
            .I(N__14483));
    LocalMux I__3116 (
            .O(N__14489),
            .I(N__14480));
    LocalMux I__3115 (
            .O(N__14486),
            .I(N__14477));
    LocalMux I__3114 (
            .O(N__14483),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    Odrv4 I__3113 (
            .O(N__14480),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    Odrv4 I__3112 (
            .O(N__14477),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ));
    CascadeMux I__3111 (
            .O(N__14470),
            .I(N__14466));
    InMux I__3110 (
            .O(N__14469),
            .I(N__14462));
    InMux I__3109 (
            .O(N__14466),
            .I(N__14457));
    InMux I__3108 (
            .O(N__14465),
            .I(N__14457));
    LocalMux I__3107 (
            .O(N__14462),
            .I(N__14454));
    LocalMux I__3106 (
            .O(N__14457),
            .I(\Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1 ));
    Odrv4 I__3105 (
            .O(N__14454),
            .I(\Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1 ));
    InMux I__3104 (
            .O(N__14449),
            .I(N__14440));
    InMux I__3103 (
            .O(N__14448),
            .I(N__14440));
    InMux I__3102 (
            .O(N__14447),
            .I(N__14437));
    InMux I__3101 (
            .O(N__14446),
            .I(N__14434));
    InMux I__3100 (
            .O(N__14445),
            .I(N__14431));
    LocalMux I__3099 (
            .O(N__14440),
            .I(\Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ));
    LocalMux I__3098 (
            .O(N__14437),
            .I(\Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ));
    LocalMux I__3097 (
            .O(N__14434),
            .I(\Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ));
    LocalMux I__3096 (
            .O(N__14431),
            .I(\Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ));
    CascadeMux I__3095 (
            .O(N__14422),
            .I(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_ ));
    InMux I__3094 (
            .O(N__14419),
            .I(N__14413));
    InMux I__3093 (
            .O(N__14418),
            .I(N__14408));
    InMux I__3092 (
            .O(N__14417),
            .I(N__14408));
    InMux I__3091 (
            .O(N__14416),
            .I(N__14405));
    LocalMux I__3090 (
            .O(N__14413),
            .I(N__14398));
    LocalMux I__3089 (
            .O(N__14408),
            .I(N__14398));
    LocalMux I__3088 (
            .O(N__14405),
            .I(N__14398));
    Odrv4 I__3087 (
            .O(N__14398),
            .I(\Lab_UT.dictrl.next_state_set_0 ));
    InMux I__3086 (
            .O(N__14395),
            .I(N__14392));
    LocalMux I__3085 (
            .O(N__14392),
            .I(\Lab_UT.dictrl.next_state_out_1 ));
    CEMux I__3084 (
            .O(N__14389),
            .I(N__14384));
    CEMux I__3083 (
            .O(N__14388),
            .I(N__14380));
    CEMux I__3082 (
            .O(N__14387),
            .I(N__14377));
    LocalMux I__3081 (
            .O(N__14384),
            .I(N__14374));
    CEMux I__3080 (
            .O(N__14383),
            .I(N__14371));
    LocalMux I__3079 (
            .O(N__14380),
            .I(N__14368));
    LocalMux I__3078 (
            .O(N__14377),
            .I(N__14365));
    Span4Mux_v I__3077 (
            .O(N__14374),
            .I(N__14362));
    LocalMux I__3076 (
            .O(N__14371),
            .I(N__14359));
    Odrv4 I__3075 (
            .O(N__14368),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    Odrv4 I__3074 (
            .O(N__14365),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    Odrv4 I__3073 (
            .O(N__14362),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    Odrv4 I__3072 (
            .O(N__14359),
            .I(\Lab_UT.dictrl.un1_state_21_reti_i ));
    InMux I__3071 (
            .O(N__14350),
            .I(N__14347));
    LocalMux I__3070 (
            .O(N__14347),
            .I(\Lab_UT.didp.countrce4.N_88_i ));
    InMux I__3069 (
            .O(N__14344),
            .I(N__14340));
    InMux I__3068 (
            .O(N__14343),
            .I(N__14337));
    LocalMux I__3067 (
            .O(N__14340),
            .I(N__14334));
    LocalMux I__3066 (
            .O(N__14337),
            .I(N__14331));
    Span4Mux_h I__3065 (
            .O(N__14334),
            .I(N__14328));
    Odrv4 I__3064 (
            .O(N__14331),
            .I(\Lab_UT.N_68_0 ));
    Odrv4 I__3063 (
            .O(N__14328),
            .I(\Lab_UT.N_68_0 ));
    InMux I__3062 (
            .O(N__14323),
            .I(N__14320));
    LocalMux I__3061 (
            .O(N__14320),
            .I(N__14317));
    Span4Mux_v I__3060 (
            .O(N__14317),
            .I(N__14314));
    Odrv4 I__3059 (
            .O(N__14314),
            .I(\Lab_UT.didp.un31_reset_i_a4_1 ));
    InMux I__3058 (
            .O(N__14311),
            .I(N__14305));
    InMux I__3057 (
            .O(N__14310),
            .I(N__14300));
    InMux I__3056 (
            .O(N__14309),
            .I(N__14300));
    InMux I__3055 (
            .O(N__14308),
            .I(N__14297));
    LocalMux I__3054 (
            .O(N__14305),
            .I(N__14294));
    LocalMux I__3053 (
            .O(N__14300),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    LocalMux I__3052 (
            .O(N__14297),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    Odrv4 I__3051 (
            .O(N__14294),
            .I(\Lab_UT.dictrl.next_state_set_1 ));
    CascadeMux I__3050 (
            .O(N__14287),
            .I(N__14283));
    InMux I__3049 (
            .O(N__14286),
            .I(N__14276));
    InMux I__3048 (
            .O(N__14283),
            .I(N__14276));
    InMux I__3047 (
            .O(N__14282),
            .I(N__14273));
    InMux I__3046 (
            .O(N__14281),
            .I(N__14270));
    LocalMux I__3045 (
            .O(N__14276),
            .I(\Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2 ));
    LocalMux I__3044 (
            .O(N__14273),
            .I(\Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2 ));
    LocalMux I__3043 (
            .O(N__14270),
            .I(\Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2 ));
    InMux I__3042 (
            .O(N__14263),
            .I(N__14255));
    InMux I__3041 (
            .O(N__14262),
            .I(N__14255));
    InMux I__3040 (
            .O(N__14261),
            .I(N__14252));
    InMux I__3039 (
            .O(N__14260),
            .I(N__14249));
    LocalMux I__3038 (
            .O(N__14255),
            .I(\Lab_UT.m37_ns ));
    LocalMux I__3037 (
            .O(N__14252),
            .I(\Lab_UT.m37_ns ));
    LocalMux I__3036 (
            .O(N__14249),
            .I(\Lab_UT.m37_ns ));
    InMux I__3035 (
            .O(N__14242),
            .I(N__14218));
    InMux I__3034 (
            .O(N__14241),
            .I(N__14218));
    InMux I__3033 (
            .O(N__14240),
            .I(N__14212));
    InMux I__3032 (
            .O(N__14239),
            .I(N__14204));
    InMux I__3031 (
            .O(N__14238),
            .I(N__14199));
    InMux I__3030 (
            .O(N__14237),
            .I(N__14199));
    InMux I__3029 (
            .O(N__14236),
            .I(N__14192));
    InMux I__3028 (
            .O(N__14235),
            .I(N__14192));
    InMux I__3027 (
            .O(N__14234),
            .I(N__14192));
    InMux I__3026 (
            .O(N__14233),
            .I(N__14187));
    InMux I__3025 (
            .O(N__14232),
            .I(N__14187));
    InMux I__3024 (
            .O(N__14231),
            .I(N__14180));
    InMux I__3023 (
            .O(N__14230),
            .I(N__14180));
    InMux I__3022 (
            .O(N__14229),
            .I(N__14180));
    InMux I__3021 (
            .O(N__14228),
            .I(N__14173));
    InMux I__3020 (
            .O(N__14227),
            .I(N__14173));
    InMux I__3019 (
            .O(N__14226),
            .I(N__14173));
    InMux I__3018 (
            .O(N__14225),
            .I(N__14166));
    InMux I__3017 (
            .O(N__14224),
            .I(N__14166));
    InMux I__3016 (
            .O(N__14223),
            .I(N__14166));
    LocalMux I__3015 (
            .O(N__14218),
            .I(N__14163));
    InMux I__3014 (
            .O(N__14217),
            .I(N__14156));
    InMux I__3013 (
            .O(N__14216),
            .I(N__14156));
    InMux I__3012 (
            .O(N__14215),
            .I(N__14156));
    LocalMux I__3011 (
            .O(N__14212),
            .I(N__14153));
    InMux I__3010 (
            .O(N__14211),
            .I(N__14146));
    InMux I__3009 (
            .O(N__14210),
            .I(N__14146));
    InMux I__3008 (
            .O(N__14209),
            .I(N__14146));
    InMux I__3007 (
            .O(N__14208),
            .I(N__14141));
    InMux I__3006 (
            .O(N__14207),
            .I(N__14141));
    LocalMux I__3005 (
            .O(N__14204),
            .I(N__14138));
    LocalMux I__3004 (
            .O(N__14199),
            .I(N__14129));
    LocalMux I__3003 (
            .O(N__14192),
            .I(N__14129));
    LocalMux I__3002 (
            .O(N__14187),
            .I(N__14129));
    LocalMux I__3001 (
            .O(N__14180),
            .I(N__14129));
    LocalMux I__3000 (
            .O(N__14173),
            .I(N__14126));
    LocalMux I__2999 (
            .O(N__14166),
            .I(N__14115));
    Span4Mux_h I__2998 (
            .O(N__14163),
            .I(N__14115));
    LocalMux I__2997 (
            .O(N__14156),
            .I(N__14115));
    Span4Mux_v I__2996 (
            .O(N__14153),
            .I(N__14115));
    LocalMux I__2995 (
            .O(N__14146),
            .I(N__14104));
    LocalMux I__2994 (
            .O(N__14141),
            .I(N__14104));
    Span4Mux_v I__2993 (
            .O(N__14138),
            .I(N__14104));
    Span4Mux_v I__2992 (
            .O(N__14129),
            .I(N__14104));
    Span4Mux_v I__2991 (
            .O(N__14126),
            .I(N__14104));
    InMux I__2990 (
            .O(N__14125),
            .I(N__14099));
    InMux I__2989 (
            .O(N__14124),
            .I(N__14099));
    Span4Mux_v I__2988 (
            .O(N__14115),
            .I(N__14096));
    Span4Mux_h I__2987 (
            .O(N__14104),
            .I(N__14093));
    LocalMux I__2986 (
            .O(N__14099),
            .I(\Lab_UT.Run ));
    Odrv4 I__2985 (
            .O(N__14096),
            .I(\Lab_UT.Run ));
    Odrv4 I__2984 (
            .O(N__14093),
            .I(\Lab_UT.Run ));
    InMux I__2983 (
            .O(N__14086),
            .I(N__14082));
    InMux I__2982 (
            .O(N__14085),
            .I(N__14079));
    LocalMux I__2981 (
            .O(N__14082),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    LocalMux I__2980 (
            .O(N__14079),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    InMux I__2979 (
            .O(N__14074),
            .I(N__14069));
    InMux I__2978 (
            .O(N__14073),
            .I(N__14064));
    InMux I__2977 (
            .O(N__14072),
            .I(N__14064));
    LocalMux I__2976 (
            .O(N__14069),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    LocalMux I__2975 (
            .O(N__14064),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    CascadeMux I__2974 (
            .O(N__14059),
            .I(\Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_ ));
    InMux I__2973 (
            .O(N__14056),
            .I(N__14053));
    LocalMux I__2972 (
            .O(N__14053),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa ));
    InMux I__2971 (
            .O(N__14050),
            .I(N__14047));
    LocalMux I__2970 (
            .O(N__14047),
            .I(N__14044));
    Odrv4 I__2969 (
            .O(N__14044),
            .I(\Lab_UT.didp.m34_nsZ0Z_1 ));
    InMux I__2968 (
            .O(N__14041),
            .I(N__14035));
    InMux I__2967 (
            .O(N__14040),
            .I(N__14035));
    LocalMux I__2966 (
            .O(N__14035),
            .I(N__14031));
    InMux I__2965 (
            .O(N__14034),
            .I(N__14028));
    Span4Mux_h I__2964 (
            .O(N__14031),
            .I(N__14025));
    LocalMux I__2963 (
            .O(N__14028),
            .I(\Lab_UT.dictrl.next_state16Z0Z_4 ));
    Odrv4 I__2962 (
            .O(N__14025),
            .I(\Lab_UT.dictrl.next_state16Z0Z_4 ));
    CascadeMux I__2961 (
            .O(N__14020),
            .I(\Lab_UT.m34_ns_cascade_ ));
    InMux I__2960 (
            .O(N__14017),
            .I(N__14014));
    LocalMux I__2959 (
            .O(N__14014),
            .I(N__14011));
    Span4Mux_s2_h I__2958 (
            .O(N__14011),
            .I(N__14008));
    Span4Mux_h I__2957 (
            .O(N__14008),
            .I(N__14003));
    InMux I__2956 (
            .O(N__14007),
            .I(N__14000));
    InMux I__2955 (
            .O(N__14006),
            .I(N__13997));
    Odrv4 I__2954 (
            .O(N__14003),
            .I(resetGen_escKey_4));
    LocalMux I__2953 (
            .O(N__14000),
            .I(resetGen_escKey_4));
    LocalMux I__2952 (
            .O(N__13997),
            .I(resetGen_escKey_4));
    InMux I__2951 (
            .O(N__13990),
            .I(N__13987));
    LocalMux I__2950 (
            .O(N__13987),
            .I(N__13984));
    Span4Mux_h I__2949 (
            .O(N__13984),
            .I(N__13975));
    InMux I__2948 (
            .O(N__13983),
            .I(N__13970));
    InMux I__2947 (
            .O(N__13982),
            .I(N__13970));
    InMux I__2946 (
            .O(N__13981),
            .I(N__13961));
    InMux I__2945 (
            .O(N__13980),
            .I(N__13961));
    InMux I__2944 (
            .O(N__13979),
            .I(N__13961));
    InMux I__2943 (
            .O(N__13978),
            .I(N__13961));
    Odrv4 I__2942 (
            .O(N__13975),
            .I(bu_rx_data_1));
    LocalMux I__2941 (
            .O(N__13970),
            .I(bu_rx_data_1));
    LocalMux I__2940 (
            .O(N__13961),
            .I(bu_rx_data_1));
    CascadeMux I__2939 (
            .O(N__13954),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__2938 (
            .O(N__13951),
            .I(N__13948));
    LocalMux I__2937 (
            .O(N__13948),
            .I(N__13943));
    CascadeMux I__2936 (
            .O(N__13947),
            .I(N__13940));
    CascadeMux I__2935 (
            .O(N__13946),
            .I(N__13934));
    Span4Mux_h I__2934 (
            .O(N__13943),
            .I(N__13931));
    InMux I__2933 (
            .O(N__13940),
            .I(N__13920));
    InMux I__2932 (
            .O(N__13939),
            .I(N__13920));
    InMux I__2931 (
            .O(N__13938),
            .I(N__13920));
    InMux I__2930 (
            .O(N__13937),
            .I(N__13920));
    InMux I__2929 (
            .O(N__13934),
            .I(N__13920));
    Span4Mux_h I__2928 (
            .O(N__13931),
            .I(N__13917));
    LocalMux I__2927 (
            .O(N__13920),
            .I(\resetGen.reset_countZ0Z_4 ));
    Odrv4 I__2926 (
            .O(N__13917),
            .I(\resetGen.reset_countZ0Z_4 ));
    InMux I__2925 (
            .O(N__13912),
            .I(N__13909));
    LocalMux I__2924 (
            .O(N__13909),
            .I(\Lab_UT.dictrl.next_state_out_3 ));
    SRMux I__2923 (
            .O(N__13906),
            .I(N__13903));
    LocalMux I__2922 (
            .O(N__13903),
            .I(N__13900));
    Odrv12 I__2921 (
            .O(N__13900),
            .I(\Lab_UT.m34_ns ));
    CascadeMux I__2920 (
            .O(N__13897),
            .I(\Lab_UT.didp.N_164_cascade_ ));
    SRMux I__2919 (
            .O(N__13894),
            .I(N__13891));
    LocalMux I__2918 (
            .O(N__13891),
            .I(N__13888));
    Span4Mux_v I__2917 (
            .O(N__13888),
            .I(N__13885));
    Span4Mux_h I__2916 (
            .O(N__13885),
            .I(N__13881));
    InMux I__2915 (
            .O(N__13884),
            .I(N__13878));
    Odrv4 I__2914 (
            .O(N__13881),
            .I(\Lab_UT.m42 ));
    LocalMux I__2913 (
            .O(N__13878),
            .I(\Lab_UT.m42 ));
    InMux I__2912 (
            .O(N__13873),
            .I(N__13870));
    LocalMux I__2911 (
            .O(N__13870),
            .I(\Lab_UT.bcd2segment2.segment_i_0Z0Z_1 ));
    CascadeMux I__2910 (
            .O(N__13867),
            .I(\Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_ ));
    InMux I__2909 (
            .O(N__13864),
            .I(N__13861));
    LocalMux I__2908 (
            .O(N__13861),
            .I(N__13858));
    Odrv4 I__2907 (
            .O(N__13858),
            .I(\uu2.bitmapZ0Z_87 ));
    CascadeMux I__2906 (
            .O(N__13855),
            .I(\Lab_UT.three_2_cascade_ ));
    InMux I__2905 (
            .O(N__13852),
            .I(N__13849));
    LocalMux I__2904 (
            .O(N__13849),
            .I(\Lab_UT.didp.countrce1.un20_qPone ));
    InMux I__2903 (
            .O(N__13846),
            .I(N__13843));
    LocalMux I__2902 (
            .O(N__13843),
            .I(\uu2.mem0.g0_7_4_0 ));
    CascadeMux I__2901 (
            .O(N__13840),
            .I(N__13835));
    CascadeMux I__2900 (
            .O(N__13839),
            .I(N__13832));
    InMux I__2899 (
            .O(N__13838),
            .I(N__13825));
    InMux I__2898 (
            .O(N__13835),
            .I(N__13817));
    InMux I__2897 (
            .O(N__13832),
            .I(N__13817));
    InMux I__2896 (
            .O(N__13831),
            .I(N__13817));
    InMux I__2895 (
            .O(N__13830),
            .I(N__13814));
    InMux I__2894 (
            .O(N__13829),
            .I(N__13811));
    InMux I__2893 (
            .O(N__13828),
            .I(N__13808));
    LocalMux I__2892 (
            .O(N__13825),
            .I(N__13805));
    InMux I__2891 (
            .O(N__13824),
            .I(N__13797));
    LocalMux I__2890 (
            .O(N__13817),
            .I(N__13792));
    LocalMux I__2889 (
            .O(N__13814),
            .I(N__13792));
    LocalMux I__2888 (
            .O(N__13811),
            .I(N__13789));
    LocalMux I__2887 (
            .O(N__13808),
            .I(N__13786));
    Span4Mux_h I__2886 (
            .O(N__13805),
            .I(N__13783));
    InMux I__2885 (
            .O(N__13804),
            .I(N__13780));
    InMux I__2884 (
            .O(N__13803),
            .I(N__13771));
    InMux I__2883 (
            .O(N__13802),
            .I(N__13771));
    InMux I__2882 (
            .O(N__13801),
            .I(N__13771));
    InMux I__2881 (
            .O(N__13800),
            .I(N__13771));
    LocalMux I__2880 (
            .O(N__13797),
            .I(N__13764));
    Span4Mux_v I__2879 (
            .O(N__13792),
            .I(N__13764));
    Span4Mux_h I__2878 (
            .O(N__13789),
            .I(N__13764));
    Odrv4 I__2877 (
            .O(N__13786),
            .I(\uu2.N_46 ));
    Odrv4 I__2876 (
            .O(N__13783),
            .I(\uu2.N_46 ));
    LocalMux I__2875 (
            .O(N__13780),
            .I(\uu2.N_46 ));
    LocalMux I__2874 (
            .O(N__13771),
            .I(\uu2.N_46 ));
    Odrv4 I__2873 (
            .O(N__13764),
            .I(\uu2.N_46 ));
    CascadeMux I__2872 (
            .O(N__13753),
            .I(N__13748));
    CascadeMux I__2871 (
            .O(N__13752),
            .I(N__13743));
    CascadeMux I__2870 (
            .O(N__13751),
            .I(N__13740));
    InMux I__2869 (
            .O(N__13748),
            .I(N__13734));
    InMux I__2868 (
            .O(N__13747),
            .I(N__13731));
    InMux I__2867 (
            .O(N__13746),
            .I(N__13728));
    InMux I__2866 (
            .O(N__13743),
            .I(N__13723));
    InMux I__2865 (
            .O(N__13740),
            .I(N__13723));
    InMux I__2864 (
            .O(N__13739),
            .I(N__13720));
    InMux I__2863 (
            .O(N__13738),
            .I(N__13717));
    InMux I__2862 (
            .O(N__13737),
            .I(N__13713));
    LocalMux I__2861 (
            .O(N__13734),
            .I(N__13703));
    LocalMux I__2860 (
            .O(N__13731),
            .I(N__13700));
    LocalMux I__2859 (
            .O(N__13728),
            .I(N__13693));
    LocalMux I__2858 (
            .O(N__13723),
            .I(N__13693));
    LocalMux I__2857 (
            .O(N__13720),
            .I(N__13693));
    LocalMux I__2856 (
            .O(N__13717),
            .I(N__13690));
    InMux I__2855 (
            .O(N__13716),
            .I(N__13687));
    LocalMux I__2854 (
            .O(N__13713),
            .I(N__13684));
    InMux I__2853 (
            .O(N__13712),
            .I(N__13671));
    InMux I__2852 (
            .O(N__13711),
            .I(N__13671));
    InMux I__2851 (
            .O(N__13710),
            .I(N__13671));
    InMux I__2850 (
            .O(N__13709),
            .I(N__13671));
    InMux I__2849 (
            .O(N__13708),
            .I(N__13664));
    InMux I__2848 (
            .O(N__13707),
            .I(N__13664));
    InMux I__2847 (
            .O(N__13706),
            .I(N__13664));
    Span4Mux_v I__2846 (
            .O(N__13703),
            .I(N__13655));
    Span4Mux_v I__2845 (
            .O(N__13700),
            .I(N__13655));
    Span4Mux_v I__2844 (
            .O(N__13693),
            .I(N__13655));
    Span4Mux_v I__2843 (
            .O(N__13690),
            .I(N__13655));
    LocalMux I__2842 (
            .O(N__13687),
            .I(N__13650));
    Span4Mux_h I__2841 (
            .O(N__13684),
            .I(N__13650));
    InMux I__2840 (
            .O(N__13683),
            .I(N__13641));
    InMux I__2839 (
            .O(N__13682),
            .I(N__13641));
    InMux I__2838 (
            .O(N__13681),
            .I(N__13641));
    InMux I__2837 (
            .O(N__13680),
            .I(N__13641));
    LocalMux I__2836 (
            .O(N__13671),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2835 (
            .O(N__13664),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2834 (
            .O(N__13655),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2833 (
            .O(N__13650),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2832 (
            .O(N__13641),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__2831 (
            .O(N__13630),
            .I(N__13620));
    InMux I__2830 (
            .O(N__13629),
            .I(N__13616));
    InMux I__2829 (
            .O(N__13628),
            .I(N__13613));
    CascadeMux I__2828 (
            .O(N__13627),
            .I(N__13610));
    CascadeMux I__2827 (
            .O(N__13626),
            .I(N__13606));
    InMux I__2826 (
            .O(N__13625),
            .I(N__13595));
    InMux I__2825 (
            .O(N__13624),
            .I(N__13595));
    InMux I__2824 (
            .O(N__13623),
            .I(N__13595));
    InMux I__2823 (
            .O(N__13620),
            .I(N__13595));
    InMux I__2822 (
            .O(N__13619),
            .I(N__13595));
    LocalMux I__2821 (
            .O(N__13616),
            .I(N__13588));
    LocalMux I__2820 (
            .O(N__13613),
            .I(N__13588));
    InMux I__2819 (
            .O(N__13610),
            .I(N__13585));
    InMux I__2818 (
            .O(N__13609),
            .I(N__13580));
    InMux I__2817 (
            .O(N__13606),
            .I(N__13580));
    LocalMux I__2816 (
            .O(N__13595),
            .I(N__13574));
    InMux I__2815 (
            .O(N__13594),
            .I(N__13569));
    InMux I__2814 (
            .O(N__13593),
            .I(N__13569));
    Span4Mux_v I__2813 (
            .O(N__13588),
            .I(N__13564));
    LocalMux I__2812 (
            .O(N__13585),
            .I(N__13564));
    LocalMux I__2811 (
            .O(N__13580),
            .I(N__13561));
    InMux I__2810 (
            .O(N__13579),
            .I(N__13554));
    InMux I__2809 (
            .O(N__13578),
            .I(N__13554));
    InMux I__2808 (
            .O(N__13577),
            .I(N__13554));
    Span4Mux_v I__2807 (
            .O(N__13574),
            .I(N__13551));
    LocalMux I__2806 (
            .O(N__13569),
            .I(N__13546));
    Span4Mux_h I__2805 (
            .O(N__13564),
            .I(N__13546));
    Span4Mux_h I__2804 (
            .O(N__13561),
            .I(N__13541));
    LocalMux I__2803 (
            .O(N__13554),
            .I(N__13541));
    Odrv4 I__2802 (
            .O(N__13551),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2801 (
            .O(N__13546),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2800 (
            .O(N__13541),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    CEMux I__2799 (
            .O(N__13534),
            .I(N__13530));
    CEMux I__2798 (
            .O(N__13533),
            .I(N__13527));
    LocalMux I__2797 (
            .O(N__13530),
            .I(N__13524));
    LocalMux I__2796 (
            .O(N__13527),
            .I(N__13520));
    Span4Mux_v I__2795 (
            .O(N__13524),
            .I(N__13517));
    CEMux I__2794 (
            .O(N__13523),
            .I(N__13514));
    Odrv4 I__2793 (
            .O(N__13520),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    Odrv4 I__2792 (
            .O(N__13517),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    LocalMux I__2791 (
            .O(N__13514),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    InMux I__2790 (
            .O(N__13507),
            .I(N__13495));
    CascadeMux I__2789 (
            .O(N__13506),
            .I(N__13491));
    CascadeMux I__2788 (
            .O(N__13505),
            .I(N__13488));
    CascadeMux I__2787 (
            .O(N__13504),
            .I(N__13485));
    CascadeMux I__2786 (
            .O(N__13503),
            .I(N__13482));
    InMux I__2785 (
            .O(N__13502),
            .I(N__13479));
    InMux I__2784 (
            .O(N__13501),
            .I(N__13476));
    InMux I__2783 (
            .O(N__13500),
            .I(N__13471));
    InMux I__2782 (
            .O(N__13499),
            .I(N__13471));
    CascadeMux I__2781 (
            .O(N__13498),
            .I(N__13468));
    LocalMux I__2780 (
            .O(N__13495),
            .I(N__13465));
    InMux I__2779 (
            .O(N__13494),
            .I(N__13459));
    InMux I__2778 (
            .O(N__13491),
            .I(N__13459));
    InMux I__2777 (
            .O(N__13488),
            .I(N__13452));
    InMux I__2776 (
            .O(N__13485),
            .I(N__13452));
    InMux I__2775 (
            .O(N__13482),
            .I(N__13452));
    LocalMux I__2774 (
            .O(N__13479),
            .I(N__13449));
    LocalMux I__2773 (
            .O(N__13476),
            .I(N__13446));
    LocalMux I__2772 (
            .O(N__13471),
            .I(N__13443));
    InMux I__2771 (
            .O(N__13468),
            .I(N__13440));
    Span4Mux_v I__2770 (
            .O(N__13465),
            .I(N__13437));
    InMux I__2769 (
            .O(N__13464),
            .I(N__13434));
    LocalMux I__2768 (
            .O(N__13459),
            .I(N__13429));
    LocalMux I__2767 (
            .O(N__13452),
            .I(N__13429));
    Span4Mux_h I__2766 (
            .O(N__13449),
            .I(N__13422));
    Span4Mux_h I__2765 (
            .O(N__13446),
            .I(N__13422));
    Span4Mux_h I__2764 (
            .O(N__13443),
            .I(N__13422));
    LocalMux I__2763 (
            .O(N__13440),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2762 (
            .O(N__13437),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2761 (
            .O(N__13434),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2760 (
            .O(N__13429),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2759 (
            .O(N__13422),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__2758 (
            .O(N__13411),
            .I(N__13406));
    InMux I__2757 (
            .O(N__13410),
            .I(N__13403));
    CascadeMux I__2756 (
            .O(N__13409),
            .I(N__13399));
    LocalMux I__2755 (
            .O(N__13406),
            .I(N__13391));
    LocalMux I__2754 (
            .O(N__13403),
            .I(N__13388));
    CascadeMux I__2753 (
            .O(N__13402),
            .I(N__13385));
    InMux I__2752 (
            .O(N__13399),
            .I(N__13377));
    InMux I__2751 (
            .O(N__13398),
            .I(N__13377));
    InMux I__2750 (
            .O(N__13397),
            .I(N__13377));
    CascadeMux I__2749 (
            .O(N__13396),
            .I(N__13370));
    CascadeMux I__2748 (
            .O(N__13395),
            .I(N__13367));
    InMux I__2747 (
            .O(N__13394),
            .I(N__13364));
    Span4Mux_h I__2746 (
            .O(N__13391),
            .I(N__13361));
    Span4Mux_h I__2745 (
            .O(N__13388),
            .I(N__13358));
    InMux I__2744 (
            .O(N__13385),
            .I(N__13353));
    InMux I__2743 (
            .O(N__13384),
            .I(N__13353));
    LocalMux I__2742 (
            .O(N__13377),
            .I(N__13350));
    InMux I__2741 (
            .O(N__13376),
            .I(N__13343));
    InMux I__2740 (
            .O(N__13375),
            .I(N__13343));
    InMux I__2739 (
            .O(N__13374),
            .I(N__13343));
    InMux I__2738 (
            .O(N__13373),
            .I(N__13340));
    InMux I__2737 (
            .O(N__13370),
            .I(N__13335));
    InMux I__2736 (
            .O(N__13367),
            .I(N__13335));
    LocalMux I__2735 (
            .O(N__13364),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2734 (
            .O(N__13361),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2733 (
            .O(N__13358),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2732 (
            .O(N__13353),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2731 (
            .O(N__13350),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2730 (
            .O(N__13343),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2729 (
            .O(N__13340),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2728 (
            .O(N__13335),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__2727 (
            .O(N__13318),
            .I(N__13313));
    InMux I__2726 (
            .O(N__13317),
            .I(N__13310));
    InMux I__2725 (
            .O(N__13316),
            .I(N__13307));
    LocalMux I__2724 (
            .O(N__13313),
            .I(N__13300));
    LocalMux I__2723 (
            .O(N__13310),
            .I(N__13297));
    LocalMux I__2722 (
            .O(N__13307),
            .I(N__13294));
    InMux I__2721 (
            .O(N__13306),
            .I(N__13291));
    CascadeMux I__2720 (
            .O(N__13305),
            .I(N__13284));
    CascadeMux I__2719 (
            .O(N__13304),
            .I(N__13281));
    InMux I__2718 (
            .O(N__13303),
            .I(N__13277));
    Span4Mux_h I__2717 (
            .O(N__13300),
            .I(N__13274));
    Span4Mux_h I__2716 (
            .O(N__13297),
            .I(N__13271));
    Span4Mux_h I__2715 (
            .O(N__13294),
            .I(N__13268));
    LocalMux I__2714 (
            .O(N__13291),
            .I(N__13265));
    InMux I__2713 (
            .O(N__13290),
            .I(N__13260));
    InMux I__2712 (
            .O(N__13289),
            .I(N__13260));
    InMux I__2711 (
            .O(N__13288),
            .I(N__13253));
    InMux I__2710 (
            .O(N__13287),
            .I(N__13253));
    InMux I__2709 (
            .O(N__13284),
            .I(N__13253));
    InMux I__2708 (
            .O(N__13281),
            .I(N__13248));
    InMux I__2707 (
            .O(N__13280),
            .I(N__13248));
    LocalMux I__2706 (
            .O(N__13277),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2705 (
            .O(N__13274),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2704 (
            .O(N__13271),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2703 (
            .O(N__13268),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2702 (
            .O(N__13265),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2701 (
            .O(N__13260),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2700 (
            .O(N__13253),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2699 (
            .O(N__13248),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    InMux I__2698 (
            .O(N__13231),
            .I(N__13226));
    InMux I__2697 (
            .O(N__13230),
            .I(N__13220));
    InMux I__2696 (
            .O(N__13229),
            .I(N__13220));
    LocalMux I__2695 (
            .O(N__13226),
            .I(N__13217));
    InMux I__2694 (
            .O(N__13225),
            .I(N__13209));
    LocalMux I__2693 (
            .O(N__13220),
            .I(N__13206));
    Span4Mux_h I__2692 (
            .O(N__13217),
            .I(N__13197));
    InMux I__2691 (
            .O(N__13216),
            .I(N__13194));
    InMux I__2690 (
            .O(N__13215),
            .I(N__13191));
    InMux I__2689 (
            .O(N__13214),
            .I(N__13186));
    InMux I__2688 (
            .O(N__13213),
            .I(N__13186));
    InMux I__2687 (
            .O(N__13212),
            .I(N__13183));
    LocalMux I__2686 (
            .O(N__13209),
            .I(N__13180));
    Span4Mux_h I__2685 (
            .O(N__13206),
            .I(N__13177));
    InMux I__2684 (
            .O(N__13205),
            .I(N__13168));
    InMux I__2683 (
            .O(N__13204),
            .I(N__13168));
    InMux I__2682 (
            .O(N__13203),
            .I(N__13168));
    InMux I__2681 (
            .O(N__13202),
            .I(N__13168));
    InMux I__2680 (
            .O(N__13201),
            .I(N__13163));
    InMux I__2679 (
            .O(N__13200),
            .I(N__13163));
    Span4Mux_v I__2678 (
            .O(N__13197),
            .I(N__13154));
    LocalMux I__2677 (
            .O(N__13194),
            .I(N__13154));
    LocalMux I__2676 (
            .O(N__13191),
            .I(N__13154));
    LocalMux I__2675 (
            .O(N__13186),
            .I(N__13154));
    LocalMux I__2674 (
            .O(N__13183),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2673 (
            .O(N__13180),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2672 (
            .O(N__13177),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2671 (
            .O(N__13168),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2670 (
            .O(N__13163),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2669 (
            .O(N__13154),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__2668 (
            .O(N__13141),
            .I(N__13138));
    LocalMux I__2667 (
            .O(N__13138),
            .I(N__13135));
    Odrv12 I__2666 (
            .O(N__13135),
            .I(\uu2.mem0.g0_16_1 ));
    CascadeMux I__2665 (
            .O(N__13132),
            .I(\Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_ ));
    CascadeMux I__2664 (
            .O(N__13129),
            .I(N__13126));
    InMux I__2663 (
            .O(N__13126),
            .I(N__13123));
    LocalMux I__2662 (
            .O(N__13123),
            .I(N__13120));
    Span4Mux_v I__2661 (
            .O(N__13120),
            .I(N__13117));
    Odrv4 I__2660 (
            .O(N__13117),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__2659 (
            .O(N__13114),
            .I(\Lab_UT.nine_cascade_ ));
    CascadeMux I__2658 (
            .O(N__13111),
            .I(N__13106));
    InMux I__2657 (
            .O(N__13110),
            .I(N__13099));
    InMux I__2656 (
            .O(N__13109),
            .I(N__13099));
    InMux I__2655 (
            .O(N__13106),
            .I(N__13099));
    LocalMux I__2654 (
            .O(N__13099),
            .I(N__13096));
    Span4Mux_h I__2653 (
            .O(N__13096),
            .I(N__13093));
    Odrv4 I__2652 (
            .O(N__13093),
            .I(\uu2.N_49 ));
    CascadeMux I__2651 (
            .O(N__13090),
            .I(\uu2.mem0.g0_7_5_0_cascade_ ));
    CascadeMux I__2650 (
            .O(N__13087),
            .I(\uu2.mem0.un31_w_data_displaying_1_0_0_cascade_ ));
    InMux I__2649 (
            .O(N__13084),
            .I(N__13081));
    LocalMux I__2648 (
            .O(N__13081),
            .I(N__13078));
    Span4Mux_v I__2647 (
            .O(N__13078),
            .I(N__13075));
    Odrv4 I__2646 (
            .O(N__13075),
            .I(\uu2.mem0.g1_0_1 ));
    CascadeMux I__2645 (
            .O(N__13072),
            .I(N__13066));
    InMux I__2644 (
            .O(N__13071),
            .I(N__13059));
    InMux I__2643 (
            .O(N__13070),
            .I(N__13056));
    InMux I__2642 (
            .O(N__13069),
            .I(N__13053));
    InMux I__2641 (
            .O(N__13066),
            .I(N__13043));
    InMux I__2640 (
            .O(N__13065),
            .I(N__13043));
    InMux I__2639 (
            .O(N__13064),
            .I(N__13043));
    InMux I__2638 (
            .O(N__13063),
            .I(N__13038));
    InMux I__2637 (
            .O(N__13062),
            .I(N__13038));
    LocalMux I__2636 (
            .O(N__13059),
            .I(N__13033));
    LocalMux I__2635 (
            .O(N__13056),
            .I(N__13033));
    LocalMux I__2634 (
            .O(N__13053),
            .I(N__13024));
    InMux I__2633 (
            .O(N__13052),
            .I(N__13021));
    InMux I__2632 (
            .O(N__13051),
            .I(N__13018));
    InMux I__2631 (
            .O(N__13050),
            .I(N__13015));
    LocalMux I__2630 (
            .O(N__13043),
            .I(N__13008));
    LocalMux I__2629 (
            .O(N__13038),
            .I(N__13008));
    Span4Mux_v I__2628 (
            .O(N__13033),
            .I(N__13008));
    InMux I__2627 (
            .O(N__13032),
            .I(N__13003));
    InMux I__2626 (
            .O(N__13031),
            .I(N__13003));
    InMux I__2625 (
            .O(N__13030),
            .I(N__12994));
    InMux I__2624 (
            .O(N__13029),
            .I(N__12994));
    InMux I__2623 (
            .O(N__13028),
            .I(N__12994));
    InMux I__2622 (
            .O(N__13027),
            .I(N__12994));
    Odrv4 I__2621 (
            .O(N__13024),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2620 (
            .O(N__13021),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2619 (
            .O(N__13018),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2618 (
            .O(N__13015),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__2617 (
            .O(N__13008),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2616 (
            .O(N__13003),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__2615 (
            .O(N__12994),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__2614 (
            .O(N__12979),
            .I(N__12975));
    InMux I__2613 (
            .O(N__12978),
            .I(N__12966));
    InMux I__2612 (
            .O(N__12975),
            .I(N__12959));
    InMux I__2611 (
            .O(N__12974),
            .I(N__12959));
    InMux I__2610 (
            .O(N__12973),
            .I(N__12959));
    CascadeMux I__2609 (
            .O(N__12972),
            .I(N__12956));
    InMux I__2608 (
            .O(N__12971),
            .I(N__12949));
    InMux I__2607 (
            .O(N__12970),
            .I(N__12949));
    InMux I__2606 (
            .O(N__12969),
            .I(N__12942));
    LocalMux I__2605 (
            .O(N__12966),
            .I(N__12937));
    LocalMux I__2604 (
            .O(N__12959),
            .I(N__12937));
    InMux I__2603 (
            .O(N__12956),
            .I(N__12934));
    InMux I__2602 (
            .O(N__12955),
            .I(N__12931));
    InMux I__2601 (
            .O(N__12954),
            .I(N__12928));
    LocalMux I__2600 (
            .O(N__12949),
            .I(N__12925));
    InMux I__2599 (
            .O(N__12948),
            .I(N__12918));
    InMux I__2598 (
            .O(N__12947),
            .I(N__12918));
    InMux I__2597 (
            .O(N__12946),
            .I(N__12918));
    InMux I__2596 (
            .O(N__12945),
            .I(N__12915));
    LocalMux I__2595 (
            .O(N__12942),
            .I(N__12910));
    Span4Mux_h I__2594 (
            .O(N__12937),
            .I(N__12910));
    LocalMux I__2593 (
            .O(N__12934),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2592 (
            .O(N__12931),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2591 (
            .O(N__12928),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__2590 (
            .O(N__12925),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2589 (
            .O(N__12918),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__2588 (
            .O(N__12915),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__2587 (
            .O(N__12910),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__2586 (
            .O(N__12895),
            .I(N__12889));
    InMux I__2585 (
            .O(N__12894),
            .I(N__12885));
    InMux I__2584 (
            .O(N__12893),
            .I(N__12869));
    InMux I__2583 (
            .O(N__12892),
            .I(N__12869));
    LocalMux I__2582 (
            .O(N__12889),
            .I(N__12861));
    InMux I__2581 (
            .O(N__12888),
            .I(N__12856));
    LocalMux I__2580 (
            .O(N__12885),
            .I(N__12853));
    InMux I__2579 (
            .O(N__12884),
            .I(N__12849));
    InMux I__2578 (
            .O(N__12883),
            .I(N__12846));
    InMux I__2577 (
            .O(N__12882),
            .I(N__12841));
    InMux I__2576 (
            .O(N__12881),
            .I(N__12841));
    InMux I__2575 (
            .O(N__12880),
            .I(N__12826));
    InMux I__2574 (
            .O(N__12879),
            .I(N__12826));
    InMux I__2573 (
            .O(N__12878),
            .I(N__12826));
    InMux I__2572 (
            .O(N__12877),
            .I(N__12826));
    InMux I__2571 (
            .O(N__12876),
            .I(N__12826));
    InMux I__2570 (
            .O(N__12875),
            .I(N__12826));
    InMux I__2569 (
            .O(N__12874),
            .I(N__12823));
    LocalMux I__2568 (
            .O(N__12869),
            .I(N__12820));
    InMux I__2567 (
            .O(N__12868),
            .I(N__12817));
    InMux I__2566 (
            .O(N__12867),
            .I(N__12810));
    InMux I__2565 (
            .O(N__12866),
            .I(N__12810));
    InMux I__2564 (
            .O(N__12865),
            .I(N__12810));
    InMux I__2563 (
            .O(N__12864),
            .I(N__12807));
    Span4Mux_h I__2562 (
            .O(N__12861),
            .I(N__12804));
    InMux I__2561 (
            .O(N__12860),
            .I(N__12799));
    InMux I__2560 (
            .O(N__12859),
            .I(N__12799));
    LocalMux I__2559 (
            .O(N__12856),
            .I(N__12794));
    Span4Mux_h I__2558 (
            .O(N__12853),
            .I(N__12794));
    InMux I__2557 (
            .O(N__12852),
            .I(N__12791));
    LocalMux I__2556 (
            .O(N__12849),
            .I(N__12784));
    LocalMux I__2555 (
            .O(N__12846),
            .I(N__12784));
    LocalMux I__2554 (
            .O(N__12841),
            .I(N__12784));
    InMux I__2553 (
            .O(N__12840),
            .I(N__12779));
    InMux I__2552 (
            .O(N__12839),
            .I(N__12779));
    LocalMux I__2551 (
            .O(N__12826),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2550 (
            .O(N__12823),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2549 (
            .O(N__12820),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2548 (
            .O(N__12817),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2547 (
            .O(N__12810),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2546 (
            .O(N__12807),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2545 (
            .O(N__12804),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2544 (
            .O(N__12799),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2543 (
            .O(N__12794),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2542 (
            .O(N__12791),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2541 (
            .O(N__12784),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2540 (
            .O(N__12779),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__2539 (
            .O(N__12754),
            .I(N__12751));
    LocalMux I__2538 (
            .O(N__12751),
            .I(\uu2.mem0.g1_0_1_1 ));
    InMux I__2537 (
            .O(N__12748),
            .I(N__12745));
    LocalMux I__2536 (
            .O(N__12745),
            .I(\uu2.mem0.g1_5_5 ));
    CascadeMux I__2535 (
            .O(N__12742),
            .I(N__12735));
    InMux I__2534 (
            .O(N__12741),
            .I(N__12730));
    InMux I__2533 (
            .O(N__12740),
            .I(N__12727));
    InMux I__2532 (
            .O(N__12739),
            .I(N__12720));
    InMux I__2531 (
            .O(N__12738),
            .I(N__12720));
    InMux I__2530 (
            .O(N__12735),
            .I(N__12720));
    InMux I__2529 (
            .O(N__12734),
            .I(N__12713));
    InMux I__2528 (
            .O(N__12733),
            .I(N__12710));
    LocalMux I__2527 (
            .O(N__12730),
            .I(N__12707));
    LocalMux I__2526 (
            .O(N__12727),
            .I(N__12704));
    LocalMux I__2525 (
            .O(N__12720),
            .I(N__12701));
    CascadeMux I__2524 (
            .O(N__12719),
            .I(N__12697));
    InMux I__2523 (
            .O(N__12718),
            .I(N__12689));
    InMux I__2522 (
            .O(N__12717),
            .I(N__12689));
    InMux I__2521 (
            .O(N__12716),
            .I(N__12689));
    LocalMux I__2520 (
            .O(N__12713),
            .I(N__12686));
    LocalMux I__2519 (
            .O(N__12710),
            .I(N__12677));
    Span4Mux_v I__2518 (
            .O(N__12707),
            .I(N__12677));
    Span4Mux_v I__2517 (
            .O(N__12704),
            .I(N__12677));
    Span4Mux_v I__2516 (
            .O(N__12701),
            .I(N__12677));
    InMux I__2515 (
            .O(N__12700),
            .I(N__12670));
    InMux I__2514 (
            .O(N__12697),
            .I(N__12670));
    InMux I__2513 (
            .O(N__12696),
            .I(N__12670));
    LocalMux I__2512 (
            .O(N__12689),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    Odrv4 I__2511 (
            .O(N__12686),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    Odrv4 I__2510 (
            .O(N__12677),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    LocalMux I__2509 (
            .O(N__12670),
            .I(\uu2.w_addr_displaying_3_repZ0Z2 ));
    InMux I__2508 (
            .O(N__12661),
            .I(N__12654));
    InMux I__2507 (
            .O(N__12660),
            .I(N__12654));
    CascadeMux I__2506 (
            .O(N__12659),
            .I(N__12650));
    LocalMux I__2505 (
            .O(N__12654),
            .I(N__12645));
    InMux I__2504 (
            .O(N__12653),
            .I(N__12642));
    InMux I__2503 (
            .O(N__12650),
            .I(N__12639));
    InMux I__2502 (
            .O(N__12649),
            .I(N__12634));
    InMux I__2501 (
            .O(N__12648),
            .I(N__12634));
    Span4Mux_v I__2500 (
            .O(N__12645),
            .I(N__12631));
    LocalMux I__2499 (
            .O(N__12642),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__2498 (
            .O(N__12639),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__2497 (
            .O(N__12634),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__2496 (
            .O(N__12631),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__2495 (
            .O(N__12622),
            .I(N__12619));
    InMux I__2494 (
            .O(N__12619),
            .I(N__12616));
    LocalMux I__2493 (
            .O(N__12616),
            .I(N__12613));
    Odrv12 I__2492 (
            .O(N__12613),
            .I(\uu2.mem0.N_74_i ));
    CascadeMux I__2491 (
            .O(N__12610),
            .I(N__12607));
    InMux I__2490 (
            .O(N__12607),
            .I(N__12604));
    LocalMux I__2489 (
            .O(N__12604),
            .I(\Lab_UT.dispString.dOutP_0_iv_3_0 ));
    CascadeMux I__2488 (
            .O(N__12601),
            .I(\uu2.N_84_cascade_ ));
    InMux I__2487 (
            .O(N__12598),
            .I(N__12589));
    InMux I__2486 (
            .O(N__12597),
            .I(N__12589));
    InMux I__2485 (
            .O(N__12596),
            .I(N__12589));
    LocalMux I__2484 (
            .O(N__12589),
            .I(N__12583));
    InMux I__2483 (
            .O(N__12588),
            .I(N__12573));
    InMux I__2482 (
            .O(N__12587),
            .I(N__12573));
    InMux I__2481 (
            .O(N__12586),
            .I(N__12573));
    Span4Mux_h I__2480 (
            .O(N__12583),
            .I(N__12570));
    InMux I__2479 (
            .O(N__12582),
            .I(N__12563));
    InMux I__2478 (
            .O(N__12581),
            .I(N__12563));
    InMux I__2477 (
            .O(N__12580),
            .I(N__12563));
    LocalMux I__2476 (
            .O(N__12573),
            .I(N__12560));
    Odrv4 I__2475 (
            .O(N__12570),
            .I(\uu2.N_97 ));
    LocalMux I__2474 (
            .O(N__12563),
            .I(\uu2.N_97 ));
    Odrv12 I__2473 (
            .O(N__12560),
            .I(\uu2.N_97 ));
    InMux I__2472 (
            .O(N__12553),
            .I(N__12549));
    CascadeMux I__2471 (
            .O(N__12552),
            .I(N__12545));
    LocalMux I__2470 (
            .O(N__12549),
            .I(N__12541));
    InMux I__2469 (
            .O(N__12548),
            .I(N__12533));
    InMux I__2468 (
            .O(N__12545),
            .I(N__12533));
    InMux I__2467 (
            .O(N__12544),
            .I(N__12533));
    Span4Mux_v I__2466 (
            .O(N__12541),
            .I(N__12530));
    InMux I__2465 (
            .O(N__12540),
            .I(N__12527));
    LocalMux I__2464 (
            .O(N__12533),
            .I(N__12520));
    Span4Mux_s3_h I__2463 (
            .O(N__12530),
            .I(N__12520));
    LocalMux I__2462 (
            .O(N__12527),
            .I(N__12520));
    Odrv4 I__2461 (
            .O(N__12520),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__2460 (
            .O(N__12517),
            .I(\uu2.N_97_cascade_ ));
    CascadeMux I__2459 (
            .O(N__12514),
            .I(N__12511));
    InMux I__2458 (
            .O(N__12511),
            .I(N__12506));
    InMux I__2457 (
            .O(N__12510),
            .I(N__12503));
    InMux I__2456 (
            .O(N__12509),
            .I(N__12500));
    LocalMux I__2455 (
            .O(N__12506),
            .I(N__12497));
    LocalMux I__2454 (
            .O(N__12503),
            .I(N__12494));
    LocalMux I__2453 (
            .O(N__12500),
            .I(\uu2.N_159 ));
    Odrv4 I__2452 (
            .O(N__12497),
            .I(\uu2.N_159 ));
    Odrv4 I__2451 (
            .O(N__12494),
            .I(\uu2.N_159 ));
    InMux I__2450 (
            .O(N__12487),
            .I(N__12478));
    InMux I__2449 (
            .O(N__12486),
            .I(N__12478));
    InMux I__2448 (
            .O(N__12485),
            .I(N__12478));
    LocalMux I__2447 (
            .O(N__12478),
            .I(N__12474));
    InMux I__2446 (
            .O(N__12477),
            .I(N__12471));
    Odrv4 I__2445 (
            .O(N__12474),
            .I(\uu2.un28_w_addr_user_i_0 ));
    LocalMux I__2444 (
            .O(N__12471),
            .I(\uu2.un28_w_addr_user_i_0 ));
    InMux I__2443 (
            .O(N__12466),
            .I(N__12463));
    LocalMux I__2442 (
            .O(N__12463),
            .I(N__12460));
    Span12Mux_s5_v I__2441 (
            .O(N__12460),
            .I(N__12454));
    InMux I__2440 (
            .O(N__12459),
            .I(N__12451));
    InMux I__2439 (
            .O(N__12458),
            .I(N__12446));
    InMux I__2438 (
            .O(N__12457),
            .I(N__12446));
    Odrv12 I__2437 (
            .O(N__12454),
            .I(L3_tx_data_0));
    LocalMux I__2436 (
            .O(N__12451),
            .I(L3_tx_data_0));
    LocalMux I__2435 (
            .O(N__12446),
            .I(L3_tx_data_0));
    InMux I__2434 (
            .O(N__12439),
            .I(N__12436));
    LocalMux I__2433 (
            .O(N__12436),
            .I(N__12432));
    CascadeMux I__2432 (
            .O(N__12435),
            .I(N__12429));
    Span4Mux_h I__2431 (
            .O(N__12432),
            .I(N__12426));
    InMux I__2430 (
            .O(N__12429),
            .I(N__12423));
    Span4Mux_h I__2429 (
            .O(N__12426),
            .I(N__12420));
    LocalMux I__2428 (
            .O(N__12423),
            .I(N__12417));
    Odrv4 I__2427 (
            .O(N__12420),
            .I(\uu2.N_86 ));
    Odrv12 I__2426 (
            .O(N__12417),
            .I(\uu2.N_86 ));
    InMux I__2425 (
            .O(N__12412),
            .I(N__12400));
    InMux I__2424 (
            .O(N__12411),
            .I(N__12400));
    InMux I__2423 (
            .O(N__12410),
            .I(N__12400));
    InMux I__2422 (
            .O(N__12409),
            .I(N__12400));
    LocalMux I__2421 (
            .O(N__12400),
            .I(N__12397));
    Span4Mux_h I__2420 (
            .O(N__12397),
            .I(N__12392));
    InMux I__2419 (
            .O(N__12396),
            .I(N__12387));
    InMux I__2418 (
            .O(N__12395),
            .I(N__12387));
    Odrv4 I__2417 (
            .O(N__12392),
            .I(L3_tx_data_rdy));
    LocalMux I__2416 (
            .O(N__12387),
            .I(L3_tx_data_rdy));
    CascadeMux I__2415 (
            .O(N__12382),
            .I(\uu2.N_86_cascade_ ));
    InMux I__2414 (
            .O(N__12379),
            .I(N__12373));
    InMux I__2413 (
            .O(N__12378),
            .I(N__12373));
    LocalMux I__2412 (
            .O(N__12373),
            .I(N__12370));
    Span4Mux_v I__2411 (
            .O(N__12370),
            .I(N__12367));
    Span4Mux_h I__2410 (
            .O(N__12367),
            .I(N__12362));
    InMux I__2409 (
            .O(N__12366),
            .I(N__12359));
    InMux I__2408 (
            .O(N__12365),
            .I(N__12356));
    Odrv4 I__2407 (
            .O(N__12362),
            .I(\uu2.N_84 ));
    LocalMux I__2406 (
            .O(N__12359),
            .I(\uu2.N_84 ));
    LocalMux I__2405 (
            .O(N__12356),
            .I(\uu2.N_84 ));
    CascadeMux I__2404 (
            .O(N__12349),
            .I(N__12345));
    CascadeMux I__2403 (
            .O(N__12348),
            .I(N__12340));
    InMux I__2402 (
            .O(N__12345),
            .I(N__12332));
    InMux I__2401 (
            .O(N__12344),
            .I(N__12332));
    InMux I__2400 (
            .O(N__12343),
            .I(N__12329));
    InMux I__2399 (
            .O(N__12340),
            .I(N__12324));
    InMux I__2398 (
            .O(N__12339),
            .I(N__12324));
    InMux I__2397 (
            .O(N__12338),
            .I(N__12318));
    InMux I__2396 (
            .O(N__12337),
            .I(N__12315));
    LocalMux I__2395 (
            .O(N__12332),
            .I(N__12308));
    LocalMux I__2394 (
            .O(N__12329),
            .I(N__12308));
    LocalMux I__2393 (
            .O(N__12324),
            .I(N__12308));
    InMux I__2392 (
            .O(N__12323),
            .I(N__12305));
    InMux I__2391 (
            .O(N__12322),
            .I(N__12302));
    InMux I__2390 (
            .O(N__12321),
            .I(N__12299));
    LocalMux I__2389 (
            .O(N__12318),
            .I(N__12296));
    LocalMux I__2388 (
            .O(N__12315),
            .I(N__12293));
    Span4Mux_v I__2387 (
            .O(N__12308),
            .I(N__12290));
    LocalMux I__2386 (
            .O(N__12305),
            .I(N__12283));
    LocalMux I__2385 (
            .O(N__12302),
            .I(N__12283));
    LocalMux I__2384 (
            .O(N__12299),
            .I(N__12283));
    Span4Mux_h I__2383 (
            .O(N__12296),
            .I(N__12277));
    Span4Mux_h I__2382 (
            .O(N__12293),
            .I(N__12270));
    Span4Mux_h I__2381 (
            .O(N__12290),
            .I(N__12270));
    Span4Mux_h I__2380 (
            .O(N__12283),
            .I(N__12270));
    InMux I__2379 (
            .O(N__12282),
            .I(N__12267));
    InMux I__2378 (
            .O(N__12281),
            .I(N__12262));
    InMux I__2377 (
            .O(N__12280),
            .I(N__12262));
    Odrv4 I__2376 (
            .O(N__12277),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    Odrv4 I__2375 (
            .O(N__12270),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    LocalMux I__2374 (
            .O(N__12267),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    LocalMux I__2373 (
            .O(N__12262),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    CascadeMux I__2372 (
            .O(N__12253),
            .I(\uu2.w_addr_i_0_tzZ0Z_0_cascade_ ));
    InMux I__2371 (
            .O(N__12250),
            .I(N__12247));
    LocalMux I__2370 (
            .O(N__12247),
            .I(N__12243));
    InMux I__2369 (
            .O(N__12246),
            .I(N__12240));
    Span4Mux_h I__2368 (
            .O(N__12243),
            .I(N__12236));
    LocalMux I__2367 (
            .O(N__12240),
            .I(N__12233));
    InMux I__2366 (
            .O(N__12239),
            .I(N__12230));
    Odrv4 I__2365 (
            .O(N__12236),
            .I(\uu2.N_61 ));
    Odrv12 I__2364 (
            .O(N__12233),
            .I(\uu2.N_61 ));
    LocalMux I__2363 (
            .O(N__12230),
            .I(\uu2.N_61 ));
    CascadeMux I__2362 (
            .O(N__12223),
            .I(N__12216));
    CascadeMux I__2361 (
            .O(N__12222),
            .I(N__12212));
    CascadeMux I__2360 (
            .O(N__12221),
            .I(N__12207));
    InMux I__2359 (
            .O(N__12220),
            .I(N__12201));
    InMux I__2358 (
            .O(N__12219),
            .I(N__12201));
    InMux I__2357 (
            .O(N__12216),
            .I(N__12198));
    InMux I__2356 (
            .O(N__12215),
            .I(N__12181));
    InMux I__2355 (
            .O(N__12212),
            .I(N__12181));
    InMux I__2354 (
            .O(N__12211),
            .I(N__12181));
    InMux I__2353 (
            .O(N__12210),
            .I(N__12181));
    InMux I__2352 (
            .O(N__12207),
            .I(N__12181));
    InMux I__2351 (
            .O(N__12206),
            .I(N__12181));
    LocalMux I__2350 (
            .O(N__12201),
            .I(N__12176));
    LocalMux I__2349 (
            .O(N__12198),
            .I(N__12176));
    InMux I__2348 (
            .O(N__12197),
            .I(N__12167));
    InMux I__2347 (
            .O(N__12196),
            .I(N__12167));
    InMux I__2346 (
            .O(N__12195),
            .I(N__12167));
    InMux I__2345 (
            .O(N__12194),
            .I(N__12167));
    LocalMux I__2344 (
            .O(N__12181),
            .I(N__12164));
    Span4Mux_v I__2343 (
            .O(N__12176),
            .I(N__12158));
    LocalMux I__2342 (
            .O(N__12167),
            .I(N__12158));
    Span4Mux_h I__2341 (
            .O(N__12164),
            .I(N__12155));
    InMux I__2340 (
            .O(N__12163),
            .I(N__12152));
    Odrv4 I__2339 (
            .O(N__12158),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__2338 (
            .O(N__12155),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__2337 (
            .O(N__12152),
            .I(\uu2.un21_w_addr_displaying_i ));
    InMux I__2336 (
            .O(N__12145),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    InMux I__2335 (
            .O(N__12142),
            .I(N__12139));
    LocalMux I__2334 (
            .O(N__12139),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ));
    CascadeMux I__2333 (
            .O(N__12136),
            .I(N__12130));
    InMux I__2332 (
            .O(N__12135),
            .I(N__12125));
    InMux I__2331 (
            .O(N__12134),
            .I(N__12125));
    InMux I__2330 (
            .O(N__12133),
            .I(N__12120));
    InMux I__2329 (
            .O(N__12130),
            .I(N__12120));
    LocalMux I__2328 (
            .O(N__12125),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2327 (
            .O(N__12120),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__2326 (
            .O(N__12115),
            .I(N__12109));
    InMux I__2325 (
            .O(N__12114),
            .I(N__12109));
    LocalMux I__2324 (
            .O(N__12109),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__2323 (
            .O(N__12106),
            .I(N__12102));
    InMux I__2322 (
            .O(N__12105),
            .I(N__12097));
    InMux I__2321 (
            .O(N__12102),
            .I(N__12097));
    LocalMux I__2320 (
            .O(N__12097),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__2319 (
            .O(N__12094),
            .I(N__12085));
    InMux I__2318 (
            .O(N__12093),
            .I(N__12085));
    InMux I__2317 (
            .O(N__12092),
            .I(N__12085));
    LocalMux I__2316 (
            .O(N__12085),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__2315 (
            .O(N__12082),
            .I(N__12077));
    CascadeMux I__2314 (
            .O(N__12081),
            .I(N__12074));
    InMux I__2313 (
            .O(N__12080),
            .I(N__12070));
    InMux I__2312 (
            .O(N__12077),
            .I(N__12063));
    InMux I__2311 (
            .O(N__12074),
            .I(N__12063));
    InMux I__2310 (
            .O(N__12073),
            .I(N__12063));
    LocalMux I__2309 (
            .O(N__12070),
            .I(\buart.Z_rx.ser_clk_2 ));
    LocalMux I__2308 (
            .O(N__12063),
            .I(\buart.Z_rx.ser_clk_2 ));
    InMux I__2307 (
            .O(N__12058),
            .I(N__12055));
    LocalMux I__2306 (
            .O(N__12055),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ));
    CascadeMux I__2305 (
            .O(N__12052),
            .I(N__12049));
    InMux I__2304 (
            .O(N__12049),
            .I(N__12042));
    InMux I__2303 (
            .O(N__12048),
            .I(N__12033));
    InMux I__2302 (
            .O(N__12047),
            .I(N__12033));
    InMux I__2301 (
            .O(N__12046),
            .I(N__12033));
    InMux I__2300 (
            .O(N__12045),
            .I(N__12033));
    LocalMux I__2299 (
            .O(N__12042),
            .I(\buart.Z_rx.ser_clk_3 ));
    LocalMux I__2298 (
            .O(N__12033),
            .I(\buart.Z_rx.ser_clk_3 ));
    InMux I__2297 (
            .O(N__12028),
            .I(N__12019));
    InMux I__2296 (
            .O(N__12027),
            .I(N__12019));
    InMux I__2295 (
            .O(N__12026),
            .I(N__12019));
    LocalMux I__2294 (
            .O(N__12019),
            .I(N__12013));
    InMux I__2293 (
            .O(N__12018),
            .I(N__12006));
    InMux I__2292 (
            .O(N__12017),
            .I(N__12006));
    InMux I__2291 (
            .O(N__12016),
            .I(N__12006));
    Span4Mux_v I__2290 (
            .O(N__12013),
            .I(N__11991));
    LocalMux I__2289 (
            .O(N__12006),
            .I(N__11991));
    InMux I__2288 (
            .O(N__12005),
            .I(N__11976));
    InMux I__2287 (
            .O(N__12004),
            .I(N__11976));
    InMux I__2286 (
            .O(N__12003),
            .I(N__11976));
    InMux I__2285 (
            .O(N__12002),
            .I(N__11976));
    InMux I__2284 (
            .O(N__12001),
            .I(N__11976));
    InMux I__2283 (
            .O(N__12000),
            .I(N__11976));
    InMux I__2282 (
            .O(N__11999),
            .I(N__11976));
    InMux I__2281 (
            .O(N__11998),
            .I(N__11971));
    InMux I__2280 (
            .O(N__11997),
            .I(N__11971));
    InMux I__2279 (
            .O(N__11996),
            .I(N__11968));
    Odrv4 I__2278 (
            .O(N__11991),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2277 (
            .O(N__11976),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2276 (
            .O(N__11971),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2275 (
            .O(N__11968),
            .I(\buart.Z_rx.startbit ));
    InMux I__2274 (
            .O(N__11959),
            .I(N__11953));
    InMux I__2273 (
            .O(N__11958),
            .I(N__11953));
    LocalMux I__2272 (
            .O(N__11953),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__2271 (
            .O(N__11950),
            .I(N__11947));
    LocalMux I__2270 (
            .O(N__11947),
            .I(N__11944));
    Span4Mux_v I__2269 (
            .O(N__11944),
            .I(N__11941));
    Odrv4 I__2268 (
            .O(N__11941),
            .I(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_2 ));
    InMux I__2267 (
            .O(N__11938),
            .I(N__11933));
    InMux I__2266 (
            .O(N__11937),
            .I(N__11927));
    InMux I__2265 (
            .O(N__11936),
            .I(N__11927));
    LocalMux I__2264 (
            .O(N__11933),
            .I(N__11924));
    InMux I__2263 (
            .O(N__11932),
            .I(N__11921));
    LocalMux I__2262 (
            .O(N__11927),
            .I(\uu2.w_addr_userZ0Z_3 ));
    Odrv4 I__2261 (
            .O(N__11924),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__2260 (
            .O(N__11921),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__2259 (
            .O(N__11914),
            .I(N__11907));
    InMux I__2258 (
            .O(N__11913),
            .I(N__11904));
    InMux I__2257 (
            .O(N__11912),
            .I(N__11899));
    InMux I__2256 (
            .O(N__11911),
            .I(N__11899));
    InMux I__2255 (
            .O(N__11910),
            .I(N__11896));
    InMux I__2254 (
            .O(N__11907),
            .I(N__11893));
    LocalMux I__2253 (
            .O(N__11904),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__2252 (
            .O(N__11899),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__2251 (
            .O(N__11896),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__2250 (
            .O(N__11893),
            .I(\uu2.w_addr_userZ0Z_5 ));
    InMux I__2249 (
            .O(N__11884),
            .I(N__11881));
    LocalMux I__2248 (
            .O(N__11881),
            .I(N__11875));
    InMux I__2247 (
            .O(N__11880),
            .I(N__11867));
    InMux I__2246 (
            .O(N__11879),
            .I(N__11867));
    InMux I__2245 (
            .O(N__11878),
            .I(N__11867));
    Span4Mux_h I__2244 (
            .O(N__11875),
            .I(N__11864));
    InMux I__2243 (
            .O(N__11874),
            .I(N__11861));
    LocalMux I__2242 (
            .O(N__11867),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__2241 (
            .O(N__11864),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__2240 (
            .O(N__11861),
            .I(\uu2.w_addr_userZ0Z_2 ));
    InMux I__2239 (
            .O(N__11854),
            .I(N__11851));
    LocalMux I__2238 (
            .O(N__11851),
            .I(\uu2.w_addr_user_3_i_a2_2_6 ));
    CascadeMux I__2237 (
            .O(N__11848),
            .I(N__11845));
    InMux I__2236 (
            .O(N__11845),
            .I(N__11842));
    LocalMux I__2235 (
            .O(N__11842),
            .I(N__11839));
    Span4Mux_h I__2234 (
            .O(N__11839),
            .I(N__11836));
    Odrv4 I__2233 (
            .O(N__11836),
            .I(\uu2.mem0.N_72_i ));
    CascadeMux I__2232 (
            .O(N__11833),
            .I(N__11830));
    InMux I__2231 (
            .O(N__11830),
            .I(N__11827));
    LocalMux I__2230 (
            .O(N__11827),
            .I(N__11822));
    InMux I__2229 (
            .O(N__11826),
            .I(N__11819));
    InMux I__2228 (
            .O(N__11825),
            .I(N__11816));
    Odrv4 I__2227 (
            .O(N__11822),
            .I(\buart.Z_rx.idle ));
    LocalMux I__2226 (
            .O(N__11819),
            .I(\buart.Z_rx.idle ));
    LocalMux I__2225 (
            .O(N__11816),
            .I(\buart.Z_rx.idle ));
    InMux I__2224 (
            .O(N__11809),
            .I(N__11806));
    LocalMux I__2223 (
            .O(N__11806),
            .I(N__11802));
    InMux I__2222 (
            .O(N__11805),
            .I(N__11799));
    Span4Mux_v I__2221 (
            .O(N__11802),
            .I(N__11796));
    LocalMux I__2220 (
            .O(N__11799),
            .I(N__11792));
    Span4Mux_v I__2219 (
            .O(N__11796),
            .I(N__11789));
    InMux I__2218 (
            .O(N__11795),
            .I(N__11786));
    Odrv4 I__2217 (
            .O(N__11792),
            .I(bu_rx_data_rdy));
    Odrv4 I__2216 (
            .O(N__11789),
            .I(bu_rx_data_rdy));
    LocalMux I__2215 (
            .O(N__11786),
            .I(bu_rx_data_rdy));
    CascadeMux I__2214 (
            .O(N__11779),
            .I(N__11776));
    InMux I__2213 (
            .O(N__11776),
            .I(N__11763));
    InMux I__2212 (
            .O(N__11775),
            .I(N__11763));
    InMux I__2211 (
            .O(N__11774),
            .I(N__11763));
    InMux I__2210 (
            .O(N__11773),
            .I(N__11763));
    InMux I__2209 (
            .O(N__11772),
            .I(N__11760));
    LocalMux I__2208 (
            .O(N__11763),
            .I(\buart.Z_rx.bitcountlde_0 ));
    LocalMux I__2207 (
            .O(N__11760),
            .I(\buart.Z_rx.bitcountlde_0 ));
    InMux I__2206 (
            .O(N__11755),
            .I(N__11752));
    LocalMux I__2205 (
            .O(N__11752),
            .I(\buart.Z_rx.un1_sample_0 ));
    CascadeMux I__2204 (
            .O(N__11749),
            .I(\buart.Z_rx.ser_clk_2_cascade_ ));
    CascadeMux I__2203 (
            .O(N__11746),
            .I(N__11740));
    InMux I__2202 (
            .O(N__11745),
            .I(N__11735));
    InMux I__2201 (
            .O(N__11744),
            .I(N__11730));
    InMux I__2200 (
            .O(N__11743),
            .I(N__11730));
    InMux I__2199 (
            .O(N__11740),
            .I(N__11727));
    InMux I__2198 (
            .O(N__11739),
            .I(N__11722));
    InMux I__2197 (
            .O(N__11738),
            .I(N__11722));
    LocalMux I__2196 (
            .O(N__11735),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2195 (
            .O(N__11730),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2194 (
            .O(N__11727),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2193 (
            .O(N__11722),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    CEMux I__2192 (
            .O(N__11713),
            .I(N__11709));
    CEMux I__2191 (
            .O(N__11712),
            .I(N__11706));
    LocalMux I__2190 (
            .O(N__11709),
            .I(N__11700));
    LocalMux I__2189 (
            .O(N__11706),
            .I(N__11700));
    CEMux I__2188 (
            .O(N__11705),
            .I(N__11697));
    Span4Mux_v I__2187 (
            .O(N__11700),
            .I(N__11694));
    LocalMux I__2186 (
            .O(N__11697),
            .I(N__11691));
    Sp12to4 I__2185 (
            .O(N__11694),
            .I(N__11688));
    Sp12to4 I__2184 (
            .O(N__11691),
            .I(N__11685));
    Span12Mux_s7_h I__2183 (
            .O(N__11688),
            .I(N__11680));
    Span12Mux_s7_v I__2182 (
            .O(N__11685),
            .I(N__11680));
    Odrv12 I__2181 (
            .O(N__11680),
            .I(\buart.Z_rx.sample ));
    InMux I__2180 (
            .O(N__11677),
            .I(N__11673));
    InMux I__2179 (
            .O(N__11676),
            .I(N__11670));
    LocalMux I__2178 (
            .O(N__11673),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__2177 (
            .O(N__11670),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__2176 (
            .O(N__11665),
            .I(N__11662));
    LocalMux I__2175 (
            .O(N__11662),
            .I(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ));
    InMux I__2174 (
            .O(N__11659),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__2173 (
            .O(N__11656),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__2172 (
            .O(N__11653),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    CascadeMux I__2171 (
            .O(N__11650),
            .I(N__11647));
    InMux I__2170 (
            .O(N__11647),
            .I(N__11644));
    LocalMux I__2169 (
            .O(N__11644),
            .I(N__11641));
    Odrv12 I__2168 (
            .O(N__11641),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    CascadeMux I__2167 (
            .O(N__11638),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ));
    InMux I__2166 (
            .O(N__11635),
            .I(N__11632));
    LocalMux I__2165 (
            .O(N__11632),
            .I(N__11629));
    Span4Mux_h I__2164 (
            .O(N__11629),
            .I(N__11626));
    Span4Mux_v I__2163 (
            .O(N__11626),
            .I(N__11622));
    InMux I__2162 (
            .O(N__11625),
            .I(N__11619));
    Odrv4 I__2161 (
            .O(N__11622),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    LocalMux I__2160 (
            .O(N__11619),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    InMux I__2159 (
            .O(N__11614),
            .I(N__11611));
    LocalMux I__2158 (
            .O(N__11611),
            .I(\Lab_UT.dictrl.next_state_out_0 ));
    CascadeMux I__2157 (
            .O(N__11608),
            .I(\Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_ ));
    CascadeMux I__2156 (
            .O(N__11605),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ));
    InMux I__2155 (
            .O(N__11602),
            .I(N__11599));
    LocalMux I__2154 (
            .O(N__11599),
            .I(N__11596));
    Span12Mux_s8_v I__2153 (
            .O(N__11596),
            .I(N__11593));
    Odrv12 I__2152 (
            .O(N__11593),
            .I(\Lab_UT.dictrl.dicRun_2_reti ));
    InMux I__2151 (
            .O(N__11590),
            .I(N__11587));
    LocalMux I__2150 (
            .O(N__11587),
            .I(N__11583));
    InMux I__2149 (
            .O(N__11586),
            .I(N__11580));
    Odrv4 I__2148 (
            .O(N__11583),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_1 ));
    LocalMux I__2147 (
            .O(N__11580),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_1 ));
    CascadeMux I__2146 (
            .O(N__11575),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_cascade_ ));
    CascadeMux I__2145 (
            .O(N__11572),
            .I(\Lab_UT.m37_ns_cascade_ ));
    InMux I__2144 (
            .O(N__11569),
            .I(N__11566));
    LocalMux I__2143 (
            .O(N__11566),
            .I(\Lab_UT.dictrl.next_state_out_2 ));
    SRMux I__2142 (
            .O(N__11563),
            .I(N__11560));
    LocalMux I__2141 (
            .O(N__11560),
            .I(N__11556));
    InMux I__2140 (
            .O(N__11559),
            .I(N__11553));
    Span4Mux_h I__2139 (
            .O(N__11556),
            .I(N__11550));
    LocalMux I__2138 (
            .O(N__11553),
            .I(N__11547));
    Odrv4 I__2137 (
            .O(N__11550),
            .I(\Lab_UT.m45 ));
    Odrv4 I__2136 (
            .O(N__11547),
            .I(\Lab_UT.m45 ));
    CascadeMux I__2135 (
            .O(N__11542),
            .I(\Lab_UT.m40_cascade_ ));
    CascadeMux I__2134 (
            .O(N__11539),
            .I(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_ ));
    CascadeMux I__2133 (
            .O(N__11536),
            .I(resetGen_escKey_4_cascade_));
    InMux I__2132 (
            .O(N__11533),
            .I(N__11525));
    InMux I__2131 (
            .O(N__11532),
            .I(N__11525));
    CascadeMux I__2130 (
            .O(N__11531),
            .I(N__11521));
    InMux I__2129 (
            .O(N__11530),
            .I(N__11518));
    LocalMux I__2128 (
            .O(N__11525),
            .I(N__11515));
    InMux I__2127 (
            .O(N__11524),
            .I(N__11510));
    InMux I__2126 (
            .O(N__11521),
            .I(N__11510));
    LocalMux I__2125 (
            .O(N__11518),
            .I(N__11505));
    Span4Mux_v I__2124 (
            .O(N__11515),
            .I(N__11505));
    LocalMux I__2123 (
            .O(N__11510),
            .I(bu_rx_data_5));
    Odrv4 I__2122 (
            .O(N__11505),
            .I(bu_rx_data_5));
    CascadeMux I__2121 (
            .O(N__11500),
            .I(N__11494));
    InMux I__2120 (
            .O(N__11499),
            .I(N__11488));
    InMux I__2119 (
            .O(N__11498),
            .I(N__11485));
    InMux I__2118 (
            .O(N__11497),
            .I(N__11474));
    InMux I__2117 (
            .O(N__11494),
            .I(N__11474));
    InMux I__2116 (
            .O(N__11493),
            .I(N__11474));
    InMux I__2115 (
            .O(N__11492),
            .I(N__11474));
    InMux I__2114 (
            .O(N__11491),
            .I(N__11474));
    LocalMux I__2113 (
            .O(N__11488),
            .I(bu_rx_data_2));
    LocalMux I__2112 (
            .O(N__11485),
            .I(bu_rx_data_2));
    LocalMux I__2111 (
            .O(N__11474),
            .I(bu_rx_data_2));
    CascadeMux I__2110 (
            .O(N__11467),
            .I(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_ ));
    InMux I__2109 (
            .O(N__11464),
            .I(N__11456));
    InMux I__2108 (
            .O(N__11463),
            .I(N__11445));
    InMux I__2107 (
            .O(N__11462),
            .I(N__11445));
    InMux I__2106 (
            .O(N__11461),
            .I(N__11445));
    InMux I__2105 (
            .O(N__11460),
            .I(N__11445));
    InMux I__2104 (
            .O(N__11459),
            .I(N__11445));
    LocalMux I__2103 (
            .O(N__11456),
            .I(bu_rx_data_4));
    LocalMux I__2102 (
            .O(N__11445),
            .I(bu_rx_data_4));
    CascadeMux I__2101 (
            .O(N__11440),
            .I(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ));
    InMux I__2100 (
            .O(N__11437),
            .I(N__11434));
    LocalMux I__2099 (
            .O(N__11434),
            .I(resetGen_escKey_2_0));
    InMux I__2098 (
            .O(N__11431),
            .I(N__11423));
    InMux I__2097 (
            .O(N__11430),
            .I(N__11423));
    CascadeMux I__2096 (
            .O(N__11429),
            .I(N__11420));
    InMux I__2095 (
            .O(N__11428),
            .I(N__11416));
    LocalMux I__2094 (
            .O(N__11423),
            .I(N__11413));
    InMux I__2093 (
            .O(N__11420),
            .I(N__11408));
    InMux I__2092 (
            .O(N__11419),
            .I(N__11408));
    LocalMux I__2091 (
            .O(N__11416),
            .I(N__11401));
    Span4Mux_v I__2090 (
            .O(N__11413),
            .I(N__11401));
    LocalMux I__2089 (
            .O(N__11408),
            .I(N__11401));
    Odrv4 I__2088 (
            .O(N__11401),
            .I(bu_rx_data_6));
    CascadeMux I__2087 (
            .O(N__11398),
            .I(N__11391));
    CascadeMux I__2086 (
            .O(N__11397),
            .I(N__11388));
    InMux I__2085 (
            .O(N__11396),
            .I(N__11383));
    InMux I__2084 (
            .O(N__11395),
            .I(N__11374));
    InMux I__2083 (
            .O(N__11394),
            .I(N__11374));
    InMux I__2082 (
            .O(N__11391),
            .I(N__11374));
    InMux I__2081 (
            .O(N__11388),
            .I(N__11374));
    InMux I__2080 (
            .O(N__11387),
            .I(N__11369));
    InMux I__2079 (
            .O(N__11386),
            .I(N__11369));
    LocalMux I__2078 (
            .O(N__11383),
            .I(bu_rx_data_3));
    LocalMux I__2077 (
            .O(N__11374),
            .I(bu_rx_data_3));
    LocalMux I__2076 (
            .O(N__11369),
            .I(bu_rx_data_3));
    CascadeMux I__2075 (
            .O(N__11362),
            .I(N__11358));
    InMux I__2074 (
            .O(N__11361),
            .I(N__11352));
    InMux I__2073 (
            .O(N__11358),
            .I(N__11352));
    CascadeMux I__2072 (
            .O(N__11357),
            .I(N__11348));
    LocalMux I__2071 (
            .O(N__11352),
            .I(N__11344));
    InMux I__2070 (
            .O(N__11351),
            .I(N__11339));
    InMux I__2069 (
            .O(N__11348),
            .I(N__11339));
    InMux I__2068 (
            .O(N__11347),
            .I(N__11336));
    Span4Mux_h I__2067 (
            .O(N__11344),
            .I(N__11333));
    LocalMux I__2066 (
            .O(N__11339),
            .I(N__11330));
    LocalMux I__2065 (
            .O(N__11336),
            .I(bu_rx_data_7));
    Odrv4 I__2064 (
            .O(N__11333),
            .I(bu_rx_data_7));
    Odrv12 I__2063 (
            .O(N__11330),
            .I(bu_rx_data_7));
    InMux I__2062 (
            .O(N__11323),
            .I(N__11320));
    LocalMux I__2061 (
            .O(N__11320),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxa_2 ));
    CascadeMux I__2060 (
            .O(N__11317),
            .I(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_ ));
    InMux I__2059 (
            .O(N__11314),
            .I(N__11311));
    LocalMux I__2058 (
            .O(N__11311),
            .I(N__11308));
    Span4Mux_v I__2057 (
            .O(N__11308),
            .I(N__11305));
    Odrv4 I__2056 (
            .O(N__11305),
            .I(\Lab_UT.didp.countrce2.N_183 ));
    InMux I__2055 (
            .O(N__11302),
            .I(N__11299));
    LocalMux I__2054 (
            .O(N__11299),
            .I(\Lab_UT.didp.countrce2.N_180 ));
    CascadeMux I__2053 (
            .O(N__11296),
            .I(\Lab_UT.didp.countrce4.N_80_i_cascade_ ));
    InMux I__2052 (
            .O(N__11293),
            .I(N__11290));
    LocalMux I__2051 (
            .O(N__11290),
            .I(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_3 ));
    InMux I__2050 (
            .O(N__11287),
            .I(N__11284));
    LocalMux I__2049 (
            .O(N__11284),
            .I(\Lab_UT.bcd2segment4.segment_i_0Z0Z_6 ));
    InMux I__2048 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__2047 (
            .O(N__11278),
            .I(\Lab_UT.dictrl.next_alarmstate4_1Z0Z_0 ));
    CascadeMux I__2046 (
            .O(N__11275),
            .I(\Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_ ));
    InMux I__2045 (
            .O(N__11272),
            .I(N__11269));
    LocalMux I__2044 (
            .O(N__11269),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__2043 (
            .O(N__11266),
            .I(N__11259));
    InMux I__2042 (
            .O(N__11265),
            .I(N__11253));
    InMux I__2041 (
            .O(N__11264),
            .I(N__11250));
    InMux I__2040 (
            .O(N__11263),
            .I(N__11247));
    InMux I__2039 (
            .O(N__11262),
            .I(N__11244));
    LocalMux I__2038 (
            .O(N__11259),
            .I(N__11241));
    InMux I__2037 (
            .O(N__11258),
            .I(N__11234));
    InMux I__2036 (
            .O(N__11257),
            .I(N__11234));
    InMux I__2035 (
            .O(N__11256),
            .I(N__11234));
    LocalMux I__2034 (
            .O(N__11253),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2033 (
            .O(N__11250),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2032 (
            .O(N__11247),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2031 (
            .O(N__11244),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    Odrv4 I__2030 (
            .O(N__11241),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__2029 (
            .O(N__11234),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    CascadeMux I__2028 (
            .O(N__11221),
            .I(\uu2.N_7_cascade_ ));
    CascadeMux I__2027 (
            .O(N__11218),
            .I(N__11215));
    InMux I__2026 (
            .O(N__11215),
            .I(N__11212));
    LocalMux I__2025 (
            .O(N__11212),
            .I(N__11209));
    Odrv4 I__2024 (
            .O(N__11209),
            .I(\uu2.N_10 ));
    InMux I__2023 (
            .O(N__11206),
            .I(N__11202));
    InMux I__2022 (
            .O(N__11205),
            .I(N__11195));
    LocalMux I__2021 (
            .O(N__11202),
            .I(N__11192));
    InMux I__2020 (
            .O(N__11201),
            .I(N__11187));
    InMux I__2019 (
            .O(N__11200),
            .I(N__11187));
    InMux I__2018 (
            .O(N__11199),
            .I(N__11182));
    InMux I__2017 (
            .O(N__11198),
            .I(N__11182));
    LocalMux I__2016 (
            .O(N__11195),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__2015 (
            .O(N__11192),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__2014 (
            .O(N__11187),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__2013 (
            .O(N__11182),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    InMux I__2012 (
            .O(N__11173),
            .I(N__11170));
    LocalMux I__2011 (
            .O(N__11170),
            .I(\uu2.N_8 ));
    InMux I__2010 (
            .O(N__11167),
            .I(N__11164));
    LocalMux I__2009 (
            .O(N__11164),
            .I(\uu2.bitmapZ0Z_84 ));
    InMux I__2008 (
            .O(N__11161),
            .I(N__11158));
    LocalMux I__2007 (
            .O(N__11158),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__2006 (
            .O(N__11155),
            .I(N__11152));
    LocalMux I__2005 (
            .O(N__11152),
            .I(\Lab_UT.didp.countrce2.N_178 ));
    InMux I__2004 (
            .O(N__11149),
            .I(N__11146));
    LocalMux I__2003 (
            .O(N__11146),
            .I(N__11143));
    Odrv12 I__2002 (
            .O(N__11143),
            .I(\Lab_UT.didp.countrce2.N_175 ));
    InMux I__2001 (
            .O(N__11140),
            .I(N__11137));
    LocalMux I__2000 (
            .O(N__11137),
            .I(N__11134));
    Span4Mux_h I__1999 (
            .O(N__11134),
            .I(N__11131));
    Odrv4 I__1998 (
            .O(N__11131),
            .I(\Lab_UT.didp.countrce2.N_170 ));
    CascadeMux I__1997 (
            .O(N__11128),
            .I(\uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_ ));
    InMux I__1996 (
            .O(N__11125),
            .I(N__11122));
    LocalMux I__1995 (
            .O(N__11122),
            .I(N__11119));
    Odrv4 I__1994 (
            .O(N__11119),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_45 ));
    InMux I__1993 (
            .O(N__11116),
            .I(N__11106));
    InMux I__1992 (
            .O(N__11115),
            .I(N__11103));
    InMux I__1991 (
            .O(N__11114),
            .I(N__11100));
    InMux I__1990 (
            .O(N__11113),
            .I(N__11095));
    InMux I__1989 (
            .O(N__11112),
            .I(N__11095));
    InMux I__1988 (
            .O(N__11111),
            .I(N__11090));
    InMux I__1987 (
            .O(N__11110),
            .I(N__11090));
    InMux I__1986 (
            .O(N__11109),
            .I(N__11087));
    LocalMux I__1985 (
            .O(N__11106),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1984 (
            .O(N__11103),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1983 (
            .O(N__11100),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1982 (
            .O(N__11095),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1981 (
            .O(N__11090),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    LocalMux I__1980 (
            .O(N__11087),
            .I(\uu2.w_addr_displaying_2_repZ0Z1 ));
    CascadeMux I__1979 (
            .O(N__11074),
            .I(N__11071));
    InMux I__1978 (
            .O(N__11071),
            .I(N__11068));
    LocalMux I__1977 (
            .O(N__11068),
            .I(N__11060));
    InMux I__1976 (
            .O(N__11067),
            .I(N__11054));
    InMux I__1975 (
            .O(N__11066),
            .I(N__11051));
    InMux I__1974 (
            .O(N__11065),
            .I(N__11048));
    InMux I__1973 (
            .O(N__11064),
            .I(N__11045));
    InMux I__1972 (
            .O(N__11063),
            .I(N__11042));
    Span4Mux_h I__1971 (
            .O(N__11060),
            .I(N__11039));
    InMux I__1970 (
            .O(N__11059),
            .I(N__11032));
    InMux I__1969 (
            .O(N__11058),
            .I(N__11032));
    InMux I__1968 (
            .O(N__11057),
            .I(N__11032));
    LocalMux I__1967 (
            .O(N__11054),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1966 (
            .O(N__11051),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1965 (
            .O(N__11048),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1964 (
            .O(N__11045),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1963 (
            .O(N__11042),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__1962 (
            .O(N__11039),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__1961 (
            .O(N__11032),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__1960 (
            .O(N__11017),
            .I(N__11014));
    LocalMux I__1959 (
            .O(N__11014),
            .I(\uu2.bitmap_pmux_sn_N_31_0 ));
    CascadeMux I__1958 (
            .O(N__11011),
            .I(\uu2.bitmap_pmux_sn_N_31_0_cascade_ ));
    InMux I__1957 (
            .O(N__11008),
            .I(N__10999));
    InMux I__1956 (
            .O(N__11007),
            .I(N__10999));
    InMux I__1955 (
            .O(N__11006),
            .I(N__10999));
    LocalMux I__1954 (
            .O(N__10999),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    InMux I__1953 (
            .O(N__10996),
            .I(N__10993));
    LocalMux I__1952 (
            .O(N__10993),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_48 ));
    CascadeMux I__1951 (
            .O(N__10990),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_ ));
    InMux I__1950 (
            .O(N__10987),
            .I(N__10984));
    LocalMux I__1949 (
            .O(N__10984),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_47 ));
    InMux I__1948 (
            .O(N__10981),
            .I(N__10978));
    LocalMux I__1947 (
            .O(N__10978),
            .I(N__10975));
    Odrv4 I__1946 (
            .O(N__10975),
            .I(\uu2.mem0.bitmap_pmux_u_ns_1 ));
    CascadeMux I__1945 (
            .O(N__10972),
            .I(\uu2.mem0.g0_5_3_cascade_ ));
    InMux I__1944 (
            .O(N__10969),
            .I(N__10966));
    LocalMux I__1943 (
            .O(N__10966),
            .I(\uu2.mem0.g0_5_6 ));
    CascadeMux I__1942 (
            .O(N__10963),
            .I(\Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_ ));
    CascadeMux I__1941 (
            .O(N__10960),
            .I(\uu2.un31_w_data_displaying_0_a2_1_cascade_ ));
    InMux I__1940 (
            .O(N__10957),
            .I(N__10950));
    InMux I__1939 (
            .O(N__10956),
            .I(N__10950));
    InMux I__1938 (
            .O(N__10955),
            .I(N__10947));
    LocalMux I__1937 (
            .O(N__10950),
            .I(N__10944));
    LocalMux I__1936 (
            .O(N__10947),
            .I(N__10941));
    Span4Mux_v I__1935 (
            .O(N__10944),
            .I(N__10936));
    Span4Mux_v I__1934 (
            .O(N__10941),
            .I(N__10936));
    Odrv4 I__1933 (
            .O(N__10936),
            .I(\uu2.un31_w_data_displaying ));
    InMux I__1932 (
            .O(N__10933),
            .I(N__10930));
    LocalMux I__1931 (
            .O(N__10930),
            .I(\uu2.un15_w_data_displaying_6 ));
    CascadeMux I__1930 (
            .O(N__10927),
            .I(\uu2.un15_w_data_displaying_6_cascade_ ));
    InMux I__1929 (
            .O(N__10924),
            .I(N__10920));
    InMux I__1928 (
            .O(N__10923),
            .I(N__10917));
    LocalMux I__1927 (
            .O(N__10920),
            .I(N__10912));
    LocalMux I__1926 (
            .O(N__10917),
            .I(N__10912));
    Odrv4 I__1925 (
            .O(N__10912),
            .I(\uu2.un49_w_data_displaying_1 ));
    InMux I__1924 (
            .O(N__10909),
            .I(N__10905));
    InMux I__1923 (
            .O(N__10908),
            .I(N__10902));
    LocalMux I__1922 (
            .O(N__10905),
            .I(N__10899));
    LocalMux I__1921 (
            .O(N__10902),
            .I(N__10896));
    Span4Mux_h I__1920 (
            .O(N__10899),
            .I(N__10893));
    Span4Mux_h I__1919 (
            .O(N__10896),
            .I(N__10890));
    Odrv4 I__1918 (
            .O(N__10893),
            .I(\uu2.un49_w_data_displaying ));
    Odrv4 I__1917 (
            .O(N__10890),
            .I(\uu2.un49_w_data_displaying ));
    CascadeMux I__1916 (
            .O(N__10885),
            .I(N__10881));
    InMux I__1915 (
            .O(N__10884),
            .I(N__10877));
    InMux I__1914 (
            .O(N__10881),
            .I(N__10872));
    InMux I__1913 (
            .O(N__10880),
            .I(N__10872));
    LocalMux I__1912 (
            .O(N__10877),
            .I(N__10869));
    LocalMux I__1911 (
            .O(N__10872),
            .I(N__10864));
    Span4Mux_h I__1910 (
            .O(N__10869),
            .I(N__10864));
    Odrv4 I__1909 (
            .O(N__10864),
            .I(\uu2.un15_w_data_displaying_i_i_o2_0 ));
    CascadeMux I__1908 (
            .O(N__10861),
            .I(\uu2.un15_w_data_displaying_i_i_o2_0_cascade_ ));
    InMux I__1907 (
            .O(N__10858),
            .I(N__10855));
    LocalMux I__1906 (
            .O(N__10855),
            .I(\uu2.mem0.un49_w_data_displaying_0 ));
    CascadeMux I__1905 (
            .O(N__10852),
            .I(N__10849));
    InMux I__1904 (
            .O(N__10849),
            .I(N__10846));
    LocalMux I__1903 (
            .O(N__10846),
            .I(N__10843));
    Odrv4 I__1902 (
            .O(N__10843),
            .I(\uu2.mem0.g0_5_5 ));
    InMux I__1901 (
            .O(N__10840),
            .I(N__10837));
    LocalMux I__1900 (
            .O(N__10837),
            .I(\uu2.mem0.un31_w_data_displaying_0 ));
    InMux I__1899 (
            .O(N__10834),
            .I(N__10831));
    LocalMux I__1898 (
            .O(N__10831),
            .I(N__10828));
    Span4Mux_h I__1897 (
            .O(N__10828),
            .I(N__10825));
    Odrv4 I__1896 (
            .O(N__10825),
            .I(\uu2.mem0.g1_1_1 ));
    InMux I__1895 (
            .O(N__10822),
            .I(N__10818));
    InMux I__1894 (
            .O(N__10821),
            .I(N__10815));
    LocalMux I__1893 (
            .O(N__10818),
            .I(N__10810));
    LocalMux I__1892 (
            .O(N__10815),
            .I(N__10807));
    CascadeMux I__1891 (
            .O(N__10814),
            .I(N__10800));
    InMux I__1890 (
            .O(N__10813),
            .I(N__10796));
    Span4Mux_h I__1889 (
            .O(N__10810),
            .I(N__10791));
    Span4Mux_h I__1888 (
            .O(N__10807),
            .I(N__10791));
    InMux I__1887 (
            .O(N__10806),
            .I(N__10788));
    InMux I__1886 (
            .O(N__10805),
            .I(N__10783));
    InMux I__1885 (
            .O(N__10804),
            .I(N__10783));
    InMux I__1884 (
            .O(N__10803),
            .I(N__10776));
    InMux I__1883 (
            .O(N__10800),
            .I(N__10776));
    InMux I__1882 (
            .O(N__10799),
            .I(N__10776));
    LocalMux I__1881 (
            .O(N__10796),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    Odrv4 I__1880 (
            .O(N__10791),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1879 (
            .O(N__10788),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1878 (
            .O(N__10783),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    LocalMux I__1877 (
            .O(N__10776),
            .I(\uu2.w_addr_displaying_7_repZ0Z1 ));
    InMux I__1876 (
            .O(N__10765),
            .I(N__10753));
    InMux I__1875 (
            .O(N__10764),
            .I(N__10753));
    InMux I__1874 (
            .O(N__10763),
            .I(N__10748));
    InMux I__1873 (
            .O(N__10762),
            .I(N__10748));
    InMux I__1872 (
            .O(N__10761),
            .I(N__10745));
    InMux I__1871 (
            .O(N__10760),
            .I(N__10742));
    InMux I__1870 (
            .O(N__10759),
            .I(N__10737));
    InMux I__1869 (
            .O(N__10758),
            .I(N__10737));
    LocalMux I__1868 (
            .O(N__10753),
            .I(N__10734));
    LocalMux I__1867 (
            .O(N__10748),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1866 (
            .O(N__10745),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1865 (
            .O(N__10742),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    LocalMux I__1864 (
            .O(N__10737),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    Odrv4 I__1863 (
            .O(N__10734),
            .I(\uu2.w_addr_displaying_8_repZ0Z1 ));
    InMux I__1862 (
            .O(N__10723),
            .I(N__10720));
    LocalMux I__1861 (
            .O(N__10720),
            .I(N__10711));
    InMux I__1860 (
            .O(N__10719),
            .I(N__10704));
    InMux I__1859 (
            .O(N__10718),
            .I(N__10704));
    InMux I__1858 (
            .O(N__10717),
            .I(N__10704));
    InMux I__1857 (
            .O(N__10716),
            .I(N__10701));
    InMux I__1856 (
            .O(N__10715),
            .I(N__10696));
    InMux I__1855 (
            .O(N__10714),
            .I(N__10696));
    Odrv4 I__1854 (
            .O(N__10711),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1853 (
            .O(N__10704),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1852 (
            .O(N__10701),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1851 (
            .O(N__10696),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__1850 (
            .O(N__10687),
            .I(N__10679));
    InMux I__1849 (
            .O(N__10686),
            .I(N__10676));
    CascadeMux I__1848 (
            .O(N__10685),
            .I(N__10673));
    CascadeMux I__1847 (
            .O(N__10684),
            .I(N__10670));
    CascadeMux I__1846 (
            .O(N__10683),
            .I(N__10667));
    CascadeMux I__1845 (
            .O(N__10682),
            .I(N__10664));
    InMux I__1844 (
            .O(N__10679),
            .I(N__10661));
    LocalMux I__1843 (
            .O(N__10676),
            .I(N__10658));
    InMux I__1842 (
            .O(N__10673),
            .I(N__10655));
    InMux I__1841 (
            .O(N__10670),
            .I(N__10648));
    InMux I__1840 (
            .O(N__10667),
            .I(N__10648));
    InMux I__1839 (
            .O(N__10664),
            .I(N__10648));
    LocalMux I__1838 (
            .O(N__10661),
            .I(N__10645));
    Span4Mux_h I__1837 (
            .O(N__10658),
            .I(N__10642));
    LocalMux I__1836 (
            .O(N__10655),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__1835 (
            .O(N__10648),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1834 (
            .O(N__10645),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1833 (
            .O(N__10642),
            .I(\uu2.w_addr_userZ0Z_1 ));
    InMux I__1832 (
            .O(N__10633),
            .I(N__10630));
    LocalMux I__1831 (
            .O(N__10630),
            .I(N__10627));
    Span4Mux_h I__1830 (
            .O(N__10627),
            .I(N__10624));
    Odrv4 I__1829 (
            .O(N__10624),
            .I(\uu2.mem0.N_111 ));
    CEMux I__1828 (
            .O(N__10621),
            .I(N__10618));
    LocalMux I__1827 (
            .O(N__10618),
            .I(N__10614));
    CEMux I__1826 (
            .O(N__10617),
            .I(N__10611));
    Span4Mux_h I__1825 (
            .O(N__10614),
            .I(N__10608));
    LocalMux I__1824 (
            .O(N__10611),
            .I(N__10605));
    Odrv4 I__1823 (
            .O(N__10608),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    Odrv12 I__1822 (
            .O(N__10605),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    CascadeMux I__1821 (
            .O(N__10600),
            .I(N__10597));
    InMux I__1820 (
            .O(N__10597),
            .I(N__10594));
    LocalMux I__1819 (
            .O(N__10594),
            .I(N__10591));
    Span4Mux_h I__1818 (
            .O(N__10591),
            .I(N__10588));
    Odrv4 I__1817 (
            .O(N__10588),
            .I(\uu2.mem0.N_73_i ));
    CascadeMux I__1816 (
            .O(N__10585),
            .I(\buart.Z_rx.bitcount_lm_2_cascade_ ));
    InMux I__1815 (
            .O(N__10582),
            .I(N__10572));
    InMux I__1814 (
            .O(N__10581),
            .I(N__10572));
    InMux I__1813 (
            .O(N__10580),
            .I(N__10569));
    InMux I__1812 (
            .O(N__10579),
            .I(N__10566));
    InMux I__1811 (
            .O(N__10578),
            .I(N__10561));
    InMux I__1810 (
            .O(N__10577),
            .I(N__10561));
    LocalMux I__1809 (
            .O(N__10572),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1808 (
            .O(N__10569),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1807 (
            .O(N__10566),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1806 (
            .O(N__10561),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    InMux I__1805 (
            .O(N__10552),
            .I(N__10549));
    LocalMux I__1804 (
            .O(N__10549),
            .I(\buart.Z_rx.bitcount_lm_4 ));
    InMux I__1803 (
            .O(N__10546),
            .I(N__10539));
    InMux I__1802 (
            .O(N__10545),
            .I(N__10536));
    InMux I__1801 (
            .O(N__10544),
            .I(N__10533));
    InMux I__1800 (
            .O(N__10543),
            .I(N__10528));
    InMux I__1799 (
            .O(N__10542),
            .I(N__10528));
    LocalMux I__1798 (
            .O(N__10539),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1797 (
            .O(N__10536),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1796 (
            .O(N__10533),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1795 (
            .O(N__10528),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__1794 (
            .O(N__10519),
            .I(N__10516));
    InMux I__1793 (
            .O(N__10516),
            .I(N__10513));
    LocalMux I__1792 (
            .O(N__10513),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__1791 (
            .O(N__10510),
            .I(N__10504));
    InMux I__1790 (
            .O(N__10509),
            .I(N__10497));
    InMux I__1789 (
            .O(N__10508),
            .I(N__10497));
    InMux I__1788 (
            .O(N__10507),
            .I(N__10497));
    InMux I__1787 (
            .O(N__10504),
            .I(N__10494));
    LocalMux I__1786 (
            .O(N__10497),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1785 (
            .O(N__10494),
            .I(\buart.Z_rx.N_27_0_i ));
    CascadeMux I__1784 (
            .O(N__10489),
            .I(\buart.Z_rx.bitcount_lm_3_cascade_ ));
    InMux I__1783 (
            .O(N__10486),
            .I(N__10476));
    InMux I__1782 (
            .O(N__10485),
            .I(N__10476));
    InMux I__1781 (
            .O(N__10484),
            .I(N__10473));
    InMux I__1780 (
            .O(N__10483),
            .I(N__10470));
    InMux I__1779 (
            .O(N__10482),
            .I(N__10465));
    InMux I__1778 (
            .O(N__10481),
            .I(N__10465));
    LocalMux I__1777 (
            .O(N__10476),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1776 (
            .O(N__10473),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1775 (
            .O(N__10470),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1774 (
            .O(N__10465),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    InMux I__1773 (
            .O(N__10456),
            .I(N__10453));
    LocalMux I__1772 (
            .O(N__10453),
            .I(\uu2.N_153 ));
    CascadeMux I__1771 (
            .O(N__10450),
            .I(\uu2.N_90_cascade_ ));
    InMux I__1770 (
            .O(N__10447),
            .I(N__10444));
    LocalMux I__1769 (
            .O(N__10444),
            .I(\uu2.N_105 ));
    CascadeMux I__1768 (
            .O(N__10441),
            .I(N__10436));
    CascadeMux I__1767 (
            .O(N__10440),
            .I(N__10432));
    InMux I__1766 (
            .O(N__10439),
            .I(N__10429));
    InMux I__1765 (
            .O(N__10436),
            .I(N__10426));
    InMux I__1764 (
            .O(N__10435),
            .I(N__10421));
    InMux I__1763 (
            .O(N__10432),
            .I(N__10421));
    LocalMux I__1762 (
            .O(N__10429),
            .I(\uu2.N_90 ));
    LocalMux I__1761 (
            .O(N__10426),
            .I(\uu2.N_90 ));
    LocalMux I__1760 (
            .O(N__10421),
            .I(\uu2.N_90 ));
    SRMux I__1759 (
            .O(N__10414),
            .I(N__10409));
    IoInMux I__1758 (
            .O(N__10413),
            .I(N__10406));
    InMux I__1757 (
            .O(N__10412),
            .I(N__10403));
    LocalMux I__1756 (
            .O(N__10409),
            .I(N__10400));
    LocalMux I__1755 (
            .O(N__10406),
            .I(N__10397));
    LocalMux I__1754 (
            .O(N__10403),
            .I(N__10394));
    Span4Mux_v I__1753 (
            .O(N__10400),
            .I(N__10391));
    Span4Mux_s2_v I__1752 (
            .O(N__10397),
            .I(N__10388));
    Span4Mux_s2_v I__1751 (
            .O(N__10394),
            .I(N__10383));
    Span4Mux_s2_v I__1750 (
            .O(N__10391),
            .I(N__10383));
    Odrv4 I__1749 (
            .O(N__10388),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1748 (
            .O(N__10383),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1747 (
            .O(N__10378),
            .I(\buart.Z_rx.N_27_0_i_cascade_ ));
    CascadeMux I__1746 (
            .O(N__10375),
            .I(\buart.Z_rx.bitcount_lm_0_cascade_ ));
    CascadeMux I__1745 (
            .O(N__10372),
            .I(N__10369));
    InMux I__1744 (
            .O(N__10369),
            .I(N__10366));
    LocalMux I__1743 (
            .O(N__10366),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    CascadeMux I__1742 (
            .O(N__10363),
            .I(\buart.Z_rx.bitcount_lm_1_cascade_ ));
    CascadeMux I__1741 (
            .O(N__10360),
            .I(N__10352));
    InMux I__1740 (
            .O(N__10359),
            .I(N__10347));
    InMux I__1739 (
            .O(N__10358),
            .I(N__10347));
    InMux I__1738 (
            .O(N__10357),
            .I(N__10344));
    InMux I__1737 (
            .O(N__10356),
            .I(N__10339));
    InMux I__1736 (
            .O(N__10355),
            .I(N__10339));
    InMux I__1735 (
            .O(N__10352),
            .I(N__10336));
    LocalMux I__1734 (
            .O(N__10347),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1733 (
            .O(N__10344),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1732 (
            .O(N__10339),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1731 (
            .O(N__10336),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    CascadeMux I__1730 (
            .O(N__10327),
            .I(N__10324));
    InMux I__1729 (
            .O(N__10324),
            .I(N__10321));
    LocalMux I__1728 (
            .O(N__10321),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    CascadeMux I__1727 (
            .O(N__10318),
            .I(\Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_ ));
    InMux I__1726 (
            .O(N__10315),
            .I(N__10312));
    LocalMux I__1725 (
            .O(N__10312),
            .I(\uu2.bitmapZ0Z_75 ));
    InMux I__1724 (
            .O(N__10309),
            .I(N__10306));
    LocalMux I__1723 (
            .O(N__10306),
            .I(\Lab_UT.bcd2segment3.segment_i_0Z0Z_1 ));
    InMux I__1722 (
            .O(N__10303),
            .I(N__10300));
    LocalMux I__1721 (
            .O(N__10300),
            .I(\Lab_UT.bcd2segment3.segment_i_0Z0Z_2 ));
    InMux I__1720 (
            .O(N__10297),
            .I(N__10294));
    LocalMux I__1719 (
            .O(N__10294),
            .I(N__10291));
    Span4Mux_h I__1718 (
            .O(N__10291),
            .I(N__10288));
    Odrv4 I__1717 (
            .O(N__10288),
            .I(\resetGen.escKeyZ0Z_3 ));
    CascadeMux I__1716 (
            .O(N__10285),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_ ));
    CascadeMux I__1715 (
            .O(N__10282),
            .I(\uu2.N_4_cascade_ ));
    InMux I__1714 (
            .O(N__10279),
            .I(N__10276));
    LocalMux I__1713 (
            .O(N__10276),
            .I(N__10273));
    Odrv4 I__1712 (
            .O(N__10273),
            .I(\uu2.g0_17_1 ));
    InMux I__1711 (
            .O(N__10270),
            .I(N__10267));
    LocalMux I__1710 (
            .O(N__10267),
            .I(\uu2.bitmapZ0Z_72 ));
    InMux I__1709 (
            .O(N__10264),
            .I(N__10261));
    LocalMux I__1708 (
            .O(N__10261),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__1707 (
            .O(N__10258),
            .I(N__10255));
    LocalMux I__1706 (
            .O(N__10255),
            .I(\uu2.N_5 ));
    InMux I__1705 (
            .O(N__10252),
            .I(N__10249));
    LocalMux I__1704 (
            .O(N__10249),
            .I(\uu2.bitmapZ0Z_203 ));
    CascadeMux I__1703 (
            .O(N__10246),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_ ));
    InMux I__1702 (
            .O(N__10243),
            .I(N__10236));
    InMux I__1701 (
            .O(N__10242),
            .I(N__10233));
    InMux I__1700 (
            .O(N__10241),
            .I(N__10226));
    InMux I__1699 (
            .O(N__10240),
            .I(N__10226));
    InMux I__1698 (
            .O(N__10239),
            .I(N__10226));
    LocalMux I__1697 (
            .O(N__10236),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__1696 (
            .O(N__10233),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__1695 (
            .O(N__10226),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__1694 (
            .O(N__10219),
            .I(N__10216));
    LocalMux I__1693 (
            .O(N__10216),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__1692 (
            .O(N__10213),
            .I(N__10210));
    LocalMux I__1691 (
            .O(N__10210),
            .I(\uu2.bitmap_RNISSSNZ0Z_162 ));
    InMux I__1690 (
            .O(N__10207),
            .I(N__10204));
    LocalMux I__1689 (
            .O(N__10204),
            .I(\uu2.bitmapZ0Z_162 ));
    CascadeMux I__1688 (
            .O(N__10201),
            .I(\uu2.N_46_cascade_ ));
    InMux I__1687 (
            .O(N__10198),
            .I(N__10193));
    InMux I__1686 (
            .O(N__10197),
            .I(N__10190));
    InMux I__1685 (
            .O(N__10196),
            .I(N__10187));
    LocalMux I__1684 (
            .O(N__10193),
            .I(N__10184));
    LocalMux I__1683 (
            .O(N__10190),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    LocalMux I__1682 (
            .O(N__10187),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    Odrv4 I__1681 (
            .O(N__10184),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    InMux I__1680 (
            .O(N__10177),
            .I(N__10171));
    InMux I__1679 (
            .O(N__10176),
            .I(N__10171));
    LocalMux I__1678 (
            .O(N__10171),
            .I(N__10168));
    Span4Mux_h I__1677 (
            .O(N__10168),
            .I(N__10165));
    Odrv4 I__1676 (
            .O(N__10165),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    CascadeMux I__1675 (
            .O(N__10162),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_ ));
    CascadeMux I__1674 (
            .O(N__10159),
            .I(N__10156));
    InMux I__1673 (
            .O(N__10156),
            .I(N__10153));
    LocalMux I__1672 (
            .O(N__10153),
            .I(N__10150));
    Span4Mux_v I__1671 (
            .O(N__10150),
            .I(N__10147));
    Odrv4 I__1670 (
            .O(N__10147),
            .I(\uu2.un426_ci ));
    InMux I__1669 (
            .O(N__10144),
            .I(N__10138));
    InMux I__1668 (
            .O(N__10143),
            .I(N__10133));
    InMux I__1667 (
            .O(N__10142),
            .I(N__10133));
    InMux I__1666 (
            .O(N__10141),
            .I(N__10130));
    LocalMux I__1665 (
            .O(N__10138),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__1664 (
            .O(N__10133),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    LocalMux I__1663 (
            .O(N__10130),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    InMux I__1662 (
            .O(N__10123),
            .I(N__10120));
    LocalMux I__1661 (
            .O(N__10120),
            .I(N__10117));
    Span4Mux_h I__1660 (
            .O(N__10117),
            .I(N__10114));
    Odrv4 I__1659 (
            .O(N__10114),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_2 ));
    InMux I__1658 (
            .O(N__10111),
            .I(N__10108));
    LocalMux I__1657 (
            .O(N__10108),
            .I(N__10105));
    Odrv4 I__1656 (
            .O(N__10105),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__1655 (
            .O(N__10102),
            .I(\uu2.mem0.g0_7_3_cascade_ ));
    InMux I__1654 (
            .O(N__10099),
            .I(N__10096));
    LocalMux I__1653 (
            .O(N__10096),
            .I(\uu2.bitmap_pmux_27_ns_1_0 ));
    InMux I__1652 (
            .O(N__10093),
            .I(N__10090));
    LocalMux I__1651 (
            .O(N__10090),
            .I(\uu2.mem0.g0_6_4 ));
    CascadeMux I__1650 (
            .O(N__10087),
            .I(\uu2.mem0.g0_6_5_cascade_ ));
    CascadeMux I__1649 (
            .O(N__10084),
            .I(\uu2.N_150_cascade_ ));
    CascadeMux I__1648 (
            .O(N__10081),
            .I(N__10078));
    InMux I__1647 (
            .O(N__10078),
            .I(N__10073));
    InMux I__1646 (
            .O(N__10077),
            .I(N__10070));
    InMux I__1645 (
            .O(N__10076),
            .I(N__10067));
    LocalMux I__1644 (
            .O(N__10073),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__1643 (
            .O(N__10070),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__1642 (
            .O(N__10067),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CascadeMux I__1641 (
            .O(N__10060),
            .I(N__10057));
    InMux I__1640 (
            .O(N__10057),
            .I(N__10054));
    LocalMux I__1639 (
            .O(N__10054),
            .I(N__10051));
    Odrv4 I__1638 (
            .O(N__10051),
            .I(\uu2.mem0.N_78_i_0 ));
    InMux I__1637 (
            .O(N__10048),
            .I(N__10044));
    CascadeMux I__1636 (
            .O(N__10047),
            .I(N__10041));
    LocalMux I__1635 (
            .O(N__10044),
            .I(N__10038));
    InMux I__1634 (
            .O(N__10041),
            .I(N__10035));
    Span4Mux_v I__1633 (
            .O(N__10038),
            .I(N__10032));
    LocalMux I__1632 (
            .O(N__10035),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__1631 (
            .O(N__10032),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    CascadeMux I__1630 (
            .O(N__10027),
            .I(N__10024));
    InMux I__1629 (
            .O(N__10024),
            .I(N__10019));
    InMux I__1628 (
            .O(N__10023),
            .I(N__10014));
    InMux I__1627 (
            .O(N__10022),
            .I(N__10014));
    LocalMux I__1626 (
            .O(N__10019),
            .I(\uu2.N_93 ));
    LocalMux I__1625 (
            .O(N__10014),
            .I(\uu2.N_93 ));
    InMux I__1624 (
            .O(N__10009),
            .I(N__10003));
    InMux I__1623 (
            .O(N__10008),
            .I(N__10000));
    InMux I__1622 (
            .O(N__10007),
            .I(N__9997));
    InMux I__1621 (
            .O(N__10006),
            .I(N__9994));
    LocalMux I__1620 (
            .O(N__10003),
            .I(N__9991));
    LocalMux I__1619 (
            .O(N__10000),
            .I(N__9988));
    LocalMux I__1618 (
            .O(N__9997),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1617 (
            .O(N__9994),
            .I(\uu2.w_addr_userZ0Z_7 ));
    Odrv4 I__1616 (
            .O(N__9991),
            .I(\uu2.w_addr_userZ0Z_7 ));
    Odrv4 I__1615 (
            .O(N__9988),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__1614 (
            .O(N__9979),
            .I(N__9976));
    LocalMux I__1613 (
            .O(N__9976),
            .I(N__9973));
    Span12Mux_s7_v I__1612 (
            .O(N__9973),
            .I(N__9969));
    InMux I__1611 (
            .O(N__9972),
            .I(N__9966));
    Odrv12 I__1610 (
            .O(N__9969),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    LocalMux I__1609 (
            .O(N__9966),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__1608 (
            .O(N__9961),
            .I(N__9957));
    InMux I__1607 (
            .O(N__9960),
            .I(N__9954));
    LocalMux I__1606 (
            .O(N__9957),
            .I(N__9951));
    LocalMux I__1605 (
            .O(N__9954),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__1604 (
            .O(N__9951),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1603 (
            .O(N__9946),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__1602 (
            .O(N__9943),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1601 (
            .O(N__9940),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1600 (
            .O(N__9937),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    InMux I__1599 (
            .O(N__9934),
            .I(N__9931));
    LocalMux I__1598 (
            .O(N__9931),
            .I(\uu2.bitmapZ0Z_111 ));
    CascadeMux I__1597 (
            .O(N__9928),
            .I(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ));
    InMux I__1596 (
            .O(N__9925),
            .I(N__9922));
    LocalMux I__1595 (
            .O(N__9922),
            .I(N__9919));
    Odrv4 I__1594 (
            .O(N__9919),
            .I(\uu2.bitmap_pmux_sn_N_15 ));
    CascadeMux I__1593 (
            .O(N__9916),
            .I(\uu2.N_395_cascade_ ));
    InMux I__1592 (
            .O(N__9913),
            .I(N__9910));
    LocalMux I__1591 (
            .O(N__9910),
            .I(\uu2.N_56 ));
    InMux I__1590 (
            .O(N__9907),
            .I(N__9904));
    LocalMux I__1589 (
            .O(N__9904),
            .I(N__9900));
    InMux I__1588 (
            .O(N__9903),
            .I(N__9897));
    Span4Mux_h I__1587 (
            .O(N__9900),
            .I(N__9894));
    LocalMux I__1586 (
            .O(N__9897),
            .I(N__9891));
    Odrv4 I__1585 (
            .O(N__9894),
            .I(\uu2.N_401 ));
    Odrv12 I__1584 (
            .O(N__9891),
            .I(\uu2.N_401 ));
    CascadeMux I__1583 (
            .O(N__9886),
            .I(\buart.Z_rx.idle_1_cascade_ ));
    CascadeMux I__1582 (
            .O(N__9883),
            .I(\buart.Z_rx.valid_1_cascade_ ));
    CascadeMux I__1581 (
            .O(N__9880),
            .I(N__9875));
    CascadeMux I__1580 (
            .O(N__9879),
            .I(N__9872));
    CascadeMux I__1579 (
            .O(N__9878),
            .I(N__9869));
    InMux I__1578 (
            .O(N__9875),
            .I(N__9864));
    InMux I__1577 (
            .O(N__9872),
            .I(N__9864));
    InMux I__1576 (
            .O(N__9869),
            .I(N__9861));
    LocalMux I__1575 (
            .O(N__9864),
            .I(\uu2.bitmapZ0Z_314 ));
    LocalMux I__1574 (
            .O(N__9861),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__1573 (
            .O(N__9856),
            .I(N__9850));
    InMux I__1572 (
            .O(N__9855),
            .I(N__9850));
    LocalMux I__1571 (
            .O(N__9850),
            .I(\uu2.N_383 ));
    InMux I__1570 (
            .O(N__9847),
            .I(N__9844));
    LocalMux I__1569 (
            .O(N__9844),
            .I(\uu2.bitmapZ0Z_180 ));
    CascadeMux I__1568 (
            .O(N__9841),
            .I(\Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ));
    CascadeMux I__1567 (
            .O(N__9838),
            .I(\Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_ ));
    InMux I__1566 (
            .O(N__9835),
            .I(N__9832));
    LocalMux I__1565 (
            .O(N__9832),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__1564 (
            .O(N__9829),
            .I(N__9826));
    LocalMux I__1563 (
            .O(N__9826),
            .I(\uu2.bitmapZ0Z_40 ));
    InMux I__1562 (
            .O(N__9823),
            .I(N__9820));
    LocalMux I__1561 (
            .O(N__9820),
            .I(\uu2.bitmap_pmux_15_i_m2_ns_1 ));
    InMux I__1560 (
            .O(N__9817),
            .I(N__9814));
    LocalMux I__1559 (
            .O(N__9814),
            .I(\uu2.mem0.g1_3_0 ));
    InMux I__1558 (
            .O(N__9811),
            .I(N__9805));
    InMux I__1557 (
            .O(N__9810),
            .I(N__9805));
    LocalMux I__1556 (
            .O(N__9805),
            .I(N__9802));
    Odrv4 I__1555 (
            .O(N__9802),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__1554 (
            .O(N__9799),
            .I(N__9793));
    InMux I__1553 (
            .O(N__9798),
            .I(N__9793));
    LocalMux I__1552 (
            .O(N__9793),
            .I(N__9790));
    Odrv4 I__1551 (
            .O(N__9790),
            .I(\uu2.bitmapZ0Z_308 ));
    CascadeMux I__1550 (
            .O(N__9787),
            .I(\uu2.N_247_cascade_ ));
    CascadeMux I__1549 (
            .O(N__9784),
            .I(N__9781));
    InMux I__1548 (
            .O(N__9781),
            .I(N__9775));
    InMux I__1547 (
            .O(N__9780),
            .I(N__9775));
    LocalMux I__1546 (
            .O(N__9775),
            .I(\uu2.N_2171_0 ));
    InMux I__1545 (
            .O(N__9772),
            .I(N__9769));
    LocalMux I__1544 (
            .O(N__9769),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_44 ));
    CascadeMux I__1543 (
            .O(N__9766),
            .I(\Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_ ));
    CascadeMux I__1542 (
            .O(N__9763),
            .I(\Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_ ));
    InMux I__1541 (
            .O(N__9760),
            .I(N__9757));
    LocalMux I__1540 (
            .O(N__9757),
            .I(\uu2.bitmapZ0Z_34 ));
    CascadeMux I__1539 (
            .O(N__9754),
            .I(N__9751));
    InMux I__1538 (
            .O(N__9751),
            .I(N__9748));
    LocalMux I__1537 (
            .O(N__9748),
            .I(\uu2.bitmapZ0Z_290 ));
    CascadeMux I__1536 (
            .O(N__9745),
            .I(\uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_ ));
    CascadeMux I__1535 (
            .O(N__9742),
            .I(N__9738));
    InMux I__1534 (
            .O(N__9741),
            .I(N__9735));
    InMux I__1533 (
            .O(N__9738),
            .I(N__9732));
    LocalMux I__1532 (
            .O(N__9735),
            .I(\uu2.g2_0_0 ));
    LocalMux I__1531 (
            .O(N__9732),
            .I(\uu2.g2_0_0 ));
    CascadeMux I__1530 (
            .O(N__9727),
            .I(\uu2.mem0.g1_6_cascade_ ));
    InMux I__1529 (
            .O(N__9724),
            .I(N__9721));
    LocalMux I__1528 (
            .O(N__9721),
            .I(\uu2.mem0.N_1201_0_0_0 ));
    InMux I__1527 (
            .O(N__9718),
            .I(N__9715));
    LocalMux I__1526 (
            .O(N__9715),
            .I(\uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0 ));
    InMux I__1525 (
            .O(N__9712),
            .I(N__9706));
    InMux I__1524 (
            .O(N__9711),
            .I(N__9706));
    LocalMux I__1523 (
            .O(N__9706),
            .I(\uu2.bitmap_pmux_sn_N_20_0 ));
    InMux I__1522 (
            .O(N__9703),
            .I(N__9700));
    LocalMux I__1521 (
            .O(N__9700),
            .I(N__9697));
    Odrv4 I__1520 (
            .O(N__9697),
            .I(\uu2.bitmap_pmux_19_i_m2_ns_1 ));
    InMux I__1519 (
            .O(N__9694),
            .I(N__9691));
    LocalMux I__1518 (
            .O(N__9691),
            .I(\uu2.N_55_0 ));
    InMux I__1517 (
            .O(N__9688),
            .I(N__9685));
    LocalMux I__1516 (
            .O(N__9685),
            .I(\uu2.mem0.bitmap_pmux_sn_N_20_1_0_1 ));
    InMux I__1515 (
            .O(N__9682),
            .I(N__9679));
    LocalMux I__1514 (
            .O(N__9679),
            .I(\uu2.mem0.N_2166_1_0_1 ));
    CascadeMux I__1513 (
            .O(N__9676),
            .I(\uu2.mem0.N_247_0_cascade_ ));
    CascadeMux I__1512 (
            .O(N__9673),
            .I(\uu2.mem0.N_2171_1_0_1_cascade_ ));
    CascadeMux I__1511 (
            .O(N__9670),
            .I(N__9667));
    InMux I__1510 (
            .O(N__9667),
            .I(N__9661));
    InMux I__1509 (
            .O(N__9666),
            .I(N__9661));
    LocalMux I__1508 (
            .O(N__9661),
            .I(N__9657));
    InMux I__1507 (
            .O(N__9660),
            .I(N__9654));
    Odrv4 I__1506 (
            .O(N__9657),
            .I(\uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7 ));
    LocalMux I__1505 (
            .O(N__9654),
            .I(\uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7 ));
    InMux I__1504 (
            .O(N__9649),
            .I(N__9646));
    LocalMux I__1503 (
            .O(N__9646),
            .I(\uu2.mem0.N_397_1_0_1 ));
    CascadeMux I__1502 (
            .O(N__9643),
            .I(\uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_ ));
    InMux I__1501 (
            .O(N__9640),
            .I(N__9637));
    LocalMux I__1500 (
            .O(N__9637),
            .I(\uu2.mem0.g1_2_0 ));
    InMux I__1499 (
            .O(N__9634),
            .I(N__9631));
    LocalMux I__1498 (
            .O(N__9631),
            .I(\uu2.N_40_0 ));
    CascadeMux I__1497 (
            .O(N__9628),
            .I(N__9625));
    InMux I__1496 (
            .O(N__9625),
            .I(N__9622));
    LocalMux I__1495 (
            .O(N__9622),
            .I(\uu2.N_48_i_0 ));
    InMux I__1494 (
            .O(N__9619),
            .I(N__9616));
    LocalMux I__1493 (
            .O(N__9616),
            .I(\uu2.N_404 ));
    InMux I__1492 (
            .O(N__9613),
            .I(N__9610));
    LocalMux I__1491 (
            .O(N__9610),
            .I(\uu2.mem0.g1_1_1_0 ));
    CascadeMux I__1490 (
            .O(N__9607),
            .I(\uu2.N_404_cascade_ ));
    InMux I__1489 (
            .O(N__9604),
            .I(N__9601));
    LocalMux I__1488 (
            .O(N__9601),
            .I(\uu2.mem0.bitmap_pmux_1_0_0 ));
    CascadeMux I__1487 (
            .O(N__9598),
            .I(\uu2.mem0.bitmap_pmux_sn_N_42_cascade_ ));
    InMux I__1486 (
            .O(N__9595),
            .I(N__9592));
    LocalMux I__1485 (
            .O(N__9592),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_46 ));
    CascadeMux I__1484 (
            .O(N__9589),
            .I(\uu2.bitmap_pmux_20_ns_1_cascade_ ));
    CascadeMux I__1483 (
            .O(N__9586),
            .I(N__9583));
    InMux I__1482 (
            .O(N__9583),
            .I(N__9580));
    LocalMux I__1481 (
            .O(N__9580),
            .I(\Lab_UT.bcd2segment4.segment_0Z0Z_2 ));
    InMux I__1480 (
            .O(N__9577),
            .I(N__9574));
    LocalMux I__1479 (
            .O(N__9574),
            .I(\uu2.bitmapZ0Z_197 ));
    CascadeMux I__1478 (
            .O(N__9571),
            .I(\Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_ ));
    InMux I__1477 (
            .O(N__9568),
            .I(N__9565));
    LocalMux I__1476 (
            .O(N__9565),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__1475 (
            .O(N__9562),
            .I(N__9559));
    LocalMux I__1474 (
            .O(N__9559),
            .I(\Lab_UT.bcd2segment4.N_217 ));
    CascadeMux I__1473 (
            .O(N__9556),
            .I(N__9553));
    InMux I__1472 (
            .O(N__9553),
            .I(N__9550));
    LocalMux I__1471 (
            .O(N__9550),
            .I(\uu2.bitmapZ0Z_194 ));
    InMux I__1470 (
            .O(N__9547),
            .I(N__9544));
    LocalMux I__1469 (
            .O(N__9544),
            .I(\Lab_UT.bcd2segment4.segment_i_1Z0Z_5 ));
    InMux I__1468 (
            .O(N__9541),
            .I(N__9538));
    LocalMux I__1467 (
            .O(N__9538),
            .I(\uu2.bitmapZ0Z_66 ));
    CascadeMux I__1466 (
            .O(N__9535),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1465 (
            .O(N__9532),
            .I(N__9529));
    InMux I__1464 (
            .O(N__9529),
            .I(N__9526));
    LocalMux I__1463 (
            .O(N__9526),
            .I(N__9523));
    Span4Mux_h I__1462 (
            .O(N__9523),
            .I(N__9516));
    InMux I__1461 (
            .O(N__9522),
            .I(N__9511));
    InMux I__1460 (
            .O(N__9521),
            .I(N__9511));
    InMux I__1459 (
            .O(N__9520),
            .I(N__9506));
    InMux I__1458 (
            .O(N__9519),
            .I(N__9506));
    Odrv4 I__1457 (
            .O(N__9516),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1456 (
            .O(N__9511),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1455 (
            .O(N__9506),
            .I(\uu2.r_addrZ0Z_4 ));
    CascadeMux I__1454 (
            .O(N__9499),
            .I(N__9496));
    InMux I__1453 (
            .O(N__9496),
            .I(N__9493));
    LocalMux I__1452 (
            .O(N__9493),
            .I(N__9490));
    Span4Mux_s3_h I__1451 (
            .O(N__9490),
            .I(N__9484));
    InMux I__1450 (
            .O(N__9489),
            .I(N__9481));
    InMux I__1449 (
            .O(N__9488),
            .I(N__9478));
    InMux I__1448 (
            .O(N__9487),
            .I(N__9475));
    Odrv4 I__1447 (
            .O(N__9484),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1446 (
            .O(N__9481),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1445 (
            .O(N__9478),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__1444 (
            .O(N__9475),
            .I(\uu2.r_addrZ0Z_5 ));
    CEMux I__1443 (
            .O(N__9466),
            .I(N__9463));
    LocalMux I__1442 (
            .O(N__9463),
            .I(N__9460));
    Odrv4 I__1441 (
            .O(N__9460),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__1440 (
            .O(N__9457),
            .I(N__9454));
    InMux I__1439 (
            .O(N__9454),
            .I(N__9451));
    LocalMux I__1438 (
            .O(N__9451),
            .I(N__9448));
    Span4Mux_s3_h I__1437 (
            .O(N__9448),
            .I(N__9445));
    Odrv4 I__1436 (
            .O(N__9445),
            .I(\uu2.mem0.N_70_i ));
    CascadeMux I__1435 (
            .O(N__9442),
            .I(N__9439));
    InMux I__1434 (
            .O(N__9439),
            .I(N__9436));
    LocalMux I__1433 (
            .O(N__9436),
            .I(N__9431));
    InMux I__1432 (
            .O(N__9435),
            .I(N__9425));
    InMux I__1431 (
            .O(N__9434),
            .I(N__9425));
    Span4Mux_h I__1430 (
            .O(N__9431),
            .I(N__9422));
    InMux I__1429 (
            .O(N__9430),
            .I(N__9419));
    LocalMux I__1428 (
            .O(N__9425),
            .I(\uu2.r_addrZ0Z_6 ));
    Odrv4 I__1427 (
            .O(N__9422),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1426 (
            .O(N__9419),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1425 (
            .O(N__9412),
            .I(N__9409));
    InMux I__1424 (
            .O(N__9409),
            .I(N__9406));
    LocalMux I__1423 (
            .O(N__9406),
            .I(N__9401));
    InMux I__1422 (
            .O(N__9405),
            .I(N__9398));
    InMux I__1421 (
            .O(N__9404),
            .I(N__9395));
    Span4Mux_v I__1420 (
            .O(N__9401),
            .I(N__9392));
    LocalMux I__1419 (
            .O(N__9398),
            .I(N__9387));
    LocalMux I__1418 (
            .O(N__9395),
            .I(N__9387));
    Odrv4 I__1417 (
            .O(N__9392),
            .I(\uu2.r_addrZ0Z_7 ));
    Odrv4 I__1416 (
            .O(N__9387),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__1415 (
            .O(N__9382),
            .I(N__9379));
    LocalMux I__1414 (
            .O(N__9379),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    InMux I__1413 (
            .O(N__9376),
            .I(N__9372));
    CascadeMux I__1412 (
            .O(N__9375),
            .I(N__9367));
    LocalMux I__1411 (
            .O(N__9372),
            .I(N__9364));
    InMux I__1410 (
            .O(N__9371),
            .I(N__9361));
    InMux I__1409 (
            .O(N__9370),
            .I(N__9358));
    InMux I__1408 (
            .O(N__9367),
            .I(N__9355));
    Span4Mux_h I__1407 (
            .O(N__9364),
            .I(N__9352));
    LocalMux I__1406 (
            .O(N__9361),
            .I(N__9347));
    LocalMux I__1405 (
            .O(N__9358),
            .I(N__9347));
    LocalMux I__1404 (
            .O(N__9355),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__1403 (
            .O(N__9352),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv12 I__1402 (
            .O(N__9347),
            .I(\uu2.r_addrZ0Z_2 ));
    InMux I__1401 (
            .O(N__9340),
            .I(N__9336));
    CascadeMux I__1400 (
            .O(N__9339),
            .I(N__9332));
    LocalMux I__1399 (
            .O(N__9336),
            .I(N__9329));
    InMux I__1398 (
            .O(N__9335),
            .I(N__9324));
    InMux I__1397 (
            .O(N__9332),
            .I(N__9321));
    Span4Mux_h I__1396 (
            .O(N__9329),
            .I(N__9318));
    InMux I__1395 (
            .O(N__9328),
            .I(N__9313));
    InMux I__1394 (
            .O(N__9327),
            .I(N__9313));
    LocalMux I__1393 (
            .O(N__9324),
            .I(N__9310));
    LocalMux I__1392 (
            .O(N__9321),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv4 I__1391 (
            .O(N__9318),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1390 (
            .O(N__9313),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv12 I__1389 (
            .O(N__9310),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1388 (
            .O(N__9301),
            .I(N__9298));
    InMux I__1387 (
            .O(N__9298),
            .I(N__9295));
    LocalMux I__1386 (
            .O(N__9295),
            .I(N__9290));
    CascadeMux I__1385 (
            .O(N__9294),
            .I(N__9287));
    CascadeMux I__1384 (
            .O(N__9293),
            .I(N__9284));
    Span4Mux_h I__1383 (
            .O(N__9290),
            .I(N__9281));
    InMux I__1382 (
            .O(N__9287),
            .I(N__9278));
    InMux I__1381 (
            .O(N__9284),
            .I(N__9275));
    Odrv4 I__1380 (
            .O(N__9281),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1379 (
            .O(N__9278),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1378 (
            .O(N__9275),
            .I(\uu2.r_addrZ0Z_3 ));
    InMux I__1377 (
            .O(N__9268),
            .I(N__9264));
    CascadeMux I__1376 (
            .O(N__9267),
            .I(N__9260));
    LocalMux I__1375 (
            .O(N__9264),
            .I(N__9257));
    InMux I__1374 (
            .O(N__9263),
            .I(N__9251));
    InMux I__1373 (
            .O(N__9260),
            .I(N__9248));
    Span4Mux_h I__1372 (
            .O(N__9257),
            .I(N__9245));
    InMux I__1371 (
            .O(N__9256),
            .I(N__9238));
    InMux I__1370 (
            .O(N__9255),
            .I(N__9238));
    InMux I__1369 (
            .O(N__9254),
            .I(N__9238));
    LocalMux I__1368 (
            .O(N__9251),
            .I(N__9235));
    LocalMux I__1367 (
            .O(N__9248),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__1366 (
            .O(N__9245),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1365 (
            .O(N__9238),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv12 I__1364 (
            .O(N__9235),
            .I(\uu2.r_addrZ0Z_0 ));
    CascadeMux I__1363 (
            .O(N__9226),
            .I(N__9223));
    InMux I__1362 (
            .O(N__9223),
            .I(N__9216));
    InMux I__1361 (
            .O(N__9222),
            .I(N__9211));
    InMux I__1360 (
            .O(N__9221),
            .I(N__9211));
    InMux I__1359 (
            .O(N__9220),
            .I(N__9206));
    InMux I__1358 (
            .O(N__9219),
            .I(N__9206));
    LocalMux I__1357 (
            .O(N__9216),
            .I(\uu2.un404_ci ));
    LocalMux I__1356 (
            .O(N__9211),
            .I(\uu2.un404_ci ));
    LocalMux I__1355 (
            .O(N__9206),
            .I(\uu2.un404_ci ));
    InMux I__1354 (
            .O(N__9199),
            .I(N__9196));
    LocalMux I__1353 (
            .O(N__9196),
            .I(N__9190));
    InMux I__1352 (
            .O(N__9195),
            .I(N__9187));
    InMux I__1351 (
            .O(N__9194),
            .I(N__9182));
    InMux I__1350 (
            .O(N__9193),
            .I(N__9182));
    Span4Mux_h I__1349 (
            .O(N__9190),
            .I(N__9179));
    LocalMux I__1348 (
            .O(N__9187),
            .I(o_One_Sec_Pulse));
    LocalMux I__1347 (
            .O(N__9182),
            .I(o_One_Sec_Pulse));
    Odrv4 I__1346 (
            .O(N__9179),
            .I(o_One_Sec_Pulse));
    InMux I__1345 (
            .O(N__9172),
            .I(N__9169));
    LocalMux I__1344 (
            .O(N__9169),
            .I(N__9165));
    InMux I__1343 (
            .O(N__9168),
            .I(N__9162));
    Span4Mux_s3_h I__1342 (
            .O(N__9165),
            .I(N__9159));
    LocalMux I__1341 (
            .O(N__9162),
            .I(N__9154));
    Span4Mux_v I__1340 (
            .O(N__9159),
            .I(N__9151));
    InMux I__1339 (
            .O(N__9158),
            .I(N__9146));
    InMux I__1338 (
            .O(N__9157),
            .I(N__9146));
    Span4Mux_v I__1337 (
            .O(N__9154),
            .I(N__9143));
    Odrv4 I__1336 (
            .O(N__9151),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__1335 (
            .O(N__9146),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__1334 (
            .O(N__9143),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__1333 (
            .O(N__9136),
            .I(N__9133));
    LocalMux I__1332 (
            .O(N__9133),
            .I(N__9129));
    InMux I__1331 (
            .O(N__9132),
            .I(N__9126));
    Span4Mux_s3_h I__1330 (
            .O(N__9129),
            .I(N__9123));
    LocalMux I__1329 (
            .O(N__9126),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__1328 (
            .O(N__9123),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__1327 (
            .O(N__9118),
            .I(N__9115));
    LocalMux I__1326 (
            .O(N__9115),
            .I(N__9112));
    Span4Mux_v I__1325 (
            .O(N__9112),
            .I(N__9109));
    Odrv4 I__1324 (
            .O(N__9109),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    CascadeMux I__1323 (
            .O(N__9106),
            .I(N__9103));
    InMux I__1322 (
            .O(N__9103),
            .I(N__9092));
    InMux I__1321 (
            .O(N__9102),
            .I(N__9092));
    InMux I__1320 (
            .O(N__9101),
            .I(N__9092));
    InMux I__1319 (
            .O(N__9100),
            .I(N__9089));
    InMux I__1318 (
            .O(N__9099),
            .I(N__9086));
    LocalMux I__1317 (
            .O(N__9092),
            .I(N__9082));
    LocalMux I__1316 (
            .O(N__9089),
            .I(N__9079));
    LocalMux I__1315 (
            .O(N__9086),
            .I(N__9076));
    InMux I__1314 (
            .O(N__9085),
            .I(N__9073));
    Span4Mux_h I__1313 (
            .O(N__9082),
            .I(N__9070));
    Span4Mux_s3_h I__1312 (
            .O(N__9079),
            .I(N__9067));
    Span4Mux_s3_h I__1311 (
            .O(N__9076),
            .I(N__9064));
    LocalMux I__1310 (
            .O(N__9073),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__1309 (
            .O(N__9070),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__1308 (
            .O(N__9067),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__1307 (
            .O(N__9064),
            .I(\uu0.l_precountZ0Z_0 ));
    InMux I__1306 (
            .O(N__9055),
            .I(N__9052));
    LocalMux I__1305 (
            .O(N__9052),
            .I(N__9049));
    IoSpan4Mux I__1304 (
            .O(N__9049),
            .I(N__9046));
    IoSpan4Mux I__1303 (
            .O(N__9046),
            .I(N__9043));
    IoSpan4Mux I__1302 (
            .O(N__9043),
            .I(N__9040));
    Odrv4 I__1301 (
            .O(N__9040),
            .I(uart_RXD));
    CascadeMux I__1300 (
            .O(N__9037),
            .I(N__9034));
    InMux I__1299 (
            .O(N__9034),
            .I(N__9031));
    LocalMux I__1298 (
            .O(N__9031),
            .I(N__9028));
    Span4Mux_h I__1297 (
            .O(N__9028),
            .I(N__9024));
    InMux I__1296 (
            .O(N__9027),
            .I(N__9021));
    Odrv4 I__1295 (
            .O(N__9024),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1294 (
            .O(N__9021),
            .I(\uu2.r_addrZ0Z_8 ));
    CascadeMux I__1293 (
            .O(N__9016),
            .I(N__9013));
    InMux I__1292 (
            .O(N__9013),
            .I(N__9010));
    LocalMux I__1291 (
            .O(N__9010),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    InMux I__1290 (
            .O(N__9007),
            .I(N__9004));
    LocalMux I__1289 (
            .O(N__9004),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__1288 (
            .O(N__9001),
            .I(N__8998));
    LocalMux I__1287 (
            .O(N__8998),
            .I(\uu2.bitmap_RNI8LB51Z0Z_186 ));
    CascadeMux I__1286 (
            .O(N__8995),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ));
    CascadeMux I__1285 (
            .O(N__8992),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ));
    CascadeMux I__1284 (
            .O(N__8989),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_ ));
    InMux I__1283 (
            .O(N__8986),
            .I(N__8983));
    LocalMux I__1282 (
            .O(N__8983),
            .I(\uu2.bitmapZ0Z_90 ));
    CascadeMux I__1281 (
            .O(N__8980),
            .I(N__8977));
    InMux I__1280 (
            .O(N__8977),
            .I(N__8974));
    LocalMux I__1279 (
            .O(N__8974),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__1278 (
            .O(N__8971),
            .I(N__8968));
    LocalMux I__1277 (
            .O(N__8968),
            .I(\uu2.mem0.bitmap_pmux_sn_i7_mux_0 ));
    InMux I__1276 (
            .O(N__8965),
            .I(N__8962));
    LocalMux I__1275 (
            .O(N__8962),
            .I(N__8959));
    Odrv4 I__1274 (
            .O(N__8959),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ));
    CascadeMux I__1273 (
            .O(N__8956),
            .I(\Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_ ));
    CascadeMux I__1272 (
            .O(N__8953),
            .I(\uu2.bitmap_RNIMQ601Z0Z_58_cascade_ ));
    CascadeMux I__1271 (
            .O(N__8950),
            .I(\Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_ ));
    InMux I__1270 (
            .O(N__8947),
            .I(N__8944));
    LocalMux I__1269 (
            .O(N__8944),
            .I(\uu2.bitmapZ0Z_58 ));
    CascadeMux I__1268 (
            .O(N__8941),
            .I(N__8938));
    InMux I__1267 (
            .O(N__8938),
            .I(N__8935));
    LocalMux I__1266 (
            .O(N__8935),
            .I(\uu2.mem0.N_71_i ));
    InMux I__1265 (
            .O(N__8932),
            .I(N__8929));
    LocalMux I__1264 (
            .O(N__8929),
            .I(\uu2.mem0.w_data_1 ));
    CascadeMux I__1263 (
            .O(N__8926),
            .I(N__8923));
    InMux I__1262 (
            .O(N__8923),
            .I(N__8920));
    LocalMux I__1261 (
            .O(N__8920),
            .I(N__8917));
    Odrv4 I__1260 (
            .O(N__8917),
            .I(\uu2.mem0.N_76_i_0 ));
    CascadeMux I__1259 (
            .O(N__8914),
            .I(\uu2.mem0.N_2166_0_cascade_ ));
    CascadeMux I__1258 (
            .O(N__8911),
            .I(\uu2.mem0.bitmap_pmux_0_cascade_ ));
    InMux I__1257 (
            .O(N__8908),
            .I(N__8905));
    LocalMux I__1256 (
            .O(N__8905),
            .I(N__8902));
    Span4Mux_s3_h I__1255 (
            .O(N__8902),
            .I(N__8899));
    Odrv4 I__1254 (
            .O(N__8899),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1253 (
            .O(N__8896),
            .I(N__8893));
    LocalMux I__1252 (
            .O(N__8893),
            .I(\uu2.mem0.ram512X8_inst_RNOZ0Z_42 ));
    CascadeMux I__1251 (
            .O(N__8890),
            .I(N__8887));
    InMux I__1250 (
            .O(N__8887),
            .I(N__8884));
    LocalMux I__1249 (
            .O(N__8884),
            .I(N__8881));
    Odrv4 I__1248 (
            .O(N__8881),
            .I(\uu2.mem0.N_75_i ));
    InMux I__1247 (
            .O(N__8878),
            .I(N__8875));
    LocalMux I__1246 (
            .O(N__8875),
            .I(\uu2.N_361 ));
    CascadeMux I__1245 (
            .O(N__8872),
            .I(\uu2.N_361_cascade_ ));
    InMux I__1244 (
            .O(N__8869),
            .I(N__8866));
    LocalMux I__1243 (
            .O(N__8866),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1242 (
            .O(N__8863),
            .I(N__8860));
    LocalMux I__1241 (
            .O(N__8860),
            .I(N__8857));
    Odrv4 I__1240 (
            .O(N__8857),
            .I(\uu2.mem0.N_69_i ));
    InMux I__1239 (
            .O(N__8854),
            .I(N__8851));
    LocalMux I__1238 (
            .O(N__8851),
            .I(\uu2.mem0.w_data_0_a3_0_4 ));
    CascadeMux I__1237 (
            .O(N__8848),
            .I(\uu2.N_61_cascade_ ));
    CascadeMux I__1236 (
            .O(N__8845),
            .I(\uu2.mem0.un51_w_data_displaying_cascade_ ));
    InMux I__1235 (
            .O(N__8842),
            .I(N__8839));
    LocalMux I__1234 (
            .O(N__8839),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1233 (
            .O(N__8836),
            .I(N__8833));
    LocalMux I__1232 (
            .O(N__8833),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__1231 (
            .O(N__8830),
            .I(N__8826));
    InMux I__1230 (
            .O(N__8829),
            .I(N__8823));
    LocalMux I__1229 (
            .O(N__8826),
            .I(N__8820));
    LocalMux I__1228 (
            .O(N__8823),
            .I(N__8817));
    Span4Mux_h I__1227 (
            .O(N__8820),
            .I(N__8814));
    Odrv12 I__1226 (
            .O(N__8817),
            .I(\uu2.un1_l_count_1_0 ));
    Odrv4 I__1225 (
            .O(N__8814),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1224 (
            .O(N__8809),
            .I(N__8806));
    LocalMux I__1223 (
            .O(N__8806),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1222 (
            .O(N__8803),
            .I(N__8797));
    InMux I__1221 (
            .O(N__8802),
            .I(N__8797));
    LocalMux I__1220 (
            .O(N__8797),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    CascadeMux I__1219 (
            .O(N__8794),
            .I(N__8791));
    InMux I__1218 (
            .O(N__8791),
            .I(N__8783));
    InMux I__1217 (
            .O(N__8790),
            .I(N__8783));
    InMux I__1216 (
            .O(N__8789),
            .I(N__8780));
    CascadeMux I__1215 (
            .O(N__8788),
            .I(N__8777));
    LocalMux I__1214 (
            .O(N__8783),
            .I(N__8771));
    LocalMux I__1213 (
            .O(N__8780),
            .I(N__8771));
    InMux I__1212 (
            .O(N__8777),
            .I(N__8766));
    InMux I__1211 (
            .O(N__8776),
            .I(N__8766));
    Span4Mux_v I__1210 (
            .O(N__8771),
            .I(N__8763));
    LocalMux I__1209 (
            .O(N__8766),
            .I(\uu2.trig_rd_is_det ));
    Odrv4 I__1208 (
            .O(N__8763),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__1207 (
            .O(N__8758),
            .I(\uu2.trig_rd_is_det_cascade_ ));
    InMux I__1206 (
            .O(N__8755),
            .I(N__8750));
    InMux I__1205 (
            .O(N__8754),
            .I(N__8745));
    InMux I__1204 (
            .O(N__8753),
            .I(N__8745));
    LocalMux I__1203 (
            .O(N__8750),
            .I(N__8742));
    LocalMux I__1202 (
            .O(N__8745),
            .I(N__8737));
    Span4Mux_v I__1201 (
            .O(N__8742),
            .I(N__8737));
    Odrv4 I__1200 (
            .O(N__8737),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__1199 (
            .O(N__8734),
            .I(N__8731));
    InMux I__1198 (
            .O(N__8731),
            .I(N__8728));
    LocalMux I__1197 (
            .O(N__8728),
            .I(\uu2.mem0.N_77_i ));
    CascadeMux I__1196 (
            .O(N__8725),
            .I(\uu2.mem0.w_data_i_a3_1_0_cascade_ ));
    InMux I__1195 (
            .O(N__8722),
            .I(N__8719));
    LocalMux I__1194 (
            .O(N__8719),
            .I(\uu2.mem0.N_79_i_0 ));
    CascadeMux I__1193 (
            .O(N__8716),
            .I(N__8713));
    InMux I__1192 (
            .O(N__8713),
            .I(N__8709));
    IoInMux I__1191 (
            .O(N__8712),
            .I(N__8706));
    LocalMux I__1190 (
            .O(N__8709),
            .I(N__8703));
    LocalMux I__1189 (
            .O(N__8706),
            .I(N__8700));
    Span4Mux_h I__1188 (
            .O(N__8703),
            .I(N__8697));
    Span12Mux_s9_v I__1187 (
            .O(N__8700),
            .I(N__8692));
    Sp12to4 I__1186 (
            .O(N__8697),
            .I(N__8692));
    Odrv12 I__1185 (
            .O(N__8692),
            .I(clk));
    SRMux I__1184 (
            .O(N__8689),
            .I(N__8686));
    LocalMux I__1183 (
            .O(N__8686),
            .I(N__8683));
    Span4Mux_s3_h I__1182 (
            .O(N__8683),
            .I(N__8680));
    Span4Mux_h I__1181 (
            .O(N__8680),
            .I(N__8676));
    CEMux I__1180 (
            .O(N__8679),
            .I(N__8673));
    Odrv4 I__1179 (
            .O(N__8676),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    LocalMux I__1178 (
            .O(N__8673),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1177 (
            .O(N__8668),
            .I(\uu0.un110_ci_cascade_ ));
    CascadeMux I__1176 (
            .O(N__8665),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__1175 (
            .O(N__8662),
            .I(N__8658));
    InMux I__1174 (
            .O(N__8661),
            .I(N__8655));
    LocalMux I__1173 (
            .O(N__8658),
            .I(N__8652));
    LocalMux I__1172 (
            .O(N__8655),
            .I(\uu0.l_countZ0Z_18 ));
    Odrv4 I__1171 (
            .O(N__8652),
            .I(\uu0.l_countZ0Z_18 ));
    CascadeMux I__1170 (
            .O(N__8647),
            .I(N__8644));
    InMux I__1169 (
            .O(N__8644),
            .I(N__8641));
    LocalMux I__1168 (
            .O(N__8641),
            .I(N__8638));
    Odrv4 I__1167 (
            .O(N__8638),
            .I(\uu0.un99_ci_0 ));
    InMux I__1166 (
            .O(N__8635),
            .I(N__8626));
    InMux I__1165 (
            .O(N__8634),
            .I(N__8626));
    InMux I__1164 (
            .O(N__8633),
            .I(N__8626));
    LocalMux I__1163 (
            .O(N__8626),
            .I(\uu0.l_countZ0Z_7 ));
    CascadeMux I__1162 (
            .O(N__8623),
            .I(N__8619));
    CascadeMux I__1161 (
            .O(N__8622),
            .I(N__8616));
    InMux I__1160 (
            .O(N__8619),
            .I(N__8613));
    InMux I__1159 (
            .O(N__8616),
            .I(N__8610));
    LocalMux I__1158 (
            .O(N__8613),
            .I(N__8607));
    LocalMux I__1157 (
            .O(N__8610),
            .I(N__8604));
    Odrv12 I__1156 (
            .O(N__8607),
            .I(\uu0.un88_ci_3 ));
    Odrv4 I__1155 (
            .O(N__8604),
            .I(\uu0.un88_ci_3 ));
    InMux I__1154 (
            .O(N__8599),
            .I(N__8585));
    InMux I__1153 (
            .O(N__8598),
            .I(N__8578));
    InMux I__1152 (
            .O(N__8597),
            .I(N__8578));
    InMux I__1151 (
            .O(N__8596),
            .I(N__8578));
    InMux I__1150 (
            .O(N__8595),
            .I(N__8569));
    InMux I__1149 (
            .O(N__8594),
            .I(N__8569));
    InMux I__1148 (
            .O(N__8593),
            .I(N__8569));
    InMux I__1147 (
            .O(N__8592),
            .I(N__8569));
    InMux I__1146 (
            .O(N__8591),
            .I(N__8566));
    InMux I__1145 (
            .O(N__8590),
            .I(N__8559));
    InMux I__1144 (
            .O(N__8589),
            .I(N__8559));
    InMux I__1143 (
            .O(N__8588),
            .I(N__8559));
    LocalMux I__1142 (
            .O(N__8585),
            .I(N__8556));
    LocalMux I__1141 (
            .O(N__8578),
            .I(N__8551));
    LocalMux I__1140 (
            .O(N__8569),
            .I(N__8551));
    LocalMux I__1139 (
            .O(N__8566),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1138 (
            .O(N__8559),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1137 (
            .O(N__8556),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1136 (
            .O(N__8551),
            .I(\uu0.un4_l_count_0 ));
    InMux I__1135 (
            .O(N__8542),
            .I(N__8536));
    InMux I__1134 (
            .O(N__8541),
            .I(N__8533));
    InMux I__1133 (
            .O(N__8540),
            .I(N__8528));
    InMux I__1132 (
            .O(N__8539),
            .I(N__8528));
    LocalMux I__1131 (
            .O(N__8536),
            .I(N__8523));
    LocalMux I__1130 (
            .O(N__8533),
            .I(N__8523));
    LocalMux I__1129 (
            .O(N__8528),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1128 (
            .O(N__8523),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__1127 (
            .O(N__8518),
            .I(N__8511));
    InMux I__1126 (
            .O(N__8517),
            .I(N__8508));
    InMux I__1125 (
            .O(N__8516),
            .I(N__8501));
    InMux I__1124 (
            .O(N__8515),
            .I(N__8501));
    InMux I__1123 (
            .O(N__8514),
            .I(N__8501));
    LocalMux I__1122 (
            .O(N__8511),
            .I(N__8494));
    LocalMux I__1121 (
            .O(N__8508),
            .I(N__8494));
    LocalMux I__1120 (
            .O(N__8501),
            .I(N__8494));
    Odrv4 I__1119 (
            .O(N__8494),
            .I(\uu0.un66_ci ));
    InMux I__1118 (
            .O(N__8491),
            .I(N__8488));
    LocalMux I__1117 (
            .O(N__8488),
            .I(N__8482));
    InMux I__1116 (
            .O(N__8487),
            .I(N__8479));
    InMux I__1115 (
            .O(N__8486),
            .I(N__8476));
    InMux I__1114 (
            .O(N__8485),
            .I(N__8473));
    Span4Mux_h I__1113 (
            .O(N__8482),
            .I(N__8470));
    LocalMux I__1112 (
            .O(N__8479),
            .I(N__8467));
    LocalMux I__1111 (
            .O(N__8476),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__1110 (
            .O(N__8473),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__1109 (
            .O(N__8470),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__1108 (
            .O(N__8467),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__1107 (
            .O(N__8458),
            .I(N__8453));
    InMux I__1106 (
            .O(N__8457),
            .I(N__8450));
    InMux I__1105 (
            .O(N__8456),
            .I(N__8447));
    LocalMux I__1104 (
            .O(N__8453),
            .I(N__8442));
    LocalMux I__1103 (
            .O(N__8450),
            .I(N__8442));
    LocalMux I__1102 (
            .O(N__8447),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv4 I__1101 (
            .O(N__8442),
            .I(\uu0.l_countZ0Z_5 ));
    InMux I__1100 (
            .O(N__8437),
            .I(N__8432));
    InMux I__1099 (
            .O(N__8436),
            .I(N__8427));
    InMux I__1098 (
            .O(N__8435),
            .I(N__8427));
    LocalMux I__1097 (
            .O(N__8432),
            .I(\uu0.un198_ci_2 ));
    LocalMux I__1096 (
            .O(N__8427),
            .I(\uu0.un198_ci_2 ));
    CascadeMux I__1095 (
            .O(N__8422),
            .I(N__8417));
    InMux I__1094 (
            .O(N__8421),
            .I(N__8413));
    InMux I__1093 (
            .O(N__8420),
            .I(N__8408));
    InMux I__1092 (
            .O(N__8417),
            .I(N__8408));
    CascadeMux I__1091 (
            .O(N__8416),
            .I(N__8401));
    LocalMux I__1090 (
            .O(N__8413),
            .I(N__8396));
    LocalMux I__1089 (
            .O(N__8408),
            .I(N__8396));
    CascadeMux I__1088 (
            .O(N__8407),
            .I(N__8393));
    CascadeMux I__1087 (
            .O(N__8406),
            .I(N__8390));
    CascadeMux I__1086 (
            .O(N__8405),
            .I(N__8387));
    CascadeMux I__1085 (
            .O(N__8404),
            .I(N__8384));
    InMux I__1084 (
            .O(N__8401),
            .I(N__8379));
    Span4Mux_s2_h I__1083 (
            .O(N__8396),
            .I(N__8376));
    InMux I__1082 (
            .O(N__8393),
            .I(N__8373));
    InMux I__1081 (
            .O(N__8390),
            .I(N__8370));
    InMux I__1080 (
            .O(N__8387),
            .I(N__8361));
    InMux I__1079 (
            .O(N__8384),
            .I(N__8361));
    InMux I__1078 (
            .O(N__8383),
            .I(N__8361));
    InMux I__1077 (
            .O(N__8382),
            .I(N__8361));
    LocalMux I__1076 (
            .O(N__8379),
            .I(N__8358));
    Odrv4 I__1075 (
            .O(N__8376),
            .I(\uu0.un110_ci ));
    LocalMux I__1074 (
            .O(N__8373),
            .I(\uu0.un110_ci ));
    LocalMux I__1073 (
            .O(N__8370),
            .I(\uu0.un110_ci ));
    LocalMux I__1072 (
            .O(N__8361),
            .I(\uu0.un110_ci ));
    Odrv4 I__1071 (
            .O(N__8358),
            .I(\uu0.un110_ci ));
    InMux I__1070 (
            .O(N__8347),
            .I(N__8344));
    LocalMux I__1069 (
            .O(N__8344),
            .I(N__8338));
    InMux I__1068 (
            .O(N__8343),
            .I(N__8333));
    InMux I__1067 (
            .O(N__8342),
            .I(N__8333));
    InMux I__1066 (
            .O(N__8341),
            .I(N__8330));
    Odrv4 I__1065 (
            .O(N__8338),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1064 (
            .O(N__8333),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1063 (
            .O(N__8330),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__1062 (
            .O(N__8323),
            .I(N__8319));
    InMux I__1061 (
            .O(N__8322),
            .I(N__8313));
    InMux I__1060 (
            .O(N__8319),
            .I(N__8313));
    InMux I__1059 (
            .O(N__8318),
            .I(N__8310));
    LocalMux I__1058 (
            .O(N__8313),
            .I(N__8307));
    LocalMux I__1057 (
            .O(N__8310),
            .I(\uu0.l_countZ0Z_17 ));
    Odrv4 I__1056 (
            .O(N__8307),
            .I(\uu0.l_countZ0Z_17 ));
    CEMux I__1055 (
            .O(N__8302),
            .I(N__8284));
    CEMux I__1054 (
            .O(N__8301),
            .I(N__8284));
    CEMux I__1053 (
            .O(N__8300),
            .I(N__8284));
    CEMux I__1052 (
            .O(N__8299),
            .I(N__8284));
    CEMux I__1051 (
            .O(N__8298),
            .I(N__8284));
    CEMux I__1050 (
            .O(N__8297),
            .I(N__8284));
    GlobalMux I__1049 (
            .O(N__8284),
            .I(N__8281));
    gio2CtrlBuf I__1048 (
            .O(N__8281),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__1047 (
            .O(N__8278),
            .I(\resetGen.escKeyZ0_cascade_ ));
    CascadeMux I__1046 (
            .O(N__8275),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__1045 (
            .O(N__8272),
            .I(N__8269));
    LocalMux I__1044 (
            .O(N__8269),
            .I(N__8265));
    InMux I__1043 (
            .O(N__8268),
            .I(N__8262));
    Odrv4 I__1042 (
            .O(N__8265),
            .I(\resetGen.reset_countZ0Z_3 ));
    LocalMux I__1041 (
            .O(N__8262),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__1040 (
            .O(N__8257),
            .I(N__8247));
    InMux I__1039 (
            .O(N__8256),
            .I(N__8247));
    InMux I__1038 (
            .O(N__8255),
            .I(N__8247));
    InMux I__1037 (
            .O(N__8254),
            .I(N__8244));
    LocalMux I__1036 (
            .O(N__8247),
            .I(\resetGen.reset_countZ0Z_0 ));
    LocalMux I__1035 (
            .O(N__8244),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__1034 (
            .O(N__8239),
            .I(N__8232));
    InMux I__1033 (
            .O(N__8238),
            .I(N__8232));
    InMux I__1032 (
            .O(N__8237),
            .I(N__8229));
    LocalMux I__1031 (
            .O(N__8232),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__1030 (
            .O(N__8229),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__1029 (
            .O(N__8224),
            .I(N__8221));
    InMux I__1028 (
            .O(N__8221),
            .I(N__8214));
    InMux I__1027 (
            .O(N__8220),
            .I(N__8214));
    InMux I__1026 (
            .O(N__8219),
            .I(N__8211));
    LocalMux I__1025 (
            .O(N__8214),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__1024 (
            .O(N__8211),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__1023 (
            .O(N__8206),
            .I(N__8200));
    InMux I__1022 (
            .O(N__8205),
            .I(N__8200));
    LocalMux I__1021 (
            .O(N__8200),
            .I(N__8197));
    Odrv12 I__1020 (
            .O(N__8197),
            .I(\resetGen.un241_ci ));
    InMux I__1019 (
            .O(N__8194),
            .I(N__8191));
    LocalMux I__1018 (
            .O(N__8191),
            .I(\resetGen.reset_count_2_0_4 ));
    InMux I__1017 (
            .O(N__8188),
            .I(N__8176));
    InMux I__1016 (
            .O(N__8187),
            .I(N__8176));
    InMux I__1015 (
            .O(N__8186),
            .I(N__8176));
    InMux I__1014 (
            .O(N__8185),
            .I(N__8176));
    LocalMux I__1013 (
            .O(N__8176),
            .I(\resetGen.escKeyZ0 ));
    CascadeMux I__1012 (
            .O(N__8173),
            .I(N__8167));
    CascadeMux I__1011 (
            .O(N__8172),
            .I(N__8164));
    InMux I__1010 (
            .O(N__8171),
            .I(N__8154));
    InMux I__1009 (
            .O(N__8170),
            .I(N__8154));
    InMux I__1008 (
            .O(N__8167),
            .I(N__8154));
    InMux I__1007 (
            .O(N__8164),
            .I(N__8154));
    InMux I__1006 (
            .O(N__8163),
            .I(N__8151));
    LocalMux I__1005 (
            .O(N__8154),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__1004 (
            .O(N__8151),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__1003 (
            .O(N__8146),
            .I(N__8139));
    InMux I__1002 (
            .O(N__8145),
            .I(N__8139));
    InMux I__1001 (
            .O(N__8144),
            .I(N__8136));
    LocalMux I__1000 (
            .O(N__8139),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__999 (
            .O(N__8136),
            .I(\uu0.l_countZ0Z_3 ));
    InMux I__998 (
            .O(N__8131),
            .I(N__8128));
    LocalMux I__997 (
            .O(N__8128),
            .I(N__8125));
    Odrv4 I__996 (
            .O(N__8125),
            .I(\uu0.un4_l_count_12 ));
    InMux I__995 (
            .O(N__8122),
            .I(N__8118));
    InMux I__994 (
            .O(N__8121),
            .I(N__8115));
    LocalMux I__993 (
            .O(N__8118),
            .I(N__8107));
    LocalMux I__992 (
            .O(N__8115),
            .I(N__8107));
    InMux I__991 (
            .O(N__8114),
            .I(N__8100));
    InMux I__990 (
            .O(N__8113),
            .I(N__8100));
    InMux I__989 (
            .O(N__8112),
            .I(N__8100));
    Odrv4 I__988 (
            .O(N__8107),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__987 (
            .O(N__8100),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__986 (
            .O(N__8095),
            .I(N__8090));
    InMux I__985 (
            .O(N__8094),
            .I(N__8087));
    InMux I__984 (
            .O(N__8093),
            .I(N__8084));
    LocalMux I__983 (
            .O(N__8090),
            .I(N__8081));
    LocalMux I__982 (
            .O(N__8087),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__981 (
            .O(N__8084),
            .I(\uu2.l_countZ0Z_5 ));
    Odrv4 I__980 (
            .O(N__8081),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__979 (
            .O(N__8074),
            .I(N__8067));
    InMux I__978 (
            .O(N__8073),
            .I(N__8067));
    InMux I__977 (
            .O(N__8072),
            .I(N__8064));
    LocalMux I__976 (
            .O(N__8067),
            .I(N__8061));
    LocalMux I__975 (
            .O(N__8064),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    Odrv4 I__974 (
            .O(N__8061),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    InMux I__973 (
            .O(N__8056),
            .I(N__8053));
    LocalMux I__972 (
            .O(N__8053),
            .I(N__8050));
    Odrv4 I__971 (
            .O(N__8050),
            .I(vbuf_tx_data_6));
    InMux I__970 (
            .O(N__8047),
            .I(N__8044));
    LocalMux I__969 (
            .O(N__8044),
            .I(N__8041));
    Odrv4 I__968 (
            .O(N__8041),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__967 (
            .O(N__8038),
            .I(N__8035));
    LocalMux I__966 (
            .O(N__8035),
            .I(N__8032));
    Odrv4 I__965 (
            .O(N__8032),
            .I(vbuf_tx_data_7));
    InMux I__964 (
            .O(N__8029),
            .I(N__8026));
    LocalMux I__963 (
            .O(N__8026),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__962 (
            .O(N__8023),
            .I(N__8019));
    CEMux I__961 (
            .O(N__8022),
            .I(N__8016));
    LocalMux I__960 (
            .O(N__8019),
            .I(N__8013));
    LocalMux I__959 (
            .O(N__8016),
            .I(N__8010));
    Span4Mux_v I__958 (
            .O(N__8013),
            .I(N__8006));
    Span4Mux_v I__957 (
            .O(N__8010),
            .I(N__8003));
    CEMux I__956 (
            .O(N__8009),
            .I(N__8000));
    Odrv4 I__955 (
            .O(N__8006),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__954 (
            .O(N__8003),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    LocalMux I__953 (
            .O(N__8000),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    CascadeMux I__952 (
            .O(N__7993),
            .I(\uu0.un88_ci_3_cascade_ ));
    CascadeMux I__951 (
            .O(N__7990),
            .I(N__7978));
    CascadeMux I__950 (
            .O(N__7989),
            .I(N__7975));
    InMux I__949 (
            .O(N__7988),
            .I(N__7958));
    InMux I__948 (
            .O(N__7987),
            .I(N__7958));
    InMux I__947 (
            .O(N__7986),
            .I(N__7958));
    InMux I__946 (
            .O(N__7985),
            .I(N__7958));
    InMux I__945 (
            .O(N__7984),
            .I(N__7958));
    InMux I__944 (
            .O(N__7983),
            .I(N__7958));
    InMux I__943 (
            .O(N__7982),
            .I(N__7953));
    InMux I__942 (
            .O(N__7981),
            .I(N__7953));
    InMux I__941 (
            .O(N__7978),
            .I(N__7942));
    InMux I__940 (
            .O(N__7975),
            .I(N__7942));
    InMux I__939 (
            .O(N__7974),
            .I(N__7942));
    InMux I__938 (
            .O(N__7973),
            .I(N__7942));
    InMux I__937 (
            .O(N__7972),
            .I(N__7942));
    CascadeMux I__936 (
            .O(N__7971),
            .I(N__7939));
    LocalMux I__935 (
            .O(N__7958),
            .I(N__7930));
    LocalMux I__934 (
            .O(N__7953),
            .I(N__7930));
    LocalMux I__933 (
            .O(N__7942),
            .I(N__7930));
    InMux I__932 (
            .O(N__7939),
            .I(N__7927));
    InMux I__931 (
            .O(N__7938),
            .I(N__7922));
    InMux I__930 (
            .O(N__7937),
            .I(N__7922));
    Span4Mux_v I__929 (
            .O(N__7930),
            .I(N__7919));
    LocalMux I__928 (
            .O(N__7927),
            .I(vbuf_tx_data_rdy));
    LocalMux I__927 (
            .O(N__7922),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__926 (
            .O(N__7919),
            .I(vbuf_tx_data_rdy));
    InMux I__925 (
            .O(N__7912),
            .I(N__7909));
    LocalMux I__924 (
            .O(N__7909),
            .I(N__7906));
    Odrv4 I__923 (
            .O(N__7906),
            .I(\uu2.r_data_wire_2 ));
    InMux I__922 (
            .O(N__7903),
            .I(N__7900));
    LocalMux I__921 (
            .O(N__7900),
            .I(vbuf_tx_data_2));
    InMux I__920 (
            .O(N__7897),
            .I(N__7894));
    LocalMux I__919 (
            .O(N__7894),
            .I(N__7891));
    Odrv4 I__918 (
            .O(N__7891),
            .I(\uu2.r_data_wire_3 ));
    InMux I__917 (
            .O(N__7888),
            .I(N__7885));
    LocalMux I__916 (
            .O(N__7885),
            .I(vbuf_tx_data_3));
    InMux I__915 (
            .O(N__7882),
            .I(N__7879));
    LocalMux I__914 (
            .O(N__7879),
            .I(\uu2.r_data_wire_4 ));
    InMux I__913 (
            .O(N__7876),
            .I(N__7873));
    LocalMux I__912 (
            .O(N__7873),
            .I(vbuf_tx_data_4));
    InMux I__911 (
            .O(N__7870),
            .I(N__7867));
    LocalMux I__910 (
            .O(N__7867),
            .I(\uu2.r_data_wire_5 ));
    InMux I__909 (
            .O(N__7864),
            .I(N__7861));
    LocalMux I__908 (
            .O(N__7861),
            .I(vbuf_tx_data_5));
    InMux I__907 (
            .O(N__7858),
            .I(N__7855));
    LocalMux I__906 (
            .O(N__7855),
            .I(\uu2.r_data_wire_6 ));
    InMux I__905 (
            .O(N__7852),
            .I(N__7849));
    LocalMux I__904 (
            .O(N__7849),
            .I(\uu2.r_data_wire_7 ));
    CEMux I__903 (
            .O(N__7846),
            .I(N__7843));
    LocalMux I__902 (
            .O(N__7843),
            .I(N__7840));
    Span4Mux_v I__901 (
            .O(N__7840),
            .I(N__7837));
    Odrv4 I__900 (
            .O(N__7837),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    InMux I__899 (
            .O(N__7834),
            .I(N__7831));
    LocalMux I__898 (
            .O(N__7831),
            .I(\uu0.sec_clkDZ0 ));
    CascadeMux I__897 (
            .O(N__7828),
            .I(\uu2.un1_l_count_2_2_cascade_ ));
    InMux I__896 (
            .O(N__7825),
            .I(N__7822));
    LocalMux I__895 (
            .O(N__7822),
            .I(\uu2.un284_ci ));
    CascadeMux I__894 (
            .O(N__7819),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__893 (
            .O(N__7816),
            .I(N__7809));
    InMux I__892 (
            .O(N__7815),
            .I(N__7809));
    InMux I__891 (
            .O(N__7814),
            .I(N__7806));
    LocalMux I__890 (
            .O(N__7809),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__889 (
            .O(N__7806),
            .I(\uu2.l_countZ0Z_7 ));
    CascadeMux I__888 (
            .O(N__7801),
            .I(N__7798));
    InMux I__887 (
            .O(N__7798),
            .I(N__7793));
    InMux I__886 (
            .O(N__7797),
            .I(N__7790));
    InMux I__885 (
            .O(N__7796),
            .I(N__7787));
    LocalMux I__884 (
            .O(N__7793),
            .I(N__7784));
    LocalMux I__883 (
            .O(N__7790),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__882 (
            .O(N__7787),
            .I(\uu2.l_countZ0Z_8 ));
    Odrv4 I__881 (
            .O(N__7784),
            .I(\uu2.l_countZ0Z_8 ));
    InMux I__880 (
            .O(N__7777),
            .I(N__7772));
    InMux I__879 (
            .O(N__7776),
            .I(N__7767));
    InMux I__878 (
            .O(N__7775),
            .I(N__7767));
    LocalMux I__877 (
            .O(N__7772),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__876 (
            .O(N__7767),
            .I(\uu2.l_countZ0Z_3 ));
    InMux I__875 (
            .O(N__7762),
            .I(N__7753));
    InMux I__874 (
            .O(N__7761),
            .I(N__7753));
    InMux I__873 (
            .O(N__7760),
            .I(N__7748));
    InMux I__872 (
            .O(N__7759),
            .I(N__7748));
    InMux I__871 (
            .O(N__7758),
            .I(N__7745));
    LocalMux I__870 (
            .O(N__7753),
            .I(N__7742));
    LocalMux I__869 (
            .O(N__7748),
            .I(N__7739));
    LocalMux I__868 (
            .O(N__7745),
            .I(\uu2.l_countZ0Z_6 ));
    Odrv4 I__867 (
            .O(N__7742),
            .I(\uu2.l_countZ0Z_6 ));
    Odrv4 I__866 (
            .O(N__7739),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__865 (
            .O(N__7732),
            .I(N__7727));
    CascadeMux I__864 (
            .O(N__7731),
            .I(N__7724));
    InMux I__863 (
            .O(N__7730),
            .I(N__7717));
    InMux I__862 (
            .O(N__7727),
            .I(N__7717));
    InMux I__861 (
            .O(N__7724),
            .I(N__7717));
    LocalMux I__860 (
            .O(N__7717),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__859 (
            .O(N__7714),
            .I(N__7700));
    InMux I__858 (
            .O(N__7713),
            .I(N__7700));
    InMux I__857 (
            .O(N__7712),
            .I(N__7700));
    InMux I__856 (
            .O(N__7711),
            .I(N__7700));
    InMux I__855 (
            .O(N__7710),
            .I(N__7695));
    InMux I__854 (
            .O(N__7709),
            .I(N__7695));
    LocalMux I__853 (
            .O(N__7700),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__852 (
            .O(N__7695),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__851 (
            .O(N__7690),
            .I(N__7680));
    InMux I__850 (
            .O(N__7689),
            .I(N__7680));
    InMux I__849 (
            .O(N__7688),
            .I(N__7680));
    CascadeMux I__848 (
            .O(N__7687),
            .I(N__7676));
    LocalMux I__847 (
            .O(N__7680),
            .I(N__7673));
    InMux I__846 (
            .O(N__7679),
            .I(N__7668));
    InMux I__845 (
            .O(N__7676),
            .I(N__7668));
    Odrv4 I__844 (
            .O(N__7673),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__843 (
            .O(N__7668),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__842 (
            .O(N__7663),
            .I(N__7654));
    InMux I__841 (
            .O(N__7662),
            .I(N__7654));
    InMux I__840 (
            .O(N__7661),
            .I(N__7647));
    InMux I__839 (
            .O(N__7660),
            .I(N__7647));
    InMux I__838 (
            .O(N__7659),
            .I(N__7647));
    LocalMux I__837 (
            .O(N__7654),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__836 (
            .O(N__7647),
            .I(\uu2.l_countZ0Z_1 ));
    CascadeMux I__835 (
            .O(N__7642),
            .I(\uu2.un1_l_count_1_2_0_cascade_ ));
    InMux I__834 (
            .O(N__7639),
            .I(N__7633));
    InMux I__833 (
            .O(N__7638),
            .I(N__7633));
    LocalMux I__832 (
            .O(N__7633),
            .I(\uu2.un1_l_count_1_3 ));
    CascadeMux I__831 (
            .O(N__7630),
            .I(N__7624));
    InMux I__830 (
            .O(N__7629),
            .I(N__7619));
    InMux I__829 (
            .O(N__7628),
            .I(N__7619));
    InMux I__828 (
            .O(N__7627),
            .I(N__7616));
    InMux I__827 (
            .O(N__7624),
            .I(N__7613));
    LocalMux I__826 (
            .O(N__7619),
            .I(N__7610));
    LocalMux I__825 (
            .O(N__7616),
            .I(\uu2.un306_ci ));
    LocalMux I__824 (
            .O(N__7613),
            .I(\uu2.un306_ci ));
    Odrv4 I__823 (
            .O(N__7610),
            .I(\uu2.un306_ci ));
    InMux I__822 (
            .O(N__7603),
            .I(N__7600));
    LocalMux I__821 (
            .O(N__7600),
            .I(N__7597));
    Odrv4 I__820 (
            .O(N__7597),
            .I(\uu2.r_data_wire_0 ));
    InMux I__819 (
            .O(N__7594),
            .I(N__7591));
    LocalMux I__818 (
            .O(N__7591),
            .I(vbuf_tx_data_0));
    InMux I__817 (
            .O(N__7588),
            .I(N__7585));
    LocalMux I__816 (
            .O(N__7585),
            .I(N__7582));
    Odrv4 I__815 (
            .O(N__7582),
            .I(\uu2.r_data_wire_1 ));
    InMux I__814 (
            .O(N__7579),
            .I(N__7576));
    LocalMux I__813 (
            .O(N__7576),
            .I(vbuf_tx_data_1));
    InMux I__812 (
            .O(N__7573),
            .I(N__7564));
    InMux I__811 (
            .O(N__7572),
            .I(N__7564));
    InMux I__810 (
            .O(N__7571),
            .I(N__7557));
    InMux I__809 (
            .O(N__7570),
            .I(N__7557));
    InMux I__808 (
            .O(N__7569),
            .I(N__7557));
    LocalMux I__807 (
            .O(N__7564),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__806 (
            .O(N__7557),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__805 (
            .O(N__7552),
            .I(N__7549));
    LocalMux I__804 (
            .O(N__7549),
            .I(\buart.Z_tx.un1_bitcount_c3 ));
    InMux I__803 (
            .O(N__7546),
            .I(N__7542));
    InMux I__802 (
            .O(N__7545),
            .I(N__7539));
    LocalMux I__801 (
            .O(N__7542),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__800 (
            .O(N__7539),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__799 (
            .O(N__7534),
            .I(N__7521));
    InMux I__798 (
            .O(N__7533),
            .I(N__7521));
    InMux I__797 (
            .O(N__7532),
            .I(N__7521));
    InMux I__796 (
            .O(N__7531),
            .I(N__7521));
    InMux I__795 (
            .O(N__7530),
            .I(N__7518));
    LocalMux I__794 (
            .O(N__7521),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__793 (
            .O(N__7518),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    InMux I__792 (
            .O(N__7513),
            .I(N__7510));
    LocalMux I__791 (
            .O(N__7510),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ));
    CascadeMux I__790 (
            .O(N__7507),
            .I(N__7503));
    InMux I__789 (
            .O(N__7506),
            .I(N__7495));
    InMux I__788 (
            .O(N__7503),
            .I(N__7495));
    InMux I__787 (
            .O(N__7502),
            .I(N__7495));
    LocalMux I__786 (
            .O(N__7495),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__785 (
            .O(N__7492),
            .I(N__7489));
    InMux I__784 (
            .O(N__7489),
            .I(N__7486));
    LocalMux I__783 (
            .O(N__7486),
            .I(\uu2.un350_ci ));
    CascadeMux I__782 (
            .O(N__7483),
            .I(N__7479));
    InMux I__781 (
            .O(N__7482),
            .I(N__7474));
    InMux I__780 (
            .O(N__7479),
            .I(N__7474));
    LocalMux I__779 (
            .O(N__7474),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__778 (
            .O(N__7471),
            .I(N__7465));
    InMux I__777 (
            .O(N__7470),
            .I(N__7465));
    LocalMux I__776 (
            .O(N__7465),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    InMux I__775 (
            .O(N__7462),
            .I(N__7456));
    InMux I__774 (
            .O(N__7461),
            .I(N__7456));
    LocalMux I__773 (
            .O(N__7456),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__772 (
            .O(N__7453),
            .I(N__7449));
    CascadeMux I__771 (
            .O(N__7452),
            .I(N__7446));
    InMux I__770 (
            .O(N__7449),
            .I(N__7441));
    InMux I__769 (
            .O(N__7446),
            .I(N__7441));
    LocalMux I__768 (
            .O(N__7441),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__767 (
            .O(N__7438),
            .I(N__7435));
    InMux I__766 (
            .O(N__7435),
            .I(N__7429));
    InMux I__765 (
            .O(N__7434),
            .I(N__7429));
    LocalMux I__764 (
            .O(N__7429),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__763 (
            .O(N__7426),
            .I(N__7423));
    LocalMux I__762 (
            .O(N__7423),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__761 (
            .O(N__7420),
            .I(N__7416));
    InMux I__760 (
            .O(N__7419),
            .I(N__7412));
    InMux I__759 (
            .O(N__7416),
            .I(N__7407));
    InMux I__758 (
            .O(N__7415),
            .I(N__7407));
    LocalMux I__757 (
            .O(N__7412),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__756 (
            .O(N__7407),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__755 (
            .O(N__7402),
            .I(N__7394));
    InMux I__754 (
            .O(N__7401),
            .I(N__7394));
    InMux I__753 (
            .O(N__7400),
            .I(N__7389));
    InMux I__752 (
            .O(N__7399),
            .I(N__7389));
    LocalMux I__751 (
            .O(N__7394),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__750 (
            .O(N__7389),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__749 (
            .O(N__7384),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    InMux I__748 (
            .O(N__7381),
            .I(N__7371));
    InMux I__747 (
            .O(N__7380),
            .I(N__7371));
    InMux I__746 (
            .O(N__7379),
            .I(N__7371));
    InMux I__745 (
            .O(N__7378),
            .I(N__7368));
    LocalMux I__744 (
            .O(N__7371),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__743 (
            .O(N__7368),
            .I(\buart.Z_tx.ser_clk ));
    CascadeMux I__742 (
            .O(N__7363),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    InMux I__741 (
            .O(N__7360),
            .I(N__7354));
    InMux I__740 (
            .O(N__7359),
            .I(N__7347));
    InMux I__739 (
            .O(N__7358),
            .I(N__7347));
    InMux I__738 (
            .O(N__7357),
            .I(N__7347));
    LocalMux I__737 (
            .O(N__7354),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__736 (
            .O(N__7347),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__735 (
            .O(N__7342),
            .I(N__7334));
    InMux I__734 (
            .O(N__7341),
            .I(N__7334));
    InMux I__733 (
            .O(N__7340),
            .I(N__7329));
    InMux I__732 (
            .O(N__7339),
            .I(N__7329));
    LocalMux I__731 (
            .O(N__7334),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__730 (
            .O(N__7329),
            .I(\uu0.un154_ci_9 ));
    InMux I__729 (
            .O(N__7324),
            .I(N__7319));
    InMux I__728 (
            .O(N__7323),
            .I(N__7314));
    InMux I__727 (
            .O(N__7322),
            .I(N__7314));
    LocalMux I__726 (
            .O(N__7319),
            .I(N__7311));
    LocalMux I__725 (
            .O(N__7314),
            .I(\uu0.l_countZ0Z_15 ));
    Odrv4 I__724 (
            .O(N__7311),
            .I(\uu0.l_countZ0Z_15 ));
    CascadeMux I__723 (
            .O(N__7306),
            .I(\uu0.un4_l_count_0_8_cascade_ ));
    CascadeMux I__722 (
            .O(N__7303),
            .I(N__7297));
    InMux I__721 (
            .O(N__7302),
            .I(N__7292));
    InMux I__720 (
            .O(N__7301),
            .I(N__7292));
    InMux I__719 (
            .O(N__7300),
            .I(N__7287));
    InMux I__718 (
            .O(N__7297),
            .I(N__7287));
    LocalMux I__717 (
            .O(N__7292),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__716 (
            .O(N__7287),
            .I(\uu0.l_countZ0Z_14 ));
    InMux I__715 (
            .O(N__7282),
            .I(N__7269));
    InMux I__714 (
            .O(N__7281),
            .I(N__7269));
    InMux I__713 (
            .O(N__7280),
            .I(N__7269));
    InMux I__712 (
            .O(N__7279),
            .I(N__7269));
    InMux I__711 (
            .O(N__7278),
            .I(N__7266));
    LocalMux I__710 (
            .O(N__7269),
            .I(N__7263));
    LocalMux I__709 (
            .O(N__7266),
            .I(\uu0.l_precountZ0Z_1 ));
    Odrv12 I__708 (
            .O(N__7263),
            .I(\uu0.l_precountZ0Z_1 ));
    InMux I__707 (
            .O(N__7258),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__706 (
            .O(N__7255),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__705 (
            .O(N__7252),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__704 (
            .O(N__7249),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__703 (
            .O(N__7246),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    InMux I__702 (
            .O(N__7243),
            .I(N__7231));
    InMux I__701 (
            .O(N__7242),
            .I(N__7231));
    InMux I__700 (
            .O(N__7241),
            .I(N__7231));
    InMux I__699 (
            .O(N__7240),
            .I(N__7231));
    LocalMux I__698 (
            .O(N__7231),
            .I(\uu0.l_countZ0Z_10 ));
    InMux I__697 (
            .O(N__7228),
            .I(N__7225));
    LocalMux I__696 (
            .O(N__7225),
            .I(\uu0.un143_ci_0 ));
    InMux I__695 (
            .O(N__7222),
            .I(N__7204));
    InMux I__694 (
            .O(N__7221),
            .I(N__7204));
    InMux I__693 (
            .O(N__7220),
            .I(N__7204));
    InMux I__692 (
            .O(N__7219),
            .I(N__7204));
    InMux I__691 (
            .O(N__7218),
            .I(N__7204));
    InMux I__690 (
            .O(N__7217),
            .I(N__7204));
    LocalMux I__689 (
            .O(N__7204),
            .I(\uu0.l_countZ0Z_8 ));
    CascadeMux I__688 (
            .O(N__7201),
            .I(\uu0.un187_ci_1_cascade_ ));
    CascadeMux I__687 (
            .O(N__7198),
            .I(N__7195));
    InMux I__686 (
            .O(N__7195),
            .I(N__7192));
    LocalMux I__685 (
            .O(N__7192),
            .I(\uu0.un165_ci_0 ));
    InMux I__684 (
            .O(N__7189),
            .I(N__7185));
    InMux I__683 (
            .O(N__7188),
            .I(N__7182));
    LocalMux I__682 (
            .O(N__7185),
            .I(\uu0.l_countZ0Z_13 ));
    LocalMux I__681 (
            .O(N__7182),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__680 (
            .O(N__7177),
            .I(N__7168));
    InMux I__679 (
            .O(N__7176),
            .I(N__7168));
    InMux I__678 (
            .O(N__7175),
            .I(N__7168));
    LocalMux I__677 (
            .O(N__7168),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__676 (
            .O(N__7165),
            .I(N__7160));
    InMux I__675 (
            .O(N__7164),
            .I(N__7155));
    InMux I__674 (
            .O(N__7163),
            .I(N__7155));
    LocalMux I__673 (
            .O(N__7160),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__672 (
            .O(N__7155),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__671 (
            .O(N__7150),
            .I(\uu0.un55_ci_cascade_ ));
    CascadeMux I__670 (
            .O(N__7147),
            .I(N__7140));
    InMux I__669 (
            .O(N__7146),
            .I(N__7126));
    InMux I__668 (
            .O(N__7145),
            .I(N__7126));
    InMux I__667 (
            .O(N__7144),
            .I(N__7126));
    InMux I__666 (
            .O(N__7143),
            .I(N__7126));
    InMux I__665 (
            .O(N__7140),
            .I(N__7126));
    InMux I__664 (
            .O(N__7139),
            .I(N__7126));
    LocalMux I__663 (
            .O(N__7126),
            .I(\uu0.l_countZ0Z_0 ));
    InMux I__662 (
            .O(N__7123),
            .I(N__7110));
    InMux I__661 (
            .O(N__7122),
            .I(N__7110));
    InMux I__660 (
            .O(N__7121),
            .I(N__7110));
    InMux I__659 (
            .O(N__7120),
            .I(N__7110));
    InMux I__658 (
            .O(N__7119),
            .I(N__7107));
    LocalMux I__657 (
            .O(N__7110),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__656 (
            .O(N__7107),
            .I(\uu0.l_countZ0Z_1 ));
    CascadeMux I__655 (
            .O(N__7102),
            .I(N__7098));
    CascadeMux I__654 (
            .O(N__7101),
            .I(N__7095));
    InMux I__653 (
            .O(N__7098),
            .I(N__7086));
    InMux I__652 (
            .O(N__7095),
            .I(N__7086));
    InMux I__651 (
            .O(N__7094),
            .I(N__7086));
    InMux I__650 (
            .O(N__7093),
            .I(N__7083));
    LocalMux I__649 (
            .O(N__7086),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__648 (
            .O(N__7083),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__647 (
            .O(N__7078),
            .I(\uu0.un4_l_count_14_cascade_ ));
    InMux I__646 (
            .O(N__7075),
            .I(N__7072));
    LocalMux I__645 (
            .O(N__7072),
            .I(N__7069));
    Odrv4 I__644 (
            .O(N__7069),
            .I(\uu0.un4_l_count_18 ));
    InMux I__643 (
            .O(N__7066),
            .I(N__7061));
    InMux I__642 (
            .O(N__7065),
            .I(N__7058));
    InMux I__641 (
            .O(N__7064),
            .I(N__7055));
    LocalMux I__640 (
            .O(N__7061),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__639 (
            .O(N__7058),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__638 (
            .O(N__7055),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__637 (
            .O(N__7048),
            .I(\uu0.un154_ci_9_cascade_ ));
    CascadeMux I__636 (
            .O(N__7045),
            .I(N__7040));
    CascadeMux I__635 (
            .O(N__7044),
            .I(N__7037));
    InMux I__634 (
            .O(N__7043),
            .I(N__7030));
    InMux I__633 (
            .O(N__7040),
            .I(N__7030));
    InMux I__632 (
            .O(N__7037),
            .I(N__7030));
    LocalMux I__631 (
            .O(N__7030),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__630 (
            .O(N__7027),
            .I(\uu0.un4_l_count_11_cascade_ ));
    CascadeMux I__629 (
            .O(N__7024),
            .I(\uu0.un4_l_count_16_cascade_ ));
    InMux I__628 (
            .O(N__7021),
            .I(N__7017));
    InMux I__627 (
            .O(N__7020),
            .I(N__7014));
    LocalMux I__626 (
            .O(N__7017),
            .I(\uu0.delay_lineZ0Z_0 ));
    LocalMux I__625 (
            .O(N__7014),
            .I(\uu0.delay_lineZ0Z_0 ));
    CascadeMux I__624 (
            .O(N__7009),
            .I(\uu0.un4_l_count_0_cascade_ ));
    InMux I__623 (
            .O(N__7006),
            .I(N__7003));
    LocalMux I__622 (
            .O(N__7003),
            .I(\uu0.delay_lineZ0Z_1 ));
    IoInMux I__621 (
            .O(N__7000),
            .I(N__6997));
    LocalMux I__620 (
            .O(N__6997),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__619 (
            .O(N__6994),
            .I(N__6988));
    InMux I__618 (
            .O(N__6993),
            .I(N__6981));
    InMux I__617 (
            .O(N__6992),
            .I(N__6981));
    InMux I__616 (
            .O(N__6991),
            .I(N__6981));
    InMux I__615 (
            .O(N__6988),
            .I(N__6978));
    LocalMux I__614 (
            .O(N__6981),
            .I(\uu0.l_precountZ0Z_2 ));
    LocalMux I__613 (
            .O(N__6978),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__612 (
            .O(N__6973),
            .I(N__6970));
    LocalMux I__611 (
            .O(N__6970),
            .I(\uu0.un4_l_count_13 ));
    InMux I__610 (
            .O(N__6967),
            .I(N__6964));
    LocalMux I__609 (
            .O(N__6964),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__608 (
            .O(N__6961),
            .I(N__6958));
    LocalMux I__607 (
            .O(N__6958),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__606 (
            .O(N__6955),
            .I(N__6952));
    LocalMux I__605 (
            .O(N__6952),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__604 (
            .O(N__6949),
            .I(\uu2.un284_ci_cascade_ ));
    CascadeMux I__603 (
            .O(N__6946),
            .I(\uu2.un306_ci_cascade_ ));
    CascadeMux I__602 (
            .O(N__6943),
            .I(\uu2.un350_ci_cascade_ ));
    InMux I__601 (
            .O(N__6940),
            .I(N__6937));
    LocalMux I__600 (
            .O(N__6937),
            .I(N__6934));
    Odrv4 I__599 (
            .O(N__6934),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__598 (
            .O(N__6931),
            .I(N__6928));
    LocalMux I__597 (
            .O(N__6928),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__596 (
            .O(N__6925),
            .I(N__6922));
    LocalMux I__595 (
            .O(N__6922),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__594 (
            .O(N__6919),
            .I(N__6916));
    LocalMux I__593 (
            .O(N__6916),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__592 (
            .O(N__6913),
            .I(N__6910));
    LocalMux I__591 (
            .O(N__6910),
            .I(N__6907));
    IoSpan4Mux I__590 (
            .O(N__6907),
            .I(N__6904));
    Odrv4 I__589 (
            .O(N__6904),
            .I(o_serial_data_c));
    IoInMux I__588 (
            .O(N__6901),
            .I(N__6898));
    LocalMux I__587 (
            .O(N__6898),
            .I(N__6895));
    Span12Mux_s5_h I__586 (
            .O(N__6895),
            .I(N__6892));
    Span12Mux_v I__585 (
            .O(N__6892),
            .I(N__6889));
    Odrv12 I__584 (
            .O(N__6889),
            .I(clk_in_c));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__18050));
    INV \INVuu2.w_addr_displaying_nesr_5C  (
            .O(\INVuu2.w_addr_displaying_nesr_5C_net ),
            .I(N__18056));
    INV \INVuu2.bitmap_215C  (
            .O(\INVuu2.bitmap_215C_net ),
            .I(N__18044));
    INV \INVuu2.w_addr_displaying_nesr_8C  (
            .O(\INVuu2.w_addr_displaying_nesr_8C_net ),
            .I(N__18055));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__18067));
    INV \INVuu2.bitmap_168C  (
            .O(\INVuu2.bitmap_168C_net ),
            .I(N__18024));
    INV \INVuu2.bitmap_200C  (
            .O(\INVuu2.bitmap_200C_net ),
            .I(N__18029));
    INV \INVuu2.w_addr_displaying_fast_nesr_8C  (
            .O(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .I(N__18033));
    INV \INVuu2.w_addr_displaying_2_rep1C  (
            .O(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .I(N__18040));
    INV \INVuu2.w_addr_displaying_4C  (
            .O(\INVuu2.w_addr_displaying_4C_net ),
            .I(N__18052));
    INV \INVuu2.w_addr_user_nesr_6C  (
            .O(\INVuu2.w_addr_user_nesr_6C_net ),
            .I(N__18058));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__18031));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__18036));
    INV \INVuu2.bitmap_197C  (
            .O(\INVuu2.bitmap_197C_net ),
            .I(N__18061));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__18035));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__18043));
    INV \INVuu2.bitmap_186C  (
            .O(\INVuu2.bitmap_186C_net ),
            .I(N__18049));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__18072));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__8712),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__7000),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__17647),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \buart.Z_tx.shifter_0_LC_1_5_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_1_5_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_1_5_2  (
            .in0(N__7982),
            .in1(N__6940),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18094),
            .ce(N__8009),
            .sr(N__17820));
    defparam \buart.Z_tx.uart_tx_LC_1_5_7 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_1_5_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_1_5_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.uart_tx_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__7981),
            .in2(_gnd_net_),
            .in3(N__6919),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18094),
            .ce(N__8009),
            .sr(N__17820));
    defparam \uu2.l_count_7_LC_1_6_0 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_1_6_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_1_6_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.l_count_7_LC_1_6_0  (
            .in0(N__8074),
            .in1(N__7762),
            .in2(N__7630),
            .in3(N__7816),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18088),
            .ce(),
            .sr(N__17817));
    defparam \uu2.l_count_1_LC_1_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_1_6_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_1_LC_1_6_1  (
            .in0(N__7661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7714),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18088),
            .ce(),
            .sr(N__17817));
    defparam \uu2.l_count_0_LC_1_6_2 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_1_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uu2.l_count_0_LC_1_6_2  (
            .in0(N__7713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18088),
            .ce(),
            .sr(N__17817));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_6_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_6_3  (
            .in0(N__7660),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7712),
            .lcout(\uu2.un284_ci ),
            .ltout(\uu2.un284_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_1_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_1_6_4 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_1_6_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.l_count_2_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6949),
            .in3(N__7679),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18088),
            .ce(),
            .sr(N__17817));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_5  (
            .in0(N__7659),
            .in1(N__7711),
            .in2(N__7687),
            .in3(N__7777),
            .lcout(\uu2.un306_ci ),
            .ltout(\uu2.un306_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_6_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_6_6  (
            .in0(N__8073),
            .in1(N__7761),
            .in2(N__6946),
            .in3(N__7815),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_1_6_7 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_1_6_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_1_6_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.l_count_8_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6943),
            .in3(N__7796),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18088),
            .ce(),
            .sr(N__17817));
    defparam \buart.Z_tx.shifter_1_LC_1_7_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_1_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_1_7_0  (
            .in0(N__7983),
            .in1(N__6931),
            .in2(_gnd_net_),
            .in3(N__7594),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \buart.Z_tx.shifter_2_LC_1_7_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_1_7_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_1_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_1_7_3  (
            .in0(N__6925),
            .in1(N__7986),
            .in2(_gnd_net_),
            .in3(N__7579),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \buart.Z_tx.shifter_3_LC_1_7_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_1_7_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_1_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_1_7_4  (
            .in0(N__7984),
            .in1(N__6967),
            .in2(_gnd_net_),
            .in3(N__7903),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \buart.Z_tx.shifter_4_LC_1_7_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_1_7_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_1_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \buart.Z_tx.shifter_4_LC_1_7_5  (
            .in0(N__7888),
            .in1(N__6961),
            .in2(_gnd_net_),
            .in3(N__7988),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \buart.Z_tx.shifter_5_LC_1_7_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_1_7_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_1_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_1_7_6  (
            .in0(N__7985),
            .in1(N__6955),
            .in2(_gnd_net_),
            .in3(N__7876),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \buart.Z_tx.shifter_6_LC_1_7_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_1_7_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_1_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_1_7_7  (
            .in0(N__8047),
            .in1(N__7987),
            .in2(_gnd_net_),
            .in3(N__7864),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18078),
            .ce(N__8022),
            .sr(N__17814));
    defparam \uu2.l_count_5_LC_1_8_0 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_1_8_0 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.l_count_5_LC_1_8_0  (
            .in0(N__8094),
            .in1(N__8122),
            .in2(_gnd_net_),
            .in3(N__7629),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \uu2.l_count_6_LC_1_8_1 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_1_8_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_1_8_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_6_LC_1_8_1  (
            .in0(N__7628),
            .in1(N__8072),
            .in2(_gnd_net_),
            .in3(N__7758),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \Lab_UT.dispString.cnt_1_LC_1_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_1_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_1_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_1_8_2  (
            .in0(N__15290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15206),
            .lcout(\Lab_UT.cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \Lab_UT.dispString.cnt_0_LC_1_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_1_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_1_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_1_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15289),
            .lcout(\Lab_UT.cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \uu0.sec_clk_LC_1_8_4 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_1_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__9195),
            .in2(_gnd_net_),
            .in3(N__8591),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \uu0.delay_line_1_LC_1_8_7 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_1_8_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uu0.delay_line_1_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(N__7021),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18071),
            .ce(),
            .sr(N__17805));
    defparam \uu0.delay_line_0_LC_1_9_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_9_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_9_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_9_0  (
            .in0(N__7280),
            .in1(N__9101),
            .in2(N__7045),
            .in3(N__6991),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18065),
            .ce(),
            .sr(N__17815));
    defparam \uu0.l_precount_3_LC_1_9_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_9_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_9_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_9_1  (
            .in0(N__6993),
            .in1(N__7043),
            .in2(N__9106),
            .in3(N__7282),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18065),
            .ce(),
            .sr(N__17815));
    defparam \uu0.l_precount_2_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_9_2 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_1_9_2  (
            .in0(N__7281),
            .in1(N__9102),
            .in2(_gnd_net_),
            .in3(N__6992),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18065),
            .ce(),
            .sr(N__17815));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_4 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_9_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_9_4  (
            .in0(N__7279),
            .in1(N__8457),
            .in2(N__7044),
            .in3(N__7119),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI96A32_18_LC_1_9_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI96A32_18_LC_1_9_5  (
            .in0(N__7324),
            .in1(N__8662),
            .in2(N__7027),
            .in3(N__8541),
            .lcout(),
            .ltout(\uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_9_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_11_LC_1_9_6  (
            .in0(N__6973),
            .in1(N__8131),
            .in2(N__7024),
            .in3(N__7075),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_9_7 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_9_7 .LUT_INIT=16'b1111000011111010;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_1_9_7  (
            .in0(N__7020),
            .in1(_gnd_net_),
            .in2(N__7009),
            .in3(N__7006),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2CNU_11_LC_1_10_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_10_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uu0.l_count_RNI2CNU_11_LC_1_10_0  (
            .in0(N__8341),
            .in1(N__7064),
            .in2(N__6994),
            .in3(N__7139),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_10_1  (
            .in0(N__8145),
            .in1(N__7094),
            .in2(N__7147),
            .in3(N__7120),
            .lcout(\uu0.un66_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_10_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_10_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_10_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uu0.l_count_2_LC_1_10_2  (
            .in0(N__7123),
            .in1(_gnd_net_),
            .in2(N__7102),
            .in3(N__7146),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18059),
            .ce(N__8297),
            .sr(N__17816));
    defparam \uu0.l_count_0_LC_1_10_3 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_10_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_10_3  (
            .in0(N__7144),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8588),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18059),
            .ce(N__8297),
            .sr(N__17816));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_10_4  (
            .in0(N__7121),
            .in1(_gnd_net_),
            .in2(N__7101),
            .in3(N__7143),
            .lcout(),
            .ltout(\uu0.un55_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_3_LC_1_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_10_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \uu0.l_count_3_LC_1_10_5  (
            .in0(N__8146),
            .in1(_gnd_net_),
            .in2(N__7150),
            .in3(N__8590),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18059),
            .ce(N__8297),
            .sr(N__17816));
    defparam \uu0.l_count_1_LC_1_10_6 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_10_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_1_10_6  (
            .in0(N__7122),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7145),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18059),
            .ce(N__8297),
            .sr(N__17816));
    defparam \uu0.l_count_11_LC_1_10_7 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_1_10_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_1_10_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_11_LC_1_10_7  (
            .in0(N__7228),
            .in1(N__7066),
            .in2(N__8407),
            .in3(N__8589),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18059),
            .ce(N__8297),
            .sr(N__17816));
    defparam \uu0.l_count_RNI04591_10_LC_1_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI04591_10_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI04591_10_LC_1_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_count_RNI04591_10_LC_1_11_0  (
            .in0(N__7240),
            .in1(N__7217),
            .in2(N__7303),
            .in3(N__7093),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2GS72_4_LC_1_11_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_11_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNI2GS72_4_LC_1_11_1  (
            .in0(N__9099),
            .in1(N__8487),
            .in2(N__7078),
            .in3(N__7163),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_11_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_11_2  (
            .in0(N__7241),
            .in1(N__7065),
            .in2(N__8172),
            .in3(N__7218),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_1_11_3 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_11_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_1_11_3  (
            .in0(N__8382),
            .in1(N__7300),
            .in2(N__7048),
            .in3(N__7164),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18053),
            .ce(N__8298),
            .sr(N__17819));
    defparam \uu0.l_count_8_LC_1_11_4 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_11_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_count_8_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__8383),
            .in2(_gnd_net_),
            .in3(N__7221),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18053),
            .ce(N__8298),
            .sr(N__17819));
    defparam \uu0.l_count_10_LC_1_11_5 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_11_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_10_LC_1_11_5  (
            .in0(N__7220),
            .in1(N__8170),
            .in2(N__8405),
            .in3(N__7243),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18053),
            .ce(N__8298),
            .sr(N__17819));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_11_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_11_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_11_6  (
            .in0(N__7242),
            .in1(_gnd_net_),
            .in2(N__8173),
            .in3(N__7219),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_9_LC_1_11_7 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_1_11_7 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu0.l_count_9_LC_1_11_7  (
            .in0(N__7222),
            .in1(_gnd_net_),
            .in2(N__8404),
            .in3(N__8171),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18053),
            .ce(N__8298),
            .sr(N__17819));
    defparam \uu0.l_count_13_LC_1_12_0 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_12_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_12_0 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uu0.l_count_13_LC_1_12_0  (
            .in0(N__8597),
            .in1(N__7189),
            .in2(N__7198),
            .in3(N__8420),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18047),
            .ce(N__8299),
            .sr(N__17822));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_12_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_12_1  (
            .in0(N__7302),
            .in1(N__7340),
            .in2(_gnd_net_),
            .in3(N__7165),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_12_2 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_12_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_15_LC_1_12_2  (
            .in0(N__8421),
            .in1(N__8599),
            .in2(N__7201),
            .in3(N__7323),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18047),
            .ce(N__8299),
            .sr(N__17822));
    defparam \uu0.l_count_12_LC_1_12_3 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_12_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_12_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_12_LC_1_12_3  (
            .in0(N__7342),
            .in1(N__8596),
            .in2(N__8422),
            .in3(N__7177),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18047),
            .ce(N__8299),
            .sr(N__17822));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_12_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_12_4  (
            .in0(N__7176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7341),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_12_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_12_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_1_12_5  (
            .in0(_gnd_net_),
            .in1(N__7188),
            .in2(_gnd_net_),
            .in3(N__7175),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(\uu0.un4_l_count_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_12_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_12_6  (
            .in0(N__7339),
            .in1(N__7322),
            .in2(N__7306),
            .in3(N__7301),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_4_LC_1_12_7 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_12_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \uu0.l_count_4_LC_1_12_7  (
            .in0(N__8517),
            .in1(N__8598),
            .in2(_gnd_net_),
            .in3(N__8485),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18047),
            .ce(N__8299),
            .sr(N__17822));
    defparam \uu0.l_precount_1_LC_1_13_5 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_13_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_13_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_precount_1_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__9100),
            .in2(_gnd_net_),
            .in3(N__7278),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18041),
            .ce(),
            .sr(N__17824));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_2_3_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_2_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__7400),
            .in2(N__7420),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_2_3_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_2_3_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_2_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_2_3_1  (
            .in0(_gnd_net_),
            .in1(N__7482),
            .in2(_gnd_net_),
            .in3(N__7258),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__18097),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_2_3_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_2_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_2_3_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_2_3_2  (
            .in0(N__7380),
            .in1(_gnd_net_),
            .in2(N__7438),
            .in3(N__7255),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__18097),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_2_3_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_2_3_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_2_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(N__7462),
            .in2(_gnd_net_),
            .in3(N__7252),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__18097),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_2_3_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_2_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_2_3_4  (
            .in0(N__7381),
            .in1(N__7471),
            .in2(_gnd_net_),
            .in3(N__7249),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__18097),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_2_3_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_2_3_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_2_3_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(N__7379),
            .in2(N__7453),
            .in3(N__7246),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18097),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_2_3_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_2_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_2_3_6  (
            .in0(N__7415),
            .in1(N__7399),
            .in2(N__7483),
            .in3(N__7426),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_2_3_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_2_3_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_2_3_7  (
            .in0(N__7470),
            .in1(N__7461),
            .in2(N__7452),
            .in3(N__7434),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_2_4_0 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_2_4_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_2_4_0  (
            .in0(N__7402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7419),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18095),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_2_4_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_2_4_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7401),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18095),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_4_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_2_4_3 .LUT_INIT=16'b1110000111110000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_2_4_3  (
            .in0(N__7570),
            .in1(N__7358),
            .in2(N__7507),
            .in3(N__7530),
            .lcout(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_4_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_4_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__7569),
            .in2(_gnd_net_),
            .in3(N__7545),
            .lcout(),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_4_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_4_5 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_2_4_5  (
            .in0(N__7502),
            .in1(N__7357),
            .in2(N__7384),
            .in3(N__7378),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_2_4_6  (
            .in0(N__7359),
            .in1(N__7571),
            .in2(N__7363),
            .in3(N__7506),
            .lcout(\buart.Z_tx.un1_bitcount_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_2_5_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_2_5_0 .LUT_INIT=16'b1111110111110010;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_2_5_0  (
            .in0(N__7533),
            .in1(N__7573),
            .in2(N__7989),
            .in3(N__7360),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \buart.Z_tx.bitcount_0_LC_2_5_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_2_5_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_2_5_1  (
            .in0(N__7572),
            .in1(N__7974),
            .in2(_gnd_net_),
            .in3(N__7532),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \buart.Z_tx.bitcount_3_LC_2_5_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_2_5_2 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_2_5_2  (
            .in0(N__7534),
            .in1(N__7546),
            .in2(N__7990),
            .in3(N__7552),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_5_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_5_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_2_5_3  (
            .in0(_gnd_net_),
            .in1(N__7972),
            .in2(_gnd_net_),
            .in3(N__7531),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_2_5_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_2_5_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_2_5_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_2_5_4  (
            .in0(N__7973),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7513),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \uu2.r_addr_2_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_2_5_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_2_LC_2_5_5  (
            .in0(N__9328),
            .in1(N__9371),
            .in2(N__8794),
            .in3(N__9256),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \uu2.r_addr_1_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_2_5_6 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.r_addr_1_LC_2_5_6  (
            .in0(N__9255),
            .in1(N__8790),
            .in2(_gnd_net_),
            .in3(N__9327),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \uu2.r_addr_0_LC_2_5_7 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_2_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_2_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.r_addr_0_LC_2_5_7  (
            .in0(_gnd_net_),
            .in1(N__8789),
            .in2(_gnd_net_),
            .in3(N__9254),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18089),
            .ce(),
            .sr(N__17806));
    defparam \uu2.l_count_9_LC_2_6_0 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_2_6_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_2_6_0 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \uu2.l_count_9_LC_2_6_0  (
            .in0(N__8754),
            .in1(N__7730),
            .in2(N__7492),
            .in3(N__7797),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18079),
            .ce(),
            .sr(N__17821));
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_6_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_2_6_1  (
            .in0(N__7760),
            .in1(N__8113),
            .in2(N__7732),
            .in3(N__7710),
            .lcout(),
            .ltout(\uu2.un1_l_count_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_2_6_2  (
            .in0(N__7689),
            .in1(N__7663),
            .in2(N__7828),
            .in3(N__7638),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_3_LC_2_6_3 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_2_6_3 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_2_6_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \uu2.l_count_3_LC_2_6_3  (
            .in0(N__7776),
            .in1(N__7825),
            .in2(N__7819),
            .in3(N__7690),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18079),
            .ce(),
            .sr(N__17821));
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_2_6_4  (
            .in0(N__7814),
            .in1(N__8095),
            .in2(N__7801),
            .in3(N__7775),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_6_5 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_6_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_2_6_5  (
            .in0(N__7759),
            .in1(N__8112),
            .in2(N__7731),
            .in3(N__7709),
            .lcout(),
            .ltout(\uu2.un1_l_count_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_6 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_2_6_6  (
            .in0(N__7688),
            .in1(N__7662),
            .in2(N__7642),
            .in3(N__7639),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_2_6_7 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_2_6_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_2_6_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu2.l_count_4_LC_2_6_7  (
            .in0(N__7627),
            .in1(N__8114),
            .in2(_gnd_net_),
            .in3(N__8753),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18079),
            .ce(),
            .sr(N__17821));
    defparam \uu2.r_data_reg_0_LC_2_7_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_0_LC_2_7_0  (
            .in0(N__7603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_7_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_1_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7588),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_7_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_2_LC_2_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7912),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_7_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_3_LC_2_7_3  (
            .in0(N__7897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_7_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7882),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_7_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_5_LC_2_7_5  (
            .in0(N__7870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_7_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7858),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_7_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7852),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__7846),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_8_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_8_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_2_8_1  (
            .in0(N__9118),
            .in1(N__9136),
            .in2(_gnd_net_),
            .in3(N__17852),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_2_8_2 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_2_8_2 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_2_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.sec_clkD_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9194),
            .lcout(\uu0.sec_clkDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18066),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_4 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__7834),
            .in2(_gnd_net_),
            .in3(N__9193),
            .lcout(oneSecStrb_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__8121),
            .in2(_gnd_net_),
            .in3(N__8093),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_2_9_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_9_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_9_0  (
            .in0(N__7937),
            .in1(N__8029),
            .in2(_gnd_net_),
            .in3(N__8056),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18060),
            .ce(N__8023),
            .sr(N__17818));
    defparam \buart.Z_tx.shifter_8_LC_2_9_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_9_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_9_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__7938),
            .in2(_gnd_net_),
            .in3(N__8038),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18060),
            .ce(N__8023),
            .sr(N__17818));
    defparam \resetGen.reset_count_RNO_0_4_LC_2_9_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_2_9_3  (
            .in0(N__8219),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8268),
            .lcout(\resetGen.reset_count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_9_4 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_9_4  (
            .in0(N__8237),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8254),
            .lcout(\resetGen.un241_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__8491),
            .in2(_gnd_net_),
            .in3(N__8458),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(\uu0.un88_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_9_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7993),
            .in3(N__8542),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_2_10_0 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_2_10_0 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_2_10_0  (
            .in0(N__9172),
            .in1(N__8829),
            .in2(N__7971),
            .in3(N__17855),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_2_10_1 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_2_10_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.escKey_LC_2_10_1  (
            .in0(N__10297),
            .in1(N__11809),
            .in2(_gnd_net_),
            .in3(N__14017),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(\resetGen.escKeyZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_2_10_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_2_10_2 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \resetGen.reset_count_0_LC_2_10_2  (
            .in0(N__8256),
            .in1(_gnd_net_),
            .in2(N__8278),
            .in3(N__13937),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_10_3 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_10_3  (
            .in0(N__8238),
            .in1(N__8255),
            .in2(_gnd_net_),
            .in3(N__8220),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_2_10_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_2_10_4 .LUT_INIT=16'b0100010000010100;
    LogicCell40 \resetGen.reset_count_3_LC_2_10_4  (
            .in0(N__8187),
            .in1(N__8272),
            .in2(N__8275),
            .in3(N__13939),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_2_10_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_2_10_5 .LUT_INIT=16'b0000000010100110;
    LogicCell40 \resetGen.reset_count_1_LC_2_10_5  (
            .in0(N__8239),
            .in1(N__8257),
            .in2(N__13947),
            .in3(N__8185),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_2_10_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_2_10_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_2_10_6 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \resetGen.reset_count_2_LC_2_10_6  (
            .in0(N__8186),
            .in1(N__13938),
            .in2(N__8224),
            .in3(N__8205),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_2_10_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_2_10_7 .LUT_INIT=16'b0000000011111000;
    LogicCell40 \resetGen.reset_count_4_LC_2_10_7  (
            .in0(N__8206),
            .in1(N__8194),
            .in2(N__13946),
            .in3(N__8188),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18054),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_11_0  (
            .in0(N__8163),
            .in1(N__8633),
            .in2(N__8323),
            .in3(N__8144),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_2_11_1 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_2_11_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_2_11_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_16_LC_2_11_1  (
            .in0(N__8436),
            .in1(N__8593),
            .in2(N__8406),
            .in3(N__8343),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18048),
            .ce(N__8300),
            .sr(N__17823));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2  (
            .in0(N__8514),
            .in1(N__8539),
            .in2(N__8622),
            .in3(N__8634),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3  (
            .in0(N__8435),
            .in1(N__8322),
            .in2(N__8668),
            .in3(N__8342),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_11_4 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_11_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \uu0.l_count_18_LC_2_11_4  (
            .in0(N__8592),
            .in1(_gnd_net_),
            .in2(N__8665),
            .in3(N__8661),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18048),
            .ce(N__8300),
            .sr(N__17823));
    defparam \uu0.l_count_7_LC_2_11_5 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_2_11_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_2_11_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_7_LC_2_11_5  (
            .in0(N__8635),
            .in1(N__8516),
            .in2(N__8647),
            .in3(N__8595),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18048),
            .ce(N__8300),
            .sr(N__17823));
    defparam \uu0.l_count_6_LC_2_11_7 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_2_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_2_11_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_6_LC_2_11_7  (
            .in0(N__8540),
            .in1(N__8515),
            .in2(N__8623),
            .in3(N__8594),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18048),
            .ce(N__8300),
            .sr(N__17823));
    defparam \uu0.l_count_5_LC_2_12_0 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_2_12_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_2_12_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_5_LC_2_12_0  (
            .in0(N__8518),
            .in1(N__8486),
            .in2(_gnd_net_),
            .in3(N__8456),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18042),
            .ce(N__8301),
            .sr(N__17825));
    defparam \uu0.l_count_17_LC_2_13_3 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_13_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_13_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_17_LC_2_13_3  (
            .in0(N__8437),
            .in1(N__8318),
            .in2(N__8416),
            .in3(N__8347),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18034),
            .ce(N__8302),
            .sr(N__17826));
    defparam CONSTANT_ONE_LUT4_LC_4_3_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_4_3_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_4_3_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_4_3_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_5_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_4_4_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_5_LC_4_4_0  (
            .in0(N__9219),
            .in1(N__9522),
            .in2(N__8788),
            .in3(N__9488),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18082),
            .ce(),
            .sr(N__17807));
    defparam \uu2.r_addr_4_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_4_1 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_4_4_1  (
            .in0(N__9521),
            .in1(N__8776),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18082),
            .ce(),
            .sr(N__17807));
    defparam \uu2.trig_rd_det_0_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_4_4_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__9157),
            .in2(_gnd_net_),
            .in3(N__8830),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18082),
            .ce(),
            .sr(N__17807));
    defparam \uu2.trig_rd_det_1_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_4_4_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.trig_rd_det_1_LC_4_4_3  (
            .in0(N__8803),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18082),
            .ce(),
            .sr(N__17807));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__8809),
            .in2(_gnd_net_),
            .in3(N__8802),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(\uu2.trig_rd_is_det_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_4_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8758),
            .in3(N__17854),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_4_4_6 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_4_4_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__9158),
            .in2(_gnd_net_),
            .in3(N__8755),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18082),
            .ce(),
            .sr(N__17807));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_4_5_0  (
            .in0(N__10686),
            .in1(N__12322),
            .in2(_gnd_net_),
            .in3(N__13071),
            .lcout(\uu2.mem0.N_77_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_21_LC_4_5_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_21_LC_4_5_1  (
            .in0(N__14706),
            .in1(N__14995),
            .in2(_gnd_net_),
            .in3(N__12378),
            .lcout(),
            .ltout(\uu2.mem0.w_data_i_a3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_5_2 .LUT_INIT=16'b0011101100010001;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_5_2  (
            .in0(N__12412),
            .in1(N__8878),
            .in2(N__8725),
            .in3(N__12466),
            .lcout(\uu2.mem0.N_79_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_4_5_3 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_4_5_3 .LUT_INIT=16'b1100111110001111;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_4_5_3  (
            .in0(N__12439),
            .in1(N__12409),
            .in2(N__8716),
            .in3(N__12379),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_5_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_5_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_4_5_4  (
            .in0(N__12323),
            .in1(N__11938),
            .in2(_gnd_net_),
            .in3(N__13628),
            .lcout(\uu2.mem0.N_75_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIUGNM6_2_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIUGNM6_2_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIUGNM6_2_LC_4_5_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.w_addr_displaying_RNIUGNM6_2_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__10908),
            .in2(_gnd_net_),
            .in3(N__10955),
            .lcout(\uu2.N_361 ),
            .ltout(\uu2.N_361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_5_6 .LUT_INIT=16'b1010111100001101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_5_6  (
            .in0(N__12411),
            .in1(N__8854),
            .in2(N__8872),
            .in3(N__14659),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_5_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_4_5_7  (
            .in0(N__14707),
            .in1(N__10633),
            .in2(_gnd_net_),
            .in3(N__12410),
            .lcout(\uu2.mem0.N_69_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_22_LC_4_6_0  (
            .in0(N__14685),
            .in1(N__14733),
            .in2(N__12435),
            .in3(N__14790),
            .lcout(\uu2.mem0.w_data_0_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_8_LC_4_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_8_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIFOBB3_8_LC_4_6_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIFOBB3_8_LC_4_6_1  (
            .in0(N__13317),
            .in1(N__10884),
            .in2(N__13627),
            .in3(N__13829),
            .lcout(\uu2.N_61 ),
            .ltout(\uu2.N_61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_2 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__10909),
            .in2(N__8848),
            .in3(N__10956),
            .lcout(),
            .ltout(\uu2.mem0.un51_w_data_displaying_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_6_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_6_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_6_3  (
            .in0(N__14734),
            .in1(_gnd_net_),
            .in2(N__8845),
            .in3(N__12344),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_6_4 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_4_6_4  (
            .in0(N__14686),
            .in1(N__12239),
            .in2(N__12349),
            .in3(N__10957),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_4_6_6  (
            .in0(N__10009),
            .in1(N__12339),
            .in2(_gnd_net_),
            .in3(N__13507),
            .lcout(\uu2.mem0.N_71_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_6_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_6_7 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_6_7  (
            .in0(N__13084),
            .in1(N__14991),
            .in2(N__12348),
            .in3(N__9604),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_4_7_2  (
            .in0(N__12343),
            .in1(N__11884),
            .in2(_gnd_net_),
            .in3(N__12978),
            .lcout(\uu2.mem0.N_76_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_4_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIDKOL_1_LC_4_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_RNIDKOL_1_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__13070),
            .in2(_gnd_net_),
            .in3(N__12895),
            .lcout(\uu2.N_48_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_i_m4_4_LC_4_7_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_i_m4_4_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_i_m4_4_LC_4_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.bcd2segment4.segment_i_m4_4_LC_4_7_6  (
            .in0(N__15512),
            .in1(N__17474),
            .in2(_gnd_net_),
            .in3(N__14943),
            .lcout(\Lab_UT.bcd2segment4.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_4_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_26_LC_4_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_26_LC_4_8_0  (
            .in0(N__8965),
            .in1(N__9907),
            .in2(_gnd_net_),
            .in3(N__8896),
            .lcout(),
            .ltout(\uu2.mem0.N_2166_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_8_1 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_4_8_1  (
            .in0(N__10981),
            .in1(N__8971),
            .in2(N__8914),
            .in3(N__9619),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_8_2 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_8_2  (
            .in0(N__12338),
            .in1(N__10834),
            .in2(N__8911),
            .in3(N__14794),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_4_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_42_LC_4_8_3 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_42_LC_4_8_3  (
            .in0(N__9711),
            .in1(N__10176),
            .in2(N__9670),
            .in3(N__9780),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_4_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_27_LC_4_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_27_LC_4_8_4  (
            .in0(N__9772),
            .in1(N__11125),
            .in2(_gnd_net_),
            .in3(N__9595),
            .lcout(\uu2.mem0.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_25_LC_4_8_5 .LUT_INIT=16'b0110000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_25_LC_4_8_5  (
            .in0(N__13316),
            .in1(N__13502),
            .in2(N__9742),
            .in3(N__9640),
            .lcout(\uu2.mem0.g1_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_4_8_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_43_LC_4_8_6 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_43_LC_4_8_6  (
            .in0(N__10177),
            .in1(N__9666),
            .in2(N__9784),
            .in3(N__9712),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_4_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_6_LC_4_9_0 .LUT_INIT=16'b1110110011000011;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_6_LC_4_9_0  (
            .in0(N__16500),
            .in1(N__16417),
            .in2(N__16647),
            .in3(N__16574),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_4_9_1 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_4_9_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_186_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8956),
            .in3(N__14241),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__17776));
    defparam \uu2.bitmap_RNIMQ601_58_LC_4_9_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIMQ601_58_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIMQ601_58_LC_4_9_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.bitmap_RNIMQ601_58_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__10765),
            .in2(N__9880),
            .in3(N__8947),
            .lcout(),
            .ltout(\uu2.bitmap_RNIMQ601Z0Z_58_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_nesr_RNIV0V92_7_LC_4_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIV0V92_7_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIV0V92_7_LC_4_9_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_RNIV0V92_7_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__11206),
            .in2(N__8953),
            .in3(N__9001),
            .lcout(\uu2.w_addr_displaying_fast_nesr_RNIV0V92Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_4_9_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_0_LC_4_9_4 .LUT_INIT=16'b1111011101101101;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_0_LC_4_9_4  (
            .in0(N__16501),
            .in1(N__16418),
            .in2(N__16648),
            .in3(N__16575),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segment_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_58_LC_4_9_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_4_9_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_4_9_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_58_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8950),
            .in3(N__14242),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__17776));
    defparam \uu2.bitmap_RNI8LB51_186_LC_4_9_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI8LB51_186_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI8LB51_186_LC_4_9_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.bitmap_RNI8LB51_186_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__10764),
            .in2(N__9879),
            .in3(N__9007),
            .lcout(\uu2.bitmap_RNI8LB51Z0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_4_9_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_0_2_LC_4_9_7 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \Lab_UT.bcd2segment1.segment_0_2_LC_4_9_7  (
            .in0(N__16573),
            .in1(N__16636),
            .in2(N__16420),
            .in3(N__16499),
            .lcout(\Lab_UT.bcd2segment1.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_3_LC_4_10_0 .LUT_INIT=16'b1111111010010010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_3_LC_4_10_0  (
            .in0(N__16643),
            .in1(N__16566),
            .in2(N__16502),
            .in3(N__16408),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_314_LC_4_10_1 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_4_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_4_10_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_314_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8995),
            .in3(N__14230),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__17778));
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_4_LC_4_10_2 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_4_LC_4_10_2  (
            .in0(N__16644),
            .in1(N__16567),
            .in2(N__16503),
            .in3(N__16409),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_218_LC_4_10_3 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_4_10_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_4_10_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_218_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8992),
            .in3(N__14229),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__17778));
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_4_10_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segmentUQ_5_LC_4_10_4 .LUT_INIT=16'b1110111011010100;
    LogicCell40 \Lab_UT.bcd2segment1.segmentUQ_5_LC_4_10_4  (
            .in0(N__16645),
            .in1(N__16568),
            .in2(N__16504),
            .in3(N__16410),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segmentUQ_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_90_LC_4_10_5 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_4_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_4_10_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_90_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8989),
            .in3(N__14231),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__17778));
    defparam \uu2.bitmap_RNIARM01_90_LC_4_10_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIARM01_90_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIARM01_90_LC_4_10_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNIARM01_90_LC_4_10_6  (
            .in0(N__8986),
            .in1(N__12894),
            .in2(N__8980),
            .in3(N__10822),
            .lcout(\uu2.bitmap_pmux_19_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_4_11_0 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_4_11_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_4_11_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.bitmap_308_LC_4_11_0  (
            .in0(N__14238),
            .in1(N__11314),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__17779));
    defparam \uu2.bitmap_52_LC_4_11_1 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_4_11_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.bitmap_52_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__14237),
            .in2(_gnd_net_),
            .in3(N__11140),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__17779));
    defparam \uu2.bitmap_111_LC_4_11_2 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_4_11_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9199),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__17779));
    defparam \uu2.vram_rd_clk_det_0_LC_4_11_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_4_11_3 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_4_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9168),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__17779));
    defparam \uu2.vram_rd_clk_det_1_LC_4_11_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_4_11_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_4_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9132),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__17779));
    defparam \uu0.l_precount_0_LC_4_12_3 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_4_12_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_4_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9085),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18030),
            .ce(),
            .sr(N__17827));
    defparam \buart.Z_rx.hh_1_LC_5_2_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_5_2_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_5_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18090),
            .ce(),
            .sr(N__17831));
    defparam \buart.Z_rx.hh_0_LC_5_3_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_5_3_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_5_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9055),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18083),
            .ce(),
            .sr(N__17829));
    defparam \uu2.r_addr_esr_8_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_5_4_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_esr_8_LC_5_4_1  (
            .in0(N__9382),
            .in1(N__9221),
            .in2(N__9016),
            .in3(N__9027),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18073),
            .ce(N__9466),
            .sr(N__17808));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__9519),
            .in2(_gnd_net_),
            .in3(N__9487),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_5_4_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_7_LC_5_4_3  (
            .in0(N__9405),
            .in1(N__9434),
            .in2(N__9535),
            .in3(N__9222),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18073),
            .ce(N__9466),
            .sr(N__17808));
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_5_4_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_esr_6_LC_5_4_5  (
            .in0(N__9520),
            .in1(N__9489),
            .in2(N__9226),
            .in3(N__9435),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18073),
            .ce(N__9466),
            .sr(N__17808));
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_5_4_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_5_4_6  (
            .in0(N__9376),
            .in1(N__9340),
            .in2(N__9294),
            .in3(N__9268),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18073),
            .ce(N__9466),
            .sr(N__17808));
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un426_ci_LC_5_4_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un426_ci_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un426_ci_LC_5_4_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.counter_gen_label_6__un426_ci_LC_5_4_7  (
            .in0(N__13830),
            .in1(N__13231),
            .in2(N__13753),
            .in3(N__13629),
            .lcout(\uu2.un426_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_5_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_5_5_2  (
            .in0(N__12337),
            .in1(N__10077),
            .in2(_gnd_net_),
            .in3(N__13318),
            .lcout(\uu2.mem0.N_70_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_5_3 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_5_5_3  (
            .in0(N__9430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9404),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_5_5 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_5_5_5  (
            .in0(N__9370),
            .in1(N__9335),
            .in2(N__9293),
            .in3(N__9263),
            .lcout(\uu2.un404_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_i_1_5_LC_5_5_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_i_1_5_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_i_1_5_LC_5_5_7 .LUT_INIT=16'b1110110110101100;
    LogicCell40 \Lab_UT.bcd2segment4.segment_i_1_5_LC_5_5_7  (
            .in0(N__17492),
            .in1(N__14944),
            .in2(N__15490),
            .in3(N__17252),
            .lcout(\Lab_UT.bcd2segment4.segment_i_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_0_2_LC_5_6_0 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \Lab_UT.bcd2segment4.segment_0_2_LC_5_6_0  (
            .in0(N__17488),
            .in1(N__14937),
            .in2(N__15511),
            .in3(N__17248),
            .lcout(\Lab_UT.bcd2segment4.segment_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIG4PV_66_LC_5_6_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIG4PV_66_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIG4PV_66_LC_5_6_1 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNIG4PV_66_LC_5_6_1  (
            .in0(N__9541),
            .in1(N__12881),
            .in2(N__9556),
            .in3(N__10821),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_20_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIKJFQ1_69_LC_5_6_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKJFQ1_69_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKJFQ1_69_LC_5_6_2 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.bitmap_RNIKJFQ1_69_LC_5_6_2  (
            .in0(N__12882),
            .in1(N__9577),
            .in2(N__9589),
            .in3(N__9568),
            .lcout(\uu2.N_40_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_197_LC_5_6_3 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_5_6_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.bitmap_197_LC_5_6_3  (
            .in0(N__14227),
            .in1(_gnd_net_),
            .in2(N__9586),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__17781));
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_0_1_LC_5_6_4 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \Lab_UT.bcd2segment4.segment_0_1_LC_5_6_4  (
            .in0(N__14941),
            .in1(N__17249),
            .in2(N__17494),
            .in3(N__14226),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment4.segment_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_69_LC_5_6_5 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_5_6_5 .LUT_INIT=16'b0111000010110000;
    LogicCell40 \uu2.bitmap_69_LC_5_6_5  (
            .in0(N__17251),
            .in1(N__15494),
            .in2(N__9571),
            .in3(N__14344),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__17781));
    defparam \uu2.bitmap_194_LC_5_6_6 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_5_6_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.bitmap_194_LC_5_6_6  (
            .in0(N__14239),
            .in1(N__17250),
            .in2(_gnd_net_),
            .in3(N__9562),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__17781));
    defparam \uu2.bitmap_66_LC_5_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_5_6_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_66_LC_5_6_7  (
            .in0(N__14228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9547),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__17781));
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_38_LC_5_7_0 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_38_LC_5_7_0  (
            .in0(N__13710),
            .in1(N__12974),
            .in2(_gnd_net_),
            .in3(N__13028),
            .lcout(\uu2.mem0.N_1201_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_53_LC_5_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_53_LC_5_7_1  (
            .in0(N__12840),
            .in1(N__12696),
            .in2(_gnd_net_),
            .in3(N__11114),
            .lcout(\uu2.mem0.g0_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep2_RNI1HJ81_LC_5_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep2_RNI1HJ81_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep2_RNI1HJ81_LC_5_7_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \uu2.w_addr_displaying_3_rep2_RNI1HJ81_LC_5_7_2  (
            .in0(N__13709),
            .in1(N__12973),
            .in2(N__12719),
            .in3(N__13030),
            .lcout(\uu2.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_7_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_37_LC_5_7_3 .LUT_INIT=16'b0100100011100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_37_LC_5_7_3  (
            .in0(N__13027),
            .in1(N__13711),
            .in2(N__12979),
            .in3(N__12700),
            .lcout(\uu2.mem0.bitmap_pmux_sn_N_20_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_59_LC_5_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_59_LC_5_7_4  (
            .in0(_gnd_net_),
            .in1(N__12839),
            .in2(_gnd_net_),
            .in3(N__11065),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_u_ns_1_N_2_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_41_LC_5_7_5 .LUT_INIT=16'b1001010010010010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_41_LC_5_7_5  (
            .in0(N__13029),
            .in1(N__13712),
            .in2(N__9643),
            .in3(N__12954),
            .lcout(\uu2.mem0.g1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI5R5D8_69_LC_5_7_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI5R5D8_69_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI5R5D8_69_LC_5_7_6 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \uu2.bitmap_RNI5R5D8_69_LC_5_7_6  (
            .in0(N__9694),
            .in1(N__9634),
            .in2(N__9628),
            .in3(N__10099),
            .lcout(\uu2.N_404 ),
            .ltout(\uu2.N_404_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_5_7_7 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_5_7_7  (
            .in0(N__9718),
            .in1(N__9613),
            .in2(N__9607),
            .in3(N__9682),
            .lcout(\uu2.mem0.bitmap_pmux_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_5_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_61_LC_5_8_0 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_61_LC_5_8_0  (
            .in0(N__13213),
            .in1(N__10804),
            .in2(N__13395),
            .in3(N__10762),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_46_LC_5_8_1 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_46_LC_5_8_1  (
            .in0(N__12738),
            .in1(N__12866),
            .in2(N__9598),
            .in3(N__11113),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_58_LC_5_8_2 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_58_LC_5_8_2  (
            .in0(N__13214),
            .in1(N__10805),
            .in2(N__13396),
            .in3(N__10763),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_N_42_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_3 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_40_LC_5_8_3  (
            .in0(N__12739),
            .in1(N__12955),
            .in2(N__9745),
            .in3(N__12865),
            .lcout(),
            .ltout(\uu2.mem0.g1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_24_LC_5_8_4  (
            .in0(N__9741),
            .in1(N__13141),
            .in2(N__9727),
            .in3(N__9724),
            .lcout(\uu2.mem0.bitmap_pmux_sn_i7_mux_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNIT4P31_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIT4P31_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIT4P31_LC_5_8_5 .LUT_INIT=16'b0010110010001000;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIT4P31_LC_5_8_5  (
            .in0(N__13737),
            .in1(N__11112),
            .in2(N__12742),
            .in3(N__11264),
            .lcout(\uu2.bitmap_pmux_sn_N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIVOBS1_93_LC_5_8_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIVOBS1_93_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIVOBS1_93_LC_5_8_6 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.bitmap_RNIVOBS1_93_LC_5_8_6  (
            .in0(N__12867),
            .in1(N__10111),
            .in2(N__13129),
            .in3(N__9703),
            .lcout(\uu2.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_5_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_23_LC_5_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_23_LC_5_8_7  (
            .in0(N__9688),
            .in1(N__9903),
            .in2(_gnd_net_),
            .in3(N__9649),
            .lcout(\uu2.mem0.N_2166_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNIKIVT_LC_5_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIKIVT_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIKIVT_LC_5_9_0 .LUT_INIT=16'b0000011100000110;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIKIVT_LC_5_9_0  (
            .in0(N__11256),
            .in1(N__11110),
            .in2(N__10814),
            .in3(N__11058),
            .lcout(\uu2.bitmap_pmux_sn_N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_5_9_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_62_LC_5_9_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_62_LC_5_9_1  (
            .in0(N__10143),
            .in1(N__9811),
            .in2(_gnd_net_),
            .in3(N__9798),
            .lcout(),
            .ltout(\uu2.mem0.N_247_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_9_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_56_LC_5_9_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_56_LC_5_9_2  (
            .in0(N__10799),
            .in1(N__11057),
            .in2(N__9676),
            .in3(N__9855),
            .lcout(),
            .ltout(\uu2.mem0.N_2171_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_36_LC_5_9_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_36_LC_5_9_3  (
            .in0(N__12741),
            .in1(N__9817),
            .in2(N__9673),
            .in3(N__9660),
            .lcout(\uu2.mem0.N_397_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_4 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_57_LC_5_9_4  (
            .in0(N__11257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10760),
            .lcout(\uu2.mem0.g1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI232M_52_LC_5_9_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI232M_52_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI232M_52_LC_5_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.bitmap_RNI232M_52_LC_5_9_5  (
            .in0(N__10142),
            .in1(N__9810),
            .in2(_gnd_net_),
            .in3(N__9799),
            .lcout(),
            .ltout(\uu2.N_247_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_rep1_nesr_RNI023T1_LC_5_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_nesr_RNI023T1_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_7_rep1_nesr_RNI023T1_LC_5_9_6 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_nesr_RNI023T1_LC_5_9_6  (
            .in0(N__10803),
            .in1(N__11059),
            .in2(N__9787),
            .in3(N__9856),
            .lcout(\uu2.N_2171_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_44_LC_5_9_7 .LUT_INIT=16'b0010001001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_44_LC_5_9_7  (
            .in0(N__11111),
            .in1(N__13738),
            .in2(_gnd_net_),
            .in3(N__11258),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.N_198_i_1_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.N_198_i_1_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.N_198_i_1_LC_5_10_0 .LUT_INIT=16'b0001010001000111;
    LogicCell40 \Lab_UT.bcd2segment4.N_198_i_1_LC_5_10_0  (
            .in0(N__17486),
            .in1(N__14935),
            .in2(N__15526),
            .in3(N__17253),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment4.N_198_iZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_290_LC_5_10_1 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_5_10_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_290_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9766),
            .in3(N__14235),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__17780));
    defparam \Lab_UT.bcd2segment4.segment_i_0_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_i_0_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_i_0_0_LC_5_10_2 .LUT_INIT=16'b0010100100010000;
    LogicCell40 \Lab_UT.bcd2segment4.segment_i_0_0_LC_5_10_2  (
            .in0(N__17487),
            .in1(N__14936),
            .in2(N__15527),
            .in3(N__17254),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment4.segment_i_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_34_LC_5_10_3 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_5_10_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_34_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9763),
            .in3(N__14236),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__17780));
    defparam \uu2.bitmap_RNI8LAO_34_LC_5_10_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI8LAO_34_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI8LAO_34_LC_5_10_4 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \uu2.bitmap_RNI8LAO_34_LC_5_10_4  (
            .in0(N__9760),
            .in1(N__10141),
            .in2(N__9754),
            .in3(N__10239),
            .lcout(\uu2.bitmap_pmux_15_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_3_LC_5_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_3_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_3_LC_5_10_5 .LUT_INIT=16'b1010101001011010;
    LogicCell40 \uu2.w_addr_displaying_fast_3_LC_5_10_5  (
            .in0(N__10241),
            .in1(_gnd_net_),
            .in2(N__12223),
            .in3(N__13804),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__17780));
    defparam \uu2.bitmap_RNILMVP_180_LC_5_10_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNILMVP_180_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNILMVP_180_LC_5_10_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.bitmap_RNILMVP_180_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(N__10240),
            .in2(N__9878),
            .in3(N__9847),
            .lcout(\uu2.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_180_LC_5_10_7 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_5_10_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_180_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__14234),
            .in2(_gnd_net_),
            .in3(N__11149),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__17780));
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_5_11_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_3_LC_5_11_0 .LUT_INIT=16'b1111100011100110;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_3_LC_5_11_0  (
            .in0(N__15730),
            .in1(N__15981),
            .in2(N__16080),
            .in3(N__15819),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segmentUQ_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_5_11_1 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_5_11_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_5_11_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_296_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9841),
            .in3(N__14232),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__17784));
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_5_11_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_0_0_LC_5_11_2 .LUT_INIT=16'b1101111101111001;
    LogicCell40 \Lab_UT.bcd2segment3.segment_0_0_LC_5_11_2  (
            .in0(N__15731),
            .in1(N__15982),
            .in2(N__16081),
            .in3(N__15820),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segment_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_5_11_3 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_5_11_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \uu2.bitmap_40_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9838),
            .in3(N__14233),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__17784));
    defparam \uu2.bitmap_RNI2S3H1_40_LC_5_11_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI2S3H1_40_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI2S3H1_40_LC_5_11_4 .LUT_INIT=16'b1100000010101111;
    LogicCell40 \uu2.bitmap_RNI2S3H1_40_LC_5_11_4  (
            .in0(N__9835),
            .in1(N__9829),
            .in2(N__11074),
            .in3(N__9823),
            .lcout(\uu2.N_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_5_11_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_5_11_5 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIF4D9_2_LC_5_11_5  (
            .in0(N__10048),
            .in1(N__10243),
            .in2(_gnd_net_),
            .in3(N__10198),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNITQGB1_111_LC_5_11_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNITQGB1_111_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNITQGB1_111_LC_5_11_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.bitmap_RNITQGB1_111_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(N__9934),
            .in2(N__9928),
            .in3(N__10213),
            .lcout(),
            .ltout(\uu2.N_395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNIJ9KQ3_LC_5_11_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIJ9KQ3_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIJ9KQ3_LC_5_11_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIJ9KQ3_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(N__9925),
            .in2(N__9916),
            .in3(N__9913),
            .lcout(\uu2.N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_5_LC_5_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_5_12_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_5_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_5_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18025),
            .ce(N__11713),
            .sr(N__17828));
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_5_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_5_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11347),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18025),
            .ce(N__11713),
            .sr(N__17828));
    defparam \buart.Z_rx.shifter_7_LC_5_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_5_12_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9979),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18025),
            .ce(N__11713),
            .sr(N__17828));
    defparam \buart.Z_rx.bitcount_RNI9OJJ_1_LC_6_2_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9OJJ_1_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9OJJ_1_LC_6_2_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9OJJ_1_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__10577),
            .in2(_gnd_net_),
            .in3(N__10356),
            .lcout(),
            .ltout(\buart.Z_rx.idle_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_6_2_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_4_LC_6_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_4_LC_6_2_2  (
            .in0(N__10482),
            .in1(N__10543),
            .in2(N__9886),
            .in3(N__11739),
            .lcout(\buart.Z_rx.idle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_6_2_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIAPJJ_1_LC_6_2_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIAPJJ_1_LC_6_2_3  (
            .in0(_gnd_net_),
            .in1(N__10481),
            .in2(_gnd_net_),
            .in3(N__10355),
            .lcout(),
            .ltout(\buart.Z_rx.valid_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_4_LC_6_2_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_4_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNI9F1H1_0_4_LC_6_2_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.bitcount_RNI9F1H1_0_4_LC_6_2_4  (
            .in0(N__10578),
            .in1(N__10542),
            .in2(N__9883),
            .in3(N__11738),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_6_2_7 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNI065O1_0_LC_6_2_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.hh_RNI065O1_0_LC_6_2_7  (
            .in0(N__9972),
            .in1(N__9961),
            .in2(_gnd_net_),
            .in3(N__11825),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_3_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11746),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_3_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__10357),
            .in2(_gnd_net_),
            .in3(N__9946),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_3_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__10579),
            .in2(_gnd_net_),
            .in3(N__9943),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_3_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__10484),
            .in2(_gnd_net_),
            .in3(N__9940),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_6_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_4_LC_6_3_4 .LUT_INIT=16'b0011010100111010;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_4_LC_6_3_4  (
            .in0(N__10545),
            .in1(N__11996),
            .in2(N__10510),
            .in3(N__9937),
            .lcout(\buart.Z_rx.bitcount_lm_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI8NF3_8_LC_6_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI8NF3_8_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI8NF3_8_LC_6_4_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.w_addr_user_nesr_RNI8NF3_8_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__10076),
            .in2(_gnd_net_),
            .in3(N__10008),
            .lcout(\uu2.N_153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_5_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_5_0  (
            .in0(N__12648),
            .in1(N__12544),
            .in2(N__10440),
            .in3(N__11911),
            .lcout(\uu2.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_6_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_6_5_1 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_6_LC_6_5_1  (
            .in0(N__11912),
            .in1(N__10435),
            .in2(N__12552),
            .in3(N__12649),
            .lcout(),
            .ltout(\uu2.N_150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_6_LC_6_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_6_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_6_LC_6_5_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uu2.w_addr_user_nesr_6_LC_6_5_2  (
            .in0(N__10022),
            .in1(N__12509),
            .in2(N__10084),
            .in3(N__12597),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_6C_net ),
            .ce(N__10621),
            .sr(N__17790));
    defparam \uu2.w_addr_user_nesr_8_LC_6_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_6_5_3 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_6_5_3  (
            .in0(N__12598),
            .in1(N__10023),
            .in2(N__10081),
            .in3(N__10007),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_6C_net ),
            .ce(N__10621),
            .sr(N__17790));
    defparam \uu2.w_addr_user_nesr_0_LC_6_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_0_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_0_LC_6_5_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \uu2.w_addr_user_nesr_0_LC_6_5_4  (
            .in0(N__10715),
            .in1(N__12548),
            .in2(N__12514),
            .in3(N__12596),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_6C_net ),
            .ce(N__10621),
            .sr(N__17790));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_5_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_6_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_6_5_6  (
            .in0(N__10714),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__12883),
            .lcout(\uu2.mem0.N_78_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_6_6_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_6_6_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_4_LC_6_6_0  (
            .in0(N__12196),
            .in1(N__13594),
            .in2(N__13840),
            .in3(N__13716),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_displaying_3_LC_6_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_LC_6_6_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uu2.w_addr_displaying_3_LC_6_6_1  (
            .in0(N__13593),
            .in1(N__13831),
            .in2(_gnd_net_),
            .in3(N__12194),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_displaying_3_rep2_LC_6_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep2_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep2_LC_6_6_2 .LUT_INIT=16'b1111010100001010;
    LogicCell40 \uu2.w_addr_displaying_3_rep2_LC_6_6_2  (
            .in0(N__12195),
            .in1(_gnd_net_),
            .in2(N__13839),
            .in3(N__12733),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_displaying_fast_2_LC_6_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_6_6_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_6_6_3  (
            .in0(N__13069),
            .in1(N__12884),
            .in2(N__10047),
            .in3(N__12197),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_user_1_LC_6_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_6_6_4 .LUT_INIT=16'b0001010011110000;
    LogicCell40 \uu2.w_addr_user_1_LC_6_6_4  (
            .in0(N__12586),
            .in1(N__10723),
            .in2(N__10685),
            .in3(N__12485),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_user_7_LC_6_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_7_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_7_LC_6_6_5 .LUT_INIT=16'b0111010100000010;
    LogicCell40 \uu2.w_addr_user_7_LC_6_6_5  (
            .in0(N__12487),
            .in1(N__12588),
            .in2(N__10027),
            .in3(N__10006),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.w_addr_user_4_LC_6_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_6_6_6 .LUT_INIT=16'b0100000111110000;
    LogicCell40 \uu2.w_addr_user_4_LC_6_6_6  (
            .in0(N__12587),
            .in1(N__10439),
            .in2(N__12659),
            .in3(N__12486),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.bitmap_221_LC_6_6_7 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_6_6_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_6_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.bitmap_221_LC_6_6_7  (
            .in0(N__10123),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14240),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_4C_net ),
            .ce(),
            .sr(N__17786));
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_6_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_48_LC_6_7_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_48_LC_6_7_0  (
            .in0(N__13682),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11115),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_7_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_55_LC_6_7_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_55_LC_6_7_1  (
            .in0(N__12716),
            .in1(N__12945),
            .in2(N__13506),
            .in3(N__13384),
            .lcout(),
            .ltout(\uu2.mem0.g0_7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_7_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_35_LC_6_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_35_LC_6_7_2  (
            .in0(N__13683),
            .in1(N__10923),
            .in2(N__10102),
            .in3(N__13230),
            .lcout(\uu2.mem0.un49_w_data_displaying_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_RNI5QH04_LC_6_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_RNI5QH04_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_RNI5QH04_LC_6_7_3 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_RNI5QH04_LC_6_7_3  (
            .in0(N__12718),
            .in1(N__11066),
            .in2(N__11218),
            .in3(N__10279),
            .lcout(\uu2.bitmap_pmux_27_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_6_7_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_54_LC_6_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_54_LC_6_7_4  (
            .in0(N__13681),
            .in1(N__13494),
            .in2(N__13402),
            .in3(N__13229),
            .lcout(),
            .ltout(\uu2.mem0.g0_6_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_7_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_34_LC_6_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_34_LC_6_7_5  (
            .in0(N__10093),
            .in1(N__13306),
            .in2(N__10087),
            .in3(N__13052),
            .lcout(\uu2.mem0.un31_w_data_displaying_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNIFG6E_LC_6_7_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIFG6E_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIFG6E_LC_6_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIFG6E_LC_6_7_6  (
            .in0(N__13680),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11262),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_6_7_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_47_LC_6_7_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_47_LC_6_7_7  (
            .in0(N__12717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12868),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_LC_6_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_rep1_LC_6_8_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_LC_6_8_0  (
            .in0(N__12220),
            .in1(N__12879),
            .in2(N__13072),
            .in3(N__11116),
            .lcout(\uu2.w_addr_displaying_2_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_1_LC_6_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_6_8_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_displaying_1_LC_6_8_1  (
            .in0(N__12876),
            .in1(_gnd_net_),
            .in2(N__12221),
            .in3(N__13064),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_6_LC_6_8_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_6_LC_6_8_2 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_6_LC_6_8_2 .LUT_INIT=16'b1011111111001000;
    LogicCell40 \uu2.w_addr_displaying_6_LC_6_8_2  (
            .in0(N__12250),
            .in1(N__12215),
            .in2(N__10159),
            .in3(N__13394),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_2_LC_6_8_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_6_8_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_2_LC_6_8_3  (
            .in0(N__12878),
            .in1(N__13065),
            .in2(N__12972),
            .in3(N__12219),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_0_LC_6_8_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_6_8_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__12206),
            .in2(_gnd_net_),
            .in3(N__12875),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_fast_1_LC_6_8_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_1_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_1_LC_6_8_5 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_displaying_fast_1_LC_6_8_5  (
            .in0(N__12880),
            .in1(_gnd_net_),
            .in2(N__12222),
            .in3(N__10197),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_1_rep1_LC_6_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_LC_6_8_6 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_LC_6_8_6  (
            .in0(N__11265),
            .in1(N__12877),
            .in2(_gnd_net_),
            .in3(N__12210),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_3_rep1_LC_6_8_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_LC_6_8_7 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_LC_6_8_7  (
            .in0(N__12211),
            .in1(N__13824),
            .in2(_gnd_net_),
            .in3(N__11067),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2_rep1C_net ),
            .ce(),
            .sr(N__17777));
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_6_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_8_LC_6_9_1 .LUT_INIT=16'b1111101100000100;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_8_LC_6_9_1  (
            .in0(N__13802),
            .in1(N__13624),
            .in2(N__10885),
            .in3(N__10144),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .ce(N__13533),
            .sr(N__17782));
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_6_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI50L01_2_LC_6_9_2 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uu2.w_addr_displaying_RNI50L01_2_LC_6_9_2  (
            .in0(N__12969),
            .in1(N__13050),
            .in2(_gnd_net_),
            .in3(N__12864),
            .lcout(\uu2.N_46 ),
            .ltout(\uu2.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_6_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_6_9_3 .LUT_INIT=16'b1010101010100110;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_7_LC_6_9_3  (
            .in0(N__11205),
            .in1(N__13623),
            .in2(N__10201),
            .in3(N__13109),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .ce(N__13533),
            .sr(N__17782));
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_6_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_rep1_nesr_LC_6_9_4 .LUT_INIT=16'b1010101010011010;
    LogicCell40 \uu2.w_addr_displaying_8_rep1_nesr_LC_6_9_4  (
            .in0(N__10759),
            .in1(N__10880),
            .in2(N__13630),
            .in3(N__13801),
            .lcout(\uu2.w_addr_displaying_8_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .ce(N__13533),
            .sr(N__17782));
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_7_LC_6_9_5 .LUT_INIT=16'b1111000010110100;
    LogicCell40 \uu2.w_addr_displaying_nesr_7_LC_6_9_5  (
            .in0(N__13803),
            .in1(N__13625),
            .in2(N__13498),
            .in3(N__13110),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .ce(N__13533),
            .sr(N__17782));
    defparam \uu2.w_addr_displaying_7_rep1_nesr_LC_6_9_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_rep1_nesr_LC_6_9_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_rep1_nesr_LC_6_9_6 .LUT_INIT=16'b1111110100000010;
    LogicCell40 \uu2.w_addr_displaying_7_rep1_nesr_LC_6_9_6  (
            .in0(N__13619),
            .in1(N__13800),
            .in2(N__13111),
            .in3(N__10813),
            .lcout(\uu2.w_addr_displaying_7_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_nesr_8C_net ),
            .ce(N__13533),
            .sr(N__17782));
    defparam \uu2.w_addr_displaying_fast_RNIETIP_1_LC_6_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIETIP_1_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIETIP_1_LC_6_9_7 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIETIP_1_LC_6_9_7  (
            .in0(N__11064),
            .in1(N__10196),
            .in2(_gnd_net_),
            .in3(N__10758),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_4_LC_6_10_0 .LUT_INIT=16'b1111111011110010;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_4_LC_6_10_0  (
            .in0(N__15983),
            .in1(N__15821),
            .in2(N__15738),
            .in3(N__16078),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segmentUQ_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_200_LC_6_10_1 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_6_10_1 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_200_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10162),
            .in3(N__14223),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_200C_net ),
            .ce(),
            .sr(N__17785));
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_5_LC_6_10_2 .LUT_INIT=16'b1110111011010100;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_5_LC_6_10_2  (
            .in0(N__15984),
            .in1(N__15822),
            .in2(N__15739),
            .in3(N__16079),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segmentUQ_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_72_LC_6_10_3 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_6_10_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_72_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10285),
            .in3(N__14225),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_200C_net ),
            .ce(),
            .sr(N__17785));
    defparam \uu2.bitmap_RNI011L_75_LC_6_10_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI011L_75_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI011L_75_LC_6_10_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNI011L_75_LC_6_10_4  (
            .in0(N__10315),
            .in1(N__11201),
            .in2(_gnd_net_),
            .in3(N__10252),
            .lcout(),
            .ltout(\uu2.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNI588O1_LC_6_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNI588O1_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNI588O1_LC_6_10_5 .LUT_INIT=16'b0000100000011001;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNI588O1_LC_6_10_5  (
            .in0(N__12888),
            .in1(N__11266),
            .in2(N__10282),
            .in3(N__10258),
            .lcout(\uu2.g0_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIQQ0L_72_LC_6_10_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIQQ0L_72_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIQQ0L_72_LC_6_10_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNIQQ0L_72_LC_6_10_6  (
            .in0(N__10270),
            .in1(N__10264),
            .in2(_gnd_net_),
            .in3(N__11200),
            .lcout(\uu2.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_203_LC_6_10_7 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_6_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.bitmap_203_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(N__10303),
            .in2(_gnd_net_),
            .in3(N__14224),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_200C_net ),
            .ce(),
            .sr(N__17785));
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segmentUQ_6_LC_6_11_0 .LUT_INIT=16'b1110100111100001;
    LogicCell40 \Lab_UT.bcd2segment3.segmentUQ_6_LC_6_11_0  (
            .in0(N__15980),
            .in1(N__15818),
            .in2(N__16071),
            .in3(N__15729),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segmentUQ_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_168_LC_6_11_1 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_6_11_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \uu2.bitmap_168_LC_6_11_1  (
            .in0(N__14217),
            .in1(_gnd_net_),
            .in2(N__10246),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__17789));
    defparam \uu2.bitmap_RNISSSN_162_LC_6_11_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNISSSN_162_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNISSSN_162_LC_6_11_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNISSSN_162_LC_6_11_2  (
            .in0(N__10207),
            .in1(N__10242),
            .in2(_gnd_net_),
            .in3(N__10219),
            .lcout(\uu2.bitmap_RNISSSNZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_6_11_3 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_6_11_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uu2.bitmap_162_LC_6_11_3  (
            .in0(N__14216),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11287),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__17789));
    defparam \Lab_UT.bcd2segment3.segment_i_1_1_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_i_1_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_i_1_1_LC_6_11_4 .LUT_INIT=16'b0000001011111111;
    LogicCell40 \Lab_UT.bcd2segment3.segment_i_1_1_LC_6_11_4  (
            .in0(N__15979),
            .in1(N__15898),
            .in2(N__16070),
            .in3(N__14215),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment3.segment_i_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_6_11_5 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_6_11_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \uu2.bitmap_75_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10318),
            .in3(N__10309),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__17789));
    defparam \Lab_UT.bcd2segment3.segment_i_0_1_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_i_0_1_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_i_0_1_LC_6_11_6 .LUT_INIT=16'b1100000010101000;
    LogicCell40 \Lab_UT.bcd2segment3.segment_i_0_1_LC_6_11_6  (
            .in0(N__15977),
            .in1(N__15814),
            .in2(N__16069),
            .in3(N__15728),
            .lcout(\Lab_UT.bcd2segment3.segment_i_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.segment_i_0_2_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.segment_i_0_2_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.segment_i_0_2_LC_6_11_7 .LUT_INIT=16'b1100010000010000;
    LogicCell40 \Lab_UT.bcd2segment3.segment_i_0_2_LC_6_11_7  (
            .in0(N__15727),
            .in1(N__16049),
            .in2(N__15823),
            .in3(N__15978),
            .lcout(\Lab_UT.bcd2segment3.segment_i_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_1_0_LC_6_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_1_0_LC_6_12_0  (
            .in0(N__11461),
            .in1(N__11493),
            .in2(N__11398),
            .in3(N__13980),
            .lcout(\Lab_UT.dictrl.next_alarmstate4_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_3_LC_6_12_1 .C_ON=1'b0;
    defparam \resetGen.escKey_3_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_3_LC_6_12_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \resetGen.escKey_3_LC_6_12_1  (
            .in0(N__13981),
            .in1(N__11394),
            .in2(N__11500),
            .in3(N__11462),
            .lcout(\resetGen.escKeyZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state16_4_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state16_4_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state16_4_LC_6_12_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state16_4_LC_6_12_2  (
            .in0(N__11460),
            .in1(N__11492),
            .in2(N__11397),
            .in3(N__13979),
            .lcout(\Lab_UT.dictrl.next_state16Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_6_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_6_12_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_6_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_LC_6_12_3  (
            .in0(N__11497),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18021),
            .ce(N__11712),
            .sr(N__17830));
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_2_0_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_2_0_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_2_0_LC_6_12_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_sqmuxa_2_0_LC_6_12_4  (
            .in0(N__11459),
            .in1(N__11491),
            .in2(N__11531),
            .in3(N__13978),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxa_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_6_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_6_12_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_6_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_6_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18021),
            .ce(N__11712),
            .sr(N__17830));
    defparam \buart.Z_rx.shifter_4_LC_6_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_6_12_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_6_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_4_LC_6_12_6  (
            .in0(N__11524),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18021),
            .ce(N__11712),
            .sr(N__17830));
    defparam \buart.Z_rx.shifter_3_LC_6_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_6_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_6_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11463),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18021),
            .ce(N__11712),
            .sr(N__17830));
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_7_2_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIMK771_4_LC_7_2_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_RNIMK771_4_LC_7_2_4  (
            .in0(N__10580),
            .in1(N__10483),
            .in2(N__10360),
            .in3(N__10544),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIIU223_4_LC_7_2_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIIU223_4_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIIU223_4_LC_7_2_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_rx.bitcount_RNIIU223_4_LC_7_2_5  (
            .in0(_gnd_net_),
            .in1(N__11826),
            .in2(_gnd_net_),
            .in3(N__11795),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(\buart.Z_rx.N_27_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_7_2_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_0_LC_7_2_6 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_0_LC_7_2_6  (
            .in0(N__11997),
            .in1(N__10412),
            .in2(N__10378),
            .in3(N__11743),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_0_LC_7_2_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_0_LC_7_2_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_0_LC_7_2_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_0_LC_7_2_7  (
            .in0(N__11744),
            .in1(N__11772),
            .in2(N__10375),
            .in3(N__11998),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18091),
            .ce(),
            .sr(N__17834));
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_7_3_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_1_LC_7_3_0 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_1_LC_7_3_0  (
            .in0(N__11999),
            .in1(N__10358),
            .in2(N__10372),
            .in3(N__10507),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_1_LC_7_3_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_1_LC_7_3_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_1_LC_7_3_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_1_LC_7_3_1  (
            .in0(N__10359),
            .in1(N__11773),
            .in2(N__10363),
            .in3(N__12002),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18084),
            .ce(),
            .sr(N__17833));
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_7_3_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_2_LC_7_3_2 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_2_LC_7_3_2  (
            .in0(N__12000),
            .in1(N__10581),
            .in2(N__10327),
            .in3(N__10508),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_2_LC_7_3_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_2_LC_7_3_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_2_LC_7_3_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_2_LC_7_3_3  (
            .in0(N__10582),
            .in1(N__11774),
            .in2(N__10585),
            .in3(N__12003),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18084),
            .ce(),
            .sr(N__17833));
    defparam \buart.Z_rx.bitcount_4_LC_7_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_4_LC_7_3_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_4_LC_7_3_4 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \buart.Z_rx.bitcount_4_LC_7_3_4  (
            .in0(N__12005),
            .in1(N__10546),
            .in2(N__11779),
            .in3(N__10552),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18084),
            .ce(),
            .sr(N__17833));
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_7_3_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNO_0_3_LC_7_3_6 .LUT_INIT=16'b0101010100111100;
    LogicCell40 \buart.Z_rx.bitcount_RNO_0_3_LC_7_3_6  (
            .in0(N__12001),
            .in1(N__10485),
            .in2(N__10519),
            .in3(N__10509),
            .lcout(),
            .ltout(\buart.Z_rx.bitcount_lm_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_3_LC_7_3_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_3_LC_7_3_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_3_LC_7_3_7 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \buart.Z_rx.bitcount_3_LC_7_3_7  (
            .in0(N__10486),
            .in1(N__11775),
            .in2(N__10489),
            .in3(N__12004),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18084),
            .ce(),
            .sr(N__17833));
    defparam \uu2.w_addr_user_RNIPJCC_1_LC_7_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIPJCC_1_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIPJCC_1_LC_7_4_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu2.w_addr_user_RNIPJCC_1_LC_7_4_6  (
            .in0(N__10716),
            .in1(N__11854),
            .in2(N__10687),
            .in3(N__10456),
            .lcout(\uu2.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_7_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_7_5_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIFBD5_3_LC_7_5_3  (
            .in0(N__10717),
            .in1(N__11936),
            .in2(N__10682),
            .in3(N__11878),
            .lcout(\uu2.N_90 ),
            .ltout(\uu2.N_90_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_7_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_7_5_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_7_5_4  (
            .in0(N__12581),
            .in1(_gnd_net_),
            .in2(N__10450),
            .in3(N__10447),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__10617),
            .sr(N__17792));
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_7_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_7_5_5 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_3_LC_7_5_5  (
            .in0(N__10718),
            .in1(N__11937),
            .in2(N__10683),
            .in3(N__11879),
            .lcout(\uu2.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_5_LC_7_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_5_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_5_LC_7_5_6 .LUT_INIT=16'b0100000101000100;
    LogicCell40 \uu2.w_addr_user_nesr_5_LC_7_5_6  (
            .in0(N__12582),
            .in1(N__11913),
            .in2(N__10441),
            .in3(N__12653),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__10617),
            .sr(N__17792));
    defparam \uu2.w_addr_user_nesr_2_LC_7_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_2_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_2_LC_7_5_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu2.w_addr_user_nesr_2_LC_7_5_7  (
            .in0(N__10719),
            .in1(N__11880),
            .in2(N__10684),
            .in3(N__12580),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__10617),
            .sr(N__17792));
    defparam \Lab_UT.dictrl.state_ret_4_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_4_LC_7_6_0 .LUT_INIT=16'b1111101110101011;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_LC_7_6_0  (
            .in0(N__17644),
            .in1(N__11635),
            .in2(N__11650),
            .in3(N__11602),
            .lcout(\Lab_UT.dictrl.state_retZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18062),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_1 .LUT_INIT=16'b1011101111010101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_1  (
            .in0(N__15171),
            .in1(N__15243),
            .in2(N__16255),
            .in3(N__15381),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_7_6_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_18_LC_7_6_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_18_LC_7_6_2  (
            .in0(N__14987),
            .in1(N__12459),
            .in2(_gnd_net_),
            .in3(N__12366),
            .lcout(\uu2.mem0.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI34K17_8_LC_7_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI34K17_8_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI34K17_8_LC_7_6_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI34K17_8_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__17642),
            .in2(_gnd_net_),
            .in3(N__12163),
            .lcout(\uu2.un21_w_addr_displaying_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIB4K34_6_LC_7_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIB4K34_6_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIB4K34_6_LC_7_6_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uu2.w_addr_user_nesr_RNIB4K34_6_LC_7_6_4  (
            .in0(N__17643),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12477),
            .lcout(\uu2.un28_w_addr_user_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_6_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_7_6_5  (
            .in0(N__11910),
            .in1(N__12282),
            .in2(_gnd_net_),
            .in3(N__13225),
            .lcout(\uu2.mem0.N_73_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_7_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dispString.rdy_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15316),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18062),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_7_7_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_32_LC_7_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_32_LC_7_7_0  (
            .in0(N__13376),
            .in1(N__12946),
            .in2(N__13504),
            .in3(N__13707),
            .lcout(\uu2.mem0.g0_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_8_LC_7_7_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_8_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_8_LC_7_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI25P31_0_8_LC_7_7_1  (
            .in0(N__13032),
            .in1(N__13280),
            .in2(_gnd_net_),
            .in3(N__12859),
            .lcout(\uu2.un49_w_data_displaying_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_8_LC_7_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_8_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_8_LC_7_7_2 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI25P31_8_LC_7_7_2  (
            .in0(N__12860),
            .in1(_gnd_net_),
            .in2(N__13304),
            .in3(N__13031),
            .lcout(),
            .ltout(\uu2.un31_w_data_displaying_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIFOBB3_2_LC_7_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIFOBB3_2_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIFOBB3_2_LC_7_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIFOBB3_2_LC_7_7_3  (
            .in0(N__12947),
            .in1(N__13577),
            .in2(N__10960),
            .in3(N__10933),
            .lcout(\uu2.un31_w_data_displaying ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_7_LC_7_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_7_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_7_LC_7_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNISQPH1_7_LC_7_7_4  (
            .in0(N__13374),
            .in1(N__13200),
            .in2(N__13503),
            .in3(N__13706),
            .lcout(\uu2.un15_w_data_displaying_6 ),
            .ltout(\uu2.un15_w_data_displaying_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIFOBB3_0_2_LC_7_7_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIFOBB3_0_2_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIFOBB3_0_2_LC_7_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIFOBB3_0_2_LC_7_7_5  (
            .in0(N__12948),
            .in1(N__13578),
            .in2(N__10927),
            .in3(N__10924),
            .lcout(\uu2.un49_w_data_displaying ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_0_7_LC_7_7_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_0_7_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNISQPH1_0_7_LC_7_7_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNISQPH1_0_7_LC_7_7_6  (
            .in0(N__13375),
            .in1(N__13201),
            .in2(N__13505),
            .in3(N__13708),
            .lcout(\uu2.un15_w_data_displaying_i_i_o2_0 ),
            .ltout(\uu2.un15_w_data_displaying_i_i_o2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_7_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_8_LC_7_7_7 .LUT_INIT=16'b1010101010100110;
    LogicCell40 \uu2.w_addr_displaying_nesr_8_LC_7_7_7  (
            .in0(N__13303),
            .in1(N__13579),
            .in2(N__10861),
            .in3(N__13828),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_8C_net ),
            .ce(N__13523),
            .sr(N__17787));
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_7_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_20_LC_7_8_0 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_20_LC_7_8_0  (
            .in0(N__10858),
            .in1(N__10969),
            .in2(N__10852),
            .in3(N__10840),
            .lcout(\uu2.mem0.g1_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_60_LC_7_8_1 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_60_LC_7_8_1  (
            .in0(N__13373),
            .in1(N__10806),
            .in2(_gnd_net_),
            .in3(N__10761),
            .lcout(),
            .ltout(\uu2.mem0.bitmap_pmux_sn_N_57_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_45_LC_7_8_2 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_45_LC_7_8_2  (
            .in0(N__13216),
            .in1(N__11006),
            .in2(N__11128),
            .in3(N__11017),
            .lcout(\uu2.mem0.ram512X8_inst_RNOZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_rep1_RNIDKIL_LC_7_8_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_rep1_RNIDKIL_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_2_rep1_RNIDKIL_LC_7_8_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_2_rep1_RNIDKIL_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__11109),
            .in2(_gnd_net_),
            .in3(N__11063),
            .lcout(\uu2.bitmap_pmux_sn_N_31_0 ),
            .ltout(\uu2.bitmap_pmux_sn_N_31_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_49_LC_7_8_4 .LUT_INIT=16'b0110011001100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_49_LC_7_8_4  (
            .in0(N__13464),
            .in1(N__13290),
            .in2(N__11011),
            .in3(N__11007),
            .lcout(),
            .ltout(\uu2.mem0.ram512X8_inst_RNOZ0Z_49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_28_LC_7_8_5 .LUT_INIT=16'b0101000000100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_28_LC_7_8_5  (
            .in0(N__11008),
            .in1(N__10996),
            .in2(N__10990),
            .in3(N__10987),
            .lcout(\uu2.mem0.bitmap_pmux_u_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_8_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_52_LC_7_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_52_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(N__12734),
            .in2(_gnd_net_),
            .in3(N__13215),
            .lcout(),
            .ltout(\uu2.mem0.g0_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_33_LC_7_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_33_LC_7_8_7  (
            .in0(N__13289),
            .in1(N__13051),
            .in2(N__10972),
            .in3(N__12874),
            .lcout(\uu2.mem0.g0_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_i_0_1_LC_7_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_i_0_1_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_i_0_1_LC_7_9_0 .LUT_INIT=16'b1011001010000000;
    LogicCell40 \Lab_UT.bcd2segment2.segment_i_0_1_LC_7_9_0  (
            .in0(N__17548),
            .in1(N__16243),
            .in2(N__16319),
            .in3(N__16155),
            .lcout(\Lab_UT.bcd2segment2.segment_i_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_i_0_2_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_i_0_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_i_0_2_LC_7_9_1 .LUT_INIT=16'b1000101000000100;
    LogicCell40 \Lab_UT.bcd2segment2.segment_i_0_2_LC_7_9_1  (
            .in0(N__16156),
            .in1(N__16308),
            .in2(N__16251),
            .in3(N__17549),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment2.segment_i_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_7_9_2 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_7_9_2 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \uu2.bitmap_215_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10963),
            .in3(N__14209),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__17788));
    defparam \uu2.bitmap_RNI693L_87_LC_7_9_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI693L_87_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI693L_87_LC_7_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNI693L_87_LC_7_9_3  (
            .in0(N__13864),
            .in1(N__11199),
            .in2(_gnd_net_),
            .in3(N__11272),
            .lcout(),
            .ltout(\uu2.N_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_RNIHOCO1_LC_7_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_RNIHOCO1_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_RNIHOCO1_LC_7_9_4 .LUT_INIT=16'b0110111001111111;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_RNIHOCO1_LC_7_9_4  (
            .in0(N__12852),
            .in1(N__11263),
            .in2(N__11221),
            .in3(N__11173),
            .lcout(\uu2.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI033L_84_LC_7_9_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI033L_84_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI033L_84_LC_7_9_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.bitmap_RNI033L_84_LC_7_9_5  (
            .in0(N__11161),
            .in1(N__11167),
            .in2(_gnd_net_),
            .in3(N__11198),
            .lcout(\uu2.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_84_LC_7_9_6 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_7_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.bitmap_84_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(N__14210),
            .in2(_gnd_net_),
            .in3(N__11155),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__17788));
    defparam \uu2.bitmap_212_LC_7_9_7 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_7_9_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu2.bitmap_212_LC_7_9_7  (
            .in0(N__14211),
            .in1(N__11302),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__17788));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_1_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_1_LC_7_10_0 .LUT_INIT=16'b0000001101001101;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_1_1_LC_7_10_0  (
            .in0(N__16223),
            .in1(N__16145),
            .in2(N__16311),
            .in3(N__17546),
            .lcout(\Lab_UT.didp.countrce2.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_0_1_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_0_1_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_0_1_LC_7_10_1 .LUT_INIT=16'b0001011001010110;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_0_1_LC_7_10_1  (
            .in0(N__17544),
            .in1(N__16291),
            .in2(N__16163),
            .in3(N__16222),
            .lcout(\Lab_UT.didp.countrce2.N_175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_1_LC_7_10_2 .LUT_INIT=16'b0010100000000110;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_1_LC_7_10_2  (
            .in0(N__16221),
            .in1(N__16138),
            .in2(N__16310),
            .in3(N__17543),
            .lcout(\Lab_UT.didp.countrce2.N_170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.un1_num_7_1_0_a2_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.un1_num_7_1_0_a2_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.un1_num_7_1_0_a2_LC_7_10_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.bcd2segment4.un1_num_7_1_0_a2_LC_7_10_3  (
            .in0(N__14882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17452),
            .lcout(\Lab_UT.N_68_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_2_1_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_2_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_2_1_LC_7_10_4 .LUT_INIT=16'b0000000101111001;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_2_1_LC_7_10_4  (
            .in0(N__16220),
            .in1(N__16137),
            .in2(N__16309),
            .in3(N__17542),
            .lcout(\Lab_UT.didp.countrce2.N_183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_1_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_1_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_1_LC_7_10_5 .LUT_INIT=16'b0000000001000111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_1_LC_7_10_5  (
            .in0(N__17545),
            .in1(N__16292),
            .in2(N__16164),
            .in3(N__16224),
            .lcout(\Lab_UT.didp.countrce2.N_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_10_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_7_10_6  (
            .in0(N__17453),
            .in1(N__11293),
            .in2(N__17341),
            .in3(N__17285),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18037),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_7_10_7 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_7_10_7  (
            .in0(N__16348),
            .in1(N__16296),
            .in2(N__15859),
            .in3(N__16225),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18037),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_11_0 .LUT_INIT=16'b1001010101010101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_11_0  (
            .in0(N__17473),
            .in1(N__14916),
            .in2(N__15529),
            .in3(N__17221),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.N_80_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_11_1 .LUT_INIT=16'b1010111100000101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_11_1  (
            .in0(N__17363),
            .in1(_gnd_net_),
            .in2(N__11296),
            .in3(N__11396),
            .lcout(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.segment_i_0_6_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.segment_i_0_6_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.segment_i_0_6_LC_7_11_2 .LUT_INIT=16'b1110100110101001;
    LogicCell40 \Lab_UT.bcd2segment4.segment_i_0_6_LC_7_11_2  (
            .in0(N__17472),
            .in1(N__14915),
            .in2(N__15528),
            .in3(N__17220),
            .lcout(\Lab_UT.bcd2segment4.segment_i_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_0_LC_7_11_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_0_LC_7_11_3  (
            .in0(N__11533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11361),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_alarmstate4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate4_LC_7_11_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate4_LC_7_11_4  (
            .in0(N__11431),
            .in1(N__11281),
            .in2(N__11275),
            .in3(N__17386),
            .lcout(\Lab_UT.next_alarmstate4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_11_5 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_11_5  (
            .in0(N__17362),
            .in1(N__14350),
            .in2(_gnd_net_),
            .in3(N__11499),
            .lcout(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state16_5_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state16_5_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state16_5_LC_7_11_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.next_state16_5_LC_7_11_6  (
            .in0(N__11430),
            .in1(N__11532),
            .in2(N__11362),
            .in3(N__17385),
            .lcout(resetGen_escKey_4),
            .ltout(resetGen_escKey_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_11_7 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIBITA2_2_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__14604),
            .in2(N__11536),
            .in3(N__14034),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_2_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_2_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_2_LC_7_12_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_sqmuxa_2_LC_7_12_0  (
            .in0(N__11530),
            .in1(N__11498),
            .in2(N__11429),
            .in3(N__13982),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_7_12_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_sqmuxa_4_LC_7_12_1  (
            .in0(N__11387),
            .in1(N__11437),
            .in2(N__11467),
            .in3(N__11464),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_0_sqmuxaZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNI0C5J6_2_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNI0C5J6_2_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNI0C5J6_2_LC_7_12_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNI0C5J6_2_LC_7_12_2  (
            .in0(N__14125),
            .in1(N__11590),
            .in2(N__11440),
            .in3(N__13884),
            .lcout(\Lab_UT.dictrl.next_state_set ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_2_0_LC_7_12_3 .C_ON=1'b0;
    defparam \resetGen.escKey_2_0_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_2_0_LC_7_12_3 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \resetGen.escKey_2_0_LC_7_12_3  (
            .in0(N__17388),
            .in1(N__11351),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(resetGen_escKey_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_3_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_3_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_sqmuxa_3_LC_7_12_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_sqmuxa_3_LC_7_12_4  (
            .in0(N__11419),
            .in1(N__11386),
            .in2(N__11357),
            .in3(N__17387),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_1_sqmuxaZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_RNICD593_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_RNICD593_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_RNICD593_LC_7_12_5 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_RNICD593_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__11323),
            .in2(N__11317),
            .in3(N__14124),
            .lcout(\Lab_UT.dictrl.next_state_1_sqmuxa ),
            .ltout(\Lab_UT.dictrl.next_state_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNI1GK36_2_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNI1GK36_2_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNI1GK36_2_LC_7_12_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \Lab_UT.dictrl.state_0_RNI1GK36_2_LC_7_12_6  (
            .in0(N__11586),
            .in1(_gnd_net_),
            .in2(N__11575),
            .in3(N__11559),
            .lcout(\Lab_UT.dictrl.next_state_set_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_7_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_7_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_7_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_LC_7_12_7  (
            .in0(N__13983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18026),
            .ce(N__11705),
            .sr(N__17832));
    defparam \Lab_UT.dictrl.next_state_RNIN0UD1_2_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIN0UD1_2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIN0UD1_2_LC_7_13_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIN0UD1_2_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__14260),
            .in2(_gnd_net_),
            .in3(N__11569),
            .lcout(\Lab_UT.dictrl.next_state_RNIN0UD1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m37_ns_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.m37_ns_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m37_ns_LC_7_13_1 .LUT_INIT=16'b0010001100000011;
    LogicCell40 \Lab_UT.didp.m37_ns_LC_7_13_1  (
            .in0(N__17073),
            .in1(N__14641),
            .in2(N__14603),
            .in3(N__17008),
            .lcout(\Lab_UT.m37_ns ),
            .ltout(\Lab_UT.m37_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_2_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_7_13_2 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_2_LC_7_13_2 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_7_13_2  (
            .in0(N__14492),
            .in1(N__14282),
            .in2(N__11572),
            .in3(N__14308),
            .lcout(\Lab_UT.dictrl.next_state_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18022),
            .ce(N__14389),
            .sr(N__11563));
    defparam \Lab_UT.didp.m45_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.m45_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m45_LC_7_13_3 .LUT_INIT=16'b0000100011000000;
    LogicCell40 \Lab_UT.didp.m45_LC_7_13_3  (
            .in0(N__17072),
            .in1(N__17009),
            .in2(N__14602),
            .in3(N__16786),
            .lcout(\Lab_UT.m45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m40_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.m40_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m40_LC_7_13_4 .LUT_INIT=16'b0111000001100000;
    LogicCell40 \Lab_UT.didp.m40_LC_7_13_4  (
            .in0(N__16785),
            .in1(N__14587),
            .in2(N__17018),
            .in3(N__17074),
            .lcout(\Lab_UT.m40 ),
            .ltout(\Lab_UT.m40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI970U_3_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI970U_3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI970U_3_LC_7_13_5 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI970U_3_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__13912),
            .in2(N__11542),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3 ),
            .ltout(\Lab_UT.dictrl.next_state_RNI970UZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNISML65_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNISML65_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNISML65_LC_7_13_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNISML65_LC_7_13_6  (
            .in0(N__16863),
            .in1(N__15622),
            .in2(N__11539),
            .in3(N__15569),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m34_ns_1_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.m34_ns_1_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m34_ns_1_LC_7_13_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.didp.m34_ns_1_LC_7_13_7  (
            .in0(N__17071),
            .in1(N__17004),
            .in2(_gnd_net_),
            .in3(N__16784),
            .lcout(\Lab_UT.didp.m34_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNI919D9_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNI919D9_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNI919D9_LC_7_14_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNI919D9_LC_7_14_0  (
            .in0(N__16961),
            .in1(N__16941),
            .in2(N__16911),
            .in3(N__16805),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_0 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNI4EJF21_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNI4EJF21_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNI4EJF21_LC_7_14_1 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNI4EJF21_LC_7_14_1  (
            .in0(N__11625),
            .in1(N__14085),
            .in2(N__11638),
            .in3(N__14073),
            .lcout(\Lab_UT.dictrl.un1_state_21_reti_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_7_14_2 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_0_LC_7_14_2 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_7_14_2  (
            .in0(N__16962),
            .in1(N__16942),
            .in2(N__14497),
            .in3(N__16806),
            .lcout(\Lab_UT.dictrl.next_state_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18020),
            .ce(N__14383),
            .sr(N__13894));
    defparam \Lab_UT.dictrl.state_ret_4_RNI4Q509_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNI4Q509_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNI4Q509_LC_7_14_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNI4Q509_LC_7_14_3  (
            .in0(N__14261),
            .in1(N__14281),
            .in2(N__16887),
            .in3(N__14311),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_7_14_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI95NC1_0_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__11614),
            .in2(_gnd_net_),
            .in3(N__16940),
            .lcout(\Lab_UT.dictrl.next_state_RNI95NC1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIO0LS1_1_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIO0LS1_1_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIO0LS1_1_LC_7_14_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIO0LS1_1_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__14395),
            .in2(_gnd_net_),
            .in3(N__14445),
            .lcout(\Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_state_RNIO0LS1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNIRRERA_LC_7_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNIRRERA_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNIRRERA_LC_7_14_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNIRRERA_LC_7_14_6  (
            .in0(N__14416),
            .in1(N__16867),
            .in2(N__11608),
            .in3(N__14446),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNINI42G_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNINI42G_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNINI42G_LC_7_14_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNINI42G_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11605),
            .in3(N__14072),
            .lcout(\Lab_UT.dictrl.dicRun_2_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_2_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_8_2_0 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_8_2_0  (
            .in0(N__12017),
            .in1(N__11665),
            .in2(N__12081),
            .in3(N__12048),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18096),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_8_2_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_8_2_2 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_8_2_2  (
            .in0(N__12018),
            .in1(N__12047),
            .in2(N__12082),
            .in3(N__12142),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18096),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_8_2_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_8_2_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_8_2_3  (
            .in0(N__12135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12016),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18096),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNILM873_4_LC_8_2_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNILM873_4_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNILM873_4_LC_8_2_4 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \buart.Z_rx.bitcount_RNILM873_4_LC_8_2_4  (
            .in0(N__12073),
            .in1(N__12046),
            .in2(N__11833),
            .in3(N__11805),
            .lcout(\buart.Z_rx.bitcountlde_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNIU4N1_2_LC_8_2_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNIU4N1_2_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNIU4N1_2_LC_8_2_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNIU4N1_2_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__11677),
            .in2(_gnd_net_),
            .in3(N__12134),
            .lcout(\buart.Z_rx.ser_clk_2 ),
            .ltout(\buart.Z_rx.ser_clk_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_2_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_2_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.bitcount_RNIC77M1_0_LC_8_2_7  (
            .in0(N__12045),
            .in1(N__11755),
            .in2(N__11749),
            .in3(N__11745),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_8_3_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_8_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_8_3_0  (
            .in0(_gnd_net_),
            .in1(N__12092),
            .in2(N__12136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_8_3_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_8_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_2_LC_8_3_1  (
            .in0(_gnd_net_),
            .in1(N__11676),
            .in2(_gnd_net_),
            .in3(N__11659),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_8_3_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_8_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_8_3_2  (
            .in0(N__12026),
            .in1(N__12114),
            .in2(_gnd_net_),
            .in3(N__11656),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__18092),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_8_3_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_8_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_4_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__11959),
            .in2(_gnd_net_),
            .in3(N__11653),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_8_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_8_3_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNO_0_5_LC_8_3_4  (
            .in0(N__12105),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12145),
            .lcout(\buart.Z_rx.Z_baudgen.counter_RNO_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_3_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_8_3_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_8_3_5  (
            .in0(N__12094),
            .in1(N__12133),
            .in2(_gnd_net_),
            .in3(N__12028),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18092),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_8_3_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_8_3_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_8_3_6  (
            .in0(N__11958),
            .in1(N__12115),
            .in2(N__12106),
            .in3(N__12093),
            .lcout(\buart.Z_rx.ser_clk_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_8_3_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_8_3_7 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_8_3_7  (
            .in0(N__12080),
            .in1(N__12058),
            .in2(N__12052),
            .in3(N__12027),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18092),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_8_5_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_8_5_0  (
            .in0(N__17293),
            .in1(N__11950),
            .in2(N__17336),
            .in3(N__15486),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18074),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m24_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.m24_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m24_LC_8_5_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.didp.m24_LC_8_5_1  (
            .in0(N__15382),
            .in1(N__15174),
            .in2(_gnd_net_),
            .in3(N__15271),
            .lcout(\Lab_UT.m24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_8_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_8_5_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNINJD5_3_LC_8_5_2  (
            .in0(N__12660),
            .in1(N__11932),
            .in2(N__11914),
            .in3(N__11874),
            .lcout(\uu2.w_addr_user_3_i_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_8_5_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_8_5_5  (
            .in0(N__12540),
            .in1(N__12281),
            .in2(_gnd_net_),
            .in3(N__13410),
            .lcout(\uu2.mem0.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_5_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_8_5_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_8_5_7  (
            .in0(N__13747),
            .in1(N__12280),
            .in2(_gnd_net_),
            .in3(N__12661),
            .lcout(\uu2.mem0.N_74_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_8_6_0 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_8_6_0  (
            .in0(N__15029),
            .in1(N__15037),
            .in2(N__12610),
            .in3(N__16481),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18068),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_8_6_1 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_8_6_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \uu2.un28_w_addr_user_i_0_o2_0_LC_8_6_1  (
            .in0(N__14721),
            .in1(N__14655),
            .in2(N__14676),
            .in3(N__14777),
            .lcout(\uu2.N_84 ),
            .ltout(\uu2.N_84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_a3_LC_8_6_2 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a3_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a3_LC_8_6_2 .LUT_INIT=16'b0000001000000100;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a3_LC_8_6_2  (
            .in0(N__14700),
            .in1(N__14977),
            .in2(N__12601),
            .in3(N__12458),
            .lcout(\uu2.N_97 ),
            .ltout(\uu2.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI7BP14_6_LC_8_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI7BP14_6_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI7BP14_6_LC_8_6_3 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \uu2.w_addr_user_nesr_RNI7BP14_6_LC_8_6_3  (
            .in0(N__12396),
            .in1(N__12553),
            .in2(N__12517),
            .in3(N__12510),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_data_0_o2_0_4_LC_8_6_4 .C_ON=1'b0;
    defparam \uu2.w_data_0_o2_0_4_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_data_0_o2_0_4_LC_8_6_4 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \uu2.w_data_0_o2_0_4_LC_8_6_4  (
            .in0(N__14699),
            .in1(N__14976),
            .in2(_gnd_net_),
            .in3(N__12457),
            .lcout(\uu2.N_86 ),
            .ltout(\uu2.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_i_0_tz_0_LC_8_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_i_0_tz_0_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_i_0_tz_0_LC_8_6_5 .LUT_INIT=16'b0101010101011111;
    LogicCell40 \uu2.w_addr_i_0_tz_0_LC_8_6_5  (
            .in0(N__12395),
            .in1(_gnd_net_),
            .in2(N__12382),
            .in3(N__12365),
            .lcout(\uu2.w_addr_i_0_tzZ0Z_0 ),
            .ltout(\uu2.w_addr_i_0_tzZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIVAPV6_8_LC_8_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIVAPV6_8_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIVAPV6_8_LC_8_6_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIVAPV6_8_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12253),
            .in3(N__12246),
            .lcout(\uu2.un21_w_addr_displaying_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIRJ7L_3_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIRJ7L_3_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIRJ7L_3_LC_8_6_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIRJ7L_3_LC_8_6_7  (
            .in0(N__15377),
            .in1(N__15170),
            .in2(_gnd_net_),
            .in3(N__15241),
            .lcout(\Lab_UT.dispString.un22_dOutP ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_3_LC_8_7_0 .LUT_INIT=16'b1111101010101010;
    LogicCell40 \Lab_UT.didp.reset_3_LC_8_7_0  (
            .in0(N__17638),
            .in1(_gnd_net_),
            .in2(N__15655),
            .in3(N__14323),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18063),
            .ce(),
            .sr(N__17126));
    defparam \Lab_UT.didp.reset_2_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_2_LC_8_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.reset_2_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__15651),
            .in2(_gnd_net_),
            .in3(N__17637),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18063),
            .ce(),
            .sr(N__17126));
    defparam \uu2.w_addr_displaying_RNI8BP31_6_LC_8_7_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8BP31_6_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8BP31_6_LC_8_7_7 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \uu2.w_addr_displaying_RNI8BP31_6_LC_8_7_7  (
            .in0(N__13746),
            .in1(N__13411),
            .in2(_gnd_net_),
            .in3(N__13212),
            .lcout(\uu2.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_8_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_51_LC_8_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_51_LC_8_8_0  (
            .in0(N__13501),
            .in1(N__13062),
            .in2(N__13751),
            .in3(N__13287),
            .lcout(),
            .ltout(\uu2.mem0.g0_7_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_8_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_31_LC_8_8_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_31_LC_8_8_1  (
            .in0(N__13846),
            .in1(N__12971),
            .in2(N__13090),
            .in3(N__12893),
            .lcout(),
            .ltout(\uu2.mem0.un31_w_data_displaying_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_8_8_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_19_LC_8_8_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_19_LC_8_8_2  (
            .in0(N__12748),
            .in1(N__12754),
            .in2(N__13087),
            .in3(N__13288),
            .lcout(\uu2.mem0.g1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_29_LC_8_8_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_29_LC_8_8_3  (
            .in0(N__13063),
            .in1(N__12970),
            .in2(N__13626),
            .in3(N__12892),
            .lcout(\uu2.mem0.g1_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_30_LC_8_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_30_LC_8_8_4  (
            .in0(N__13204),
            .in1(N__13500),
            .in2(N__13409),
            .in3(N__13739),
            .lcout(\uu2.mem0.g1_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_8_8_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_50_LC_8_8_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_50_LC_8_8_5  (
            .in0(N__12740),
            .in1(N__13398),
            .in2(_gnd_net_),
            .in3(N__13203),
            .lcout(\uu2.mem0.g0_7_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_5_LC_8_8_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_5_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_5_LC_8_8_6 .LUT_INIT=16'b1001101010101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_5_LC_8_8_6  (
            .in0(N__13205),
            .in1(N__13838),
            .in2(N__13752),
            .in3(N__13609),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_5C_net ),
            .ce(N__13534),
            .sr(N__17783));
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_8_8_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_39_LC_8_8_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_39_LC_8_8_7  (
            .in0(N__13499),
            .in1(N__13397),
            .in2(N__13305),
            .in3(N__13202),
            .lcout(\uu2.mem0.g0_16_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.segment_1_1_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.segment_1_1_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.segment_1_1_LC_8_9_0 .LUT_INIT=16'b0001110111010111;
    LogicCell40 \Lab_UT.bcd2segment1.segment_1_1_LC_8_9_0  (
            .in0(N__16611),
            .in1(N__16460),
            .in2(N__16406),
            .in3(N__16548),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment1.segment_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_8_9_1 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_8_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu2.bitmap_93_LC_8_9_1  (
            .in0(N__14208),
            .in1(_gnd_net_),
            .in2(N__13132),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__17791));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_8_9_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_8_9_3  (
            .in0(N__16461),
            .in1(_gnd_net_),
            .in2(N__16569),
            .in3(N__16613),
            .lcout(\Lab_UT.didp.countrce1.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.un1_num_11_LC_8_9_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.bcd2segment1.un1_num_11_LC_8_9_4  (
            .in0(N__16612),
            .in1(N__16459),
            .in2(N__16407),
            .in3(N__16549),
            .lcout(\Lab_UT.nine ),
            .ltout(\Lab_UT.nine_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_3_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_3_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI84NN1_3_LC_8_9_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI84NN1_3_LC_8_9_5  (
            .in0(N__17551),
            .in1(N__16160),
            .in2(N__13114),
            .in3(N__16711),
            .lcout(\Lab_UT.didp.q_RNI84NN1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment2.segment_i_1_1_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment2.segment_i_1_1_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment2.segment_i_1_1_LC_8_9_6 .LUT_INIT=16'b0001000011111111;
    LogicCell40 \Lab_UT.bcd2segment2.segment_i_1_1_LC_8_9_6  (
            .in0(N__16710),
            .in1(N__17550),
            .in2(N__16172),
            .in3(N__14207),
            .lcout(),
            .ltout(\Lab_UT.bcd2segment2.segment_i_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_8_9_7 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_8_9_7 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \uu2.bitmap_87_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__13873),
            .in2(N__13867),
            .in3(_gnd_net_),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__17791));
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_10_0 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_8_10_0  (
            .in0(N__17145),
            .in1(N__16554),
            .in2(N__16671),
            .in3(N__16467),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_8_10_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_8_10_1  (
            .in0(N__16466),
            .in1(N__17143),
            .in2(_gnd_net_),
            .in3(N__16663),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment1.un1_num_5_2_LC_8_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.bcd2segment1.un1_num_5_2_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__16553),
            .in2(_gnd_net_),
            .in3(N__16465),
            .lcout(),
            .ltout(\Lab_UT.three_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_10_3 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_8_10_3  (
            .in0(N__16667),
            .in1(N__17146),
            .in2(N__13855),
            .in3(N__16617),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_10_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_8_10_4  (
            .in0(N__16341),
            .in1(N__16180),
            .in2(N__15855),
            .in3(N__16162),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_10_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_8_10_5  (
            .in0(N__16340),
            .in1(N__16087),
            .in2(N__17560),
            .in3(N__15851),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_10_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_8_10_6  (
            .in0(N__15847),
            .in1(N__16339),
            .in2(_gnd_net_),
            .in3(N__16239),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_8_10_7 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_8_10_7  (
            .in0(N__13852),
            .in1(N__17144),
            .in2(N__16672),
            .in3(N__16397),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18045),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_set_0_1_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_set_0_1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_set_0_1_LC_8_11_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.next_state_set_0_1_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__14006),
            .in2(_gnd_net_),
            .in3(N__14040),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_set_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNILGF17_3_LC_8_11_2 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNILGF17_3_LC_8_11_2  (
            .in0(N__14547),
            .in1(N__14751),
            .in2(N__14059),
            .in3(N__14056),
            .lcout(\Lab_UT.dictrl.next_state_set_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m34_ns_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.m34_ns_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m34_ns_LC_8_11_3 .LUT_INIT=16'b0100000011101010;
    LogicCell40 \Lab_UT.didp.m34_ns_LC_8_11_3  (
            .in0(N__14601),
            .in1(N__14635),
            .in2(N__14548),
            .in3(N__14050),
            .lcout(\Lab_UT.m34_ns ),
            .ltout(\Lab_UT.m34_ns_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIM00A3_3_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIM00A3_3_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIM00A3_3_LC_8_11_4 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIM00A3_3_LC_8_11_4  (
            .in0(N__14041),
            .in1(N__14546),
            .in2(N__14020),
            .in3(N__14007),
            .lcout(\Lab_UT.dictrl.next_state_set_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_11_5 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_8_11_5  (
            .in0(N__17219),
            .in1(N__14917),
            .in2(N__17365),
            .in3(N__13990),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_8_11_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_8_11_6  (
            .in0(N__14918),
            .in1(N__17335),
            .in2(N__13954),
            .in3(N__17292),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18038),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_8_11_7 .C_ON=1'b0;
    defparam \resetGen.rst_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_8_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13951),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18038),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_12_0 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_12_0 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_8_12_0  (
            .in0(N__14496),
            .in1(N__15593),
            .in2(N__15640),
            .in3(N__15565),
            .lcout(\Lab_UT.dictrl.next_state_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18032),
            .ce(N__14388),
            .sr(N__13906));
    defparam \Lab_UT.didp.m41_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.m41_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m41_LC_8_12_1 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \Lab_UT.didp.m41_LC_8_12_1  (
            .in0(N__14529),
            .in1(N__14630),
            .in2(_gnd_net_),
            .in3(N__16780),
            .lcout(),
            .ltout(\Lab_UT.didp.N_164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m42_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.m42_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m42_LC_8_12_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \Lab_UT.didp.m42_LC_8_12_2  (
            .in0(N__16781),
            .in1(N__14597),
            .in2(N__13897),
            .in3(N__17015),
            .lcout(\Lab_UT.m42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_12_3 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_2_LC_8_12_3  (
            .in0(N__15488),
            .in1(N__14914),
            .in2(_gnd_net_),
            .in3(N__17214),
            .lcout(\Lab_UT.didp.countrce4.N_88_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_RNICI8U_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_RNICI8U_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_RNICI8U_LC_8_12_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_RNICI8U_LC_8_12_5  (
            .in0(N__17016),
            .in1(N__14631),
            .in2(N__14605),
            .in3(N__16782),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_8_12_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_8_12_7  (
            .in0(N__15489),
            .in1(N__14343),
            .in2(_gnd_net_),
            .in3(N__17215),
            .lcout(\Lab_UT.didp.un31_reset_i_a4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_13_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_LC_8_13_0 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_LC_8_13_0  (
            .in0(N__14418),
            .in1(N__16897),
            .in2(N__14470),
            .in3(N__14449),
            .lcout(\Lab_UT.state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_0_1_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_LC_8_13_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_LC_8_13_1  (
            .in0(N__14448),
            .in1(N__14465),
            .in2(N__16912),
            .in3(N__14417),
            .lcout(\Lab_UT.state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_13_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_13_2 .LUT_INIT=16'b1010001111110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_8_13_2  (
            .in0(N__14263),
            .in1(N__14286),
            .in2(N__16913),
            .in3(N__14310),
            .lcout(\Lab_UT.dictrl.state_i_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_0_2_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_LC_8_13_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_LC_8_13_3  (
            .in0(N__14309),
            .in1(N__16901),
            .in2(N__14287),
            .in3(N__14262),
            .lcout(\Lab_UT.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_8_13_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_RNIGOKU_LC_8_13_4  (
            .in0(N__17041),
            .in1(N__16755),
            .in2(_gnd_net_),
            .in3(N__17162),
            .lcout(\Lab_UT.Run ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_13_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_LC_8_13_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_LC_8_13_5  (
            .in0(_gnd_net_),
            .in1(N__14086),
            .in2(_gnd_net_),
            .in3(N__14074),
            .lcout(\Lab_UT.dictrl.dicRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_0_3_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_LC_8_13_7 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_LC_8_13_7  (
            .in0(N__16896),
            .in1(N__15570),
            .in2(N__15600),
            .in3(N__15638),
            .lcout(\Lab_UT.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18027),
            .ce(),
            .sr(N__17812));
    defparam \Lab_UT.dictrl.state_ret_3_RNI2T7U_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNI2T7U_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNI2T7U_LC_8_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNI2T7U_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(N__14627),
            .in2(_gnd_net_),
            .in3(N__17042),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_state_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNITFCD1_1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNITFCD1_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNITFCD1_1_LC_8_14_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.state_0_RNITFCD1_1_LC_8_14_1  (
            .in0(N__16760),
            .in1(N__17080),
            .in2(N__14644),
            .in3(N__17019),
            .lcout(\Lab_UT.dictrl.state_0_RNITFCD1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m37_ns_1_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.m37_ns_1_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m37_ns_1_LC_8_14_2 .LUT_INIT=16'b0001000110111110;
    LogicCell40 \Lab_UT.didp.m37_ns_1_LC_8_14_2  (
            .in0(N__14583),
            .in1(N__14629),
            .in2(N__14542),
            .in3(N__16759),
            .lcout(\Lab_UT.didp.m37_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_RNI0P1V_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_RNI0P1V_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_RNI0P1V_LC_8_14_3 .LUT_INIT=16'b0001001111011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_RNI0P1V_LC_8_14_3  (
            .in0(N__14628),
            .in1(N__14582),
            .in2(N__14541),
            .in3(N__17163),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_state_24_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_RNIRB6E1_1_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_RNIRB6E1_1_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_RNIRB6E1_1_LC_8_14_4 .LUT_INIT=16'b1000100000001111;
    LogicCell40 \Lab_UT.dictrl.state_0_RNIRB6E1_1_LC_8_14_4  (
            .in0(N__17020),
            .in1(N__17079),
            .in2(N__14500),
            .in3(N__16761),
            .lcout(\Lab_UT.dictrl.state_0_RNIRB6E1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_8_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_RNINNUG_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__16914),
            .in2(_gnd_net_),
            .in3(N__17853),
            .lcout(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0 ),
            .ltout(\Lab_UT.dictrl.state_ret_4_RNINNUGZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_14_7 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_14_7 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_8_14_7  (
            .in0(N__14469),
            .in1(N__14447),
            .in2(N__14422),
            .in3(N__14419),
            .lcout(\Lab_UT.dictrl.next_state_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18023),
            .ce(N__14387),
            .sr(N__14755));
    defparam \Lab_UT.dispString.dOut_5_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_9_5_0 .LUT_INIT=16'b0010001011000100;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_9_5_0  (
            .in0(N__15375),
            .in1(N__15163),
            .in2(N__18277),
            .in3(N__15270),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18085),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m28_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.m28_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m28_LC_9_5_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.didp.m28_LC_9_5_2  (
            .in0(N__15371),
            .in1(N__15155),
            .in2(_gnd_net_),
            .in3(N__15266),
            .lcout(\Lab_UT.un29_dOutP ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_9_5_3 .LUT_INIT=16'b1110011111000111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_9_5_3  (
            .in0(N__15268),
            .in1(N__15373),
            .in2(N__15173),
            .in3(N__16174),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_9_5_4 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_9_5_4  (
            .in0(N__15028),
            .in1(N__15412),
            .in2(N__14710),
            .in3(N__16646),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18085),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_9_5_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_9_5_5  (
            .in0(N__17659),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14831),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18085),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_9_5_6 .LUT_INIT=16'b0000000011000100;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_9_5_6  (
            .in0(N__15374),
            .in1(N__15162),
            .in2(N__16723),
            .in3(N__15269),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18085),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_9_5_7 .LUT_INIT=16'b1110110111101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_9_5_7  (
            .in0(N__15267),
            .in1(N__15372),
            .in2(N__15172),
            .in3(N__15813),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_9_6_0 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_9_6_0  (
            .in0(N__15402),
            .in1(N__16419),
            .in2(N__15030),
            .in3(N__17493),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.G_64_a0_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.G_64_a0_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.G_64_a0_LC_9_6_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.bcd2segment4.G_64_a0_LC_9_6_3  (
            .in0(N__14845),
            .in1(N__17404),
            .in2(N__15487),
            .in3(N__15073),
            .lcout(\Lab_UT.alarmMatch ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_9_6_4 .LUT_INIT=16'b1110111111100101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_9_6_4  (
            .in0(N__15242),
            .in1(N__14761),
            .in2(N__15178),
            .in3(N__15726),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_9_6_5 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__15401),
            .in2(N__15040),
            .in3(N__17230),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_9_6_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_9_6_6  (
            .in0(N__15403),
            .in1(N__16576),
            .in2(N__15031),
            .in3(N__14942),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_9_6_7 .LUT_INIT=16'b0011111111111111;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__15004),
            .in2(N__14998),
            .in3(N__14953),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18075),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_9_7_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_9_7_0  (
            .in0(N__16321),
            .in1(N__14838),
            .in2(N__15087),
            .in3(N__14814),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_0_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_0_LC_9_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.bcd2segment4.G_64_a0_1_0_LC_9_7_1  (
            .in0(N__14919),
            .in1(N__16320),
            .in2(N__16173),
            .in3(N__16250),
            .lcout(\Lab_UT.bcd2segment4.G_64_a0_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_9_7_2 .LUT_INIT=16'b1111010100110001;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_9_7_2  (
            .in0(N__14839),
            .in1(N__14815),
            .in2(N__15088),
            .in3(N__17559),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_9_7_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_9_7_3  (
            .in0(N__14806),
            .in1(_gnd_net_),
            .in2(N__14797),
            .in3(N__15832),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18069),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_0_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_0_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_0_LC_9_7_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.alarmchar_0_LC_9_7_4  (
            .in0(N__18319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18262),
            .lcout(\Lab_UT.alarmcharZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18069),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_9_7_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_RNIL6V9_0_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__18261),
            .in2(_gnd_net_),
            .in3(N__18317),
            .lcout(),
            .ltout(\Lab_UT.alarmchar9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_2_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_2_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_2_LC_9_7_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.alarmchar_2_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15091),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmcharZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18069),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_1_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_1_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_1_LC_9_7_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.alarmchar_1_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__18127),
            .in2(_gnd_net_),
            .in3(N__18318),
            .lcout(\Lab_UT.alarmcharZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18069),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment3.un1_num_1_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment3.un1_num_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment3.un1_num_1_LC_9_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.bcd2segment3.un1_num_1_LC_9_8_0  (
            .in0(N__15943),
            .in1(N__15774),
            .in2(N__16047),
            .in3(N__15698),
            .lcout(\Lab_UT.zero ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_8_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_8_1  (
            .in0(N__15699),
            .in1(N__16026),
            .in2(N__15794),
            .in3(N__15945),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.qPone_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_8_2 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_9_8_2  (
            .in0(N__16698),
            .in1(N__16031),
            .in2(N__15064),
            .in3(N__15057),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18064),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_8_3 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_9_8_3  (
            .in0(N__15701),
            .in1(N__15058),
            .in2(N__15795),
            .in3(N__16699),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18064),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_8_4 .LUT_INIT=16'b1001100101010101;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_8_4  (
            .in0(N__15944),
            .in1(N__15778),
            .in2(_gnd_net_),
            .in3(N__15700),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.N_79_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_8_5 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_9_8_5  (
            .in0(N__15056),
            .in1(N__16697),
            .in2(N__15061),
            .in3(N__15946),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18064),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_8_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_9_8_6  (
            .in0(N__16696),
            .in1(N__15055),
            .in2(_gnd_net_),
            .in3(N__15702),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18064),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_9_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_9_8_7 .LUT_INIT=16'b1101111111011101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_9_8_7  (
            .in0(N__15265),
            .in1(N__15147),
            .in2(N__15376),
            .in3(N__16025),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_1_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_1_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_1_LC_9_9_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNI36SS_1_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__15773),
            .in2(_gnd_net_),
            .in3(N__15692),
            .lcout(\Lab_UT.N_207 ),
            .ltout(\Lab_UT.N_207_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIIKFH3_3_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIIKFH3_3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIIKFH3_3_LC_9_9_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIIKFH3_3_LC_9_9_1  (
            .in0(N__15879),
            .in1(N__16027),
            .in2(N__15658),
            .in3(N__15953),
            .lcout(\Lab_UT.didp.q_RNIIKFH3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_LC_9_9_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_LC_9_9_2 .LUT_INIT=16'b1000110110101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_LC_9_9_2  (
            .in0(N__16886),
            .in1(N__15639),
            .in2(N__15604),
            .in3(N__15574),
            .lcout(\Lab_UT.state_i_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18057),
            .ce(),
            .sr(N__17809));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_9_9_3 .LUT_INIT=16'b1110111011110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_9_9_3  (
            .in0(N__15541),
            .in1(N__15245),
            .in2(N__15985),
            .in3(N__15121),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_9_9_4 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_9_9_4  (
            .in0(N__15393),
            .in1(_gnd_net_),
            .in2(N__15532),
            .in3(N__15525),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.m29_LC_9_9_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.m29_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.m29_LC_9_9_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.didp.m29_LC_9_9_5  (
            .in0(N__15339),
            .in1(N__15120),
            .in2(_gnd_net_),
            .in3(N__15244),
            .lcout(\Lab_UT.un3_dOutP ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_3_LC_9_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_3_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_3_LC_9_9_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \Lab_UT.dispString.cnt_3_LC_9_9_6  (
            .in0(N__15247),
            .in1(N__15312),
            .in2(N__15148),
            .in3(N__15340),
            .lcout(\Lab_UT.cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18057),
            .ce(),
            .sr(N__17809));
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_9_9_7  (
            .in0(N__15311),
            .in1(N__15122),
            .in2(_gnd_net_),
            .in3(N__15246),
            .lcout(\Lab_UT.cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18057),
            .ce(),
            .sr(N__17809));
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_10_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__16312),
            .in2(_gnd_net_),
            .in3(N__16229),
            .lcout(\Lab_UT.N_204 ),
            .ltout(\Lab_UT.N_204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_2_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_9_10_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_9_10_1  (
            .in0(N__16681),
            .in1(N__16171),
            .in2(N__16702),
            .in3(N__17558),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18051),
            .ce(),
            .sr(N__17127));
    defparam \Lab_UT.didp.reset_0_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_0_LC_9_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.reset_0_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__16680),
            .in2(_gnd_net_),
            .in3(N__17856),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18051),
            .ce(),
            .sr(N__17127));
    defparam \Lab_UT.didp.ce_1_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_9_10_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_9_10_3  (
            .in0(N__16618),
            .in1(N__16558),
            .in2(N__16482),
            .in3(N__16398),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18051),
            .ce(),
            .sr(N__17127));
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_0_1_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_0_1_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_0_1_LC_9_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI1S78_0_1_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__16313),
            .in2(_gnd_net_),
            .in3(N__16230),
            .lcout(\Lab_UT.didp.countrce2.three_2 ),
            .ltout(\Lab_UT.didp.countrce2.three_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_10_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_10_5  (
            .in0(N__16161),
            .in1(_gnd_net_),
            .in2(N__16090),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.countrce2.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_3_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_9_10_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_9_10_6  (
            .in0(N__16048),
            .in1(N__15968),
            .in2(N__15880),
            .in3(N__15894),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18051),
            .ce(),
            .sr(N__17127));
    defparam \Lab_UT.didp.reset_1_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.reset_1_LC_9_10_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.didp.reset_1_LC_9_10_7  (
            .in0(N__17857),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15875),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18051),
            .ce(),
            .sr(N__17127));
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.G_64_a0_1_LC_9_11_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.bcd2segment4.G_64_a0_1_LC_9_11_0  (
            .in0(N__17547),
            .in1(N__17471),
            .in2(_gnd_net_),
            .in3(N__17201),
            .lcout(\Lab_UT.bcd2segment4.G_64_a0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_11_2 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_9_11_2  (
            .in0(N__17395),
            .in1(N__17202),
            .in2(_gnd_net_),
            .in3(N__17364),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_9_11_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_9_11_3  (
            .in0(N__17203),
            .in1(N__17340),
            .in2(N__17296),
            .in3(N__17275),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18046),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_0_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_9_12_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_9_12_0  (
            .in0(N__17044),
            .in1(N__16783),
            .in2(_gnd_net_),
            .in3(N__17164),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18039),
            .ce(),
            .sr(N__17128));
    defparam \Lab_UT.dictrl.state_ret_3_RNIDH8U_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNIDH8U_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNIDH8U_LC_9_13_6 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNIDH8U_LC_9_13_6  (
            .in0(N__17078),
            .in1(N__17043),
            .in2(N__17017),
            .in3(N__16772),
            .lcout(\Lab_UT.dictrl.state_ret_3_RNIDH8UZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_LC_9_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_LC_9_14_3 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_0_LC_9_14_3  (
            .in0(N__16963),
            .in1(N__16932),
            .in2(N__16918),
            .in3(N__16810),
            .lcout(\Lab_UT.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18028),
            .ce(),
            .sr(N__17813));
    defparam \Lab_UT.alarmchar_4_LC_11_5_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_4_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_4_LC_11_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.alarmchar_4_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18373),
            .lcout(\Lab_UT.alarmcharZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18093),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_11_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_11_5_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__18126),
            .in2(_gnd_net_),
            .in3(N__18316),
            .lcout(),
            .ltout(\Lab_UT.alarmchar_2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_6_LC_11_5_6 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_6_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_6_LC_11_5_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \Lab_UT.alarmchar_6_LC_11_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17662),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmcharZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18093),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_11_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_11_6_0 .LUT_INIT=16'b1100000011000101;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNIA99N6_0_LC_11_6_0  (
            .in0(N__18330),
            .in1(N__18217),
            .in2(N__18190),
            .in3(N__18353),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1 ),
            .ltout(\Lab_UT.dictrl.next_alarmstate_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_11_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_3_LC_11_6_1 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_3_LC_11_6_1  (
            .in0(N__17646),
            .in1(_gnd_net_),
            .in2(N__17650),
            .in3(N__17587),
            .lcout(\Lab_UT.un1_next_alarmstate21_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18086),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.G_3_LC_11_6_2 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.G_3_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.G_3_LC_11_6_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.bcd2segment4.G_3_LC_11_6_2  (
            .in0(N__18305),
            .in1(N__18354),
            .in2(N__18232),
            .in3(N__17645),
            .lcout(),
            .ltout(\Lab_UT.G_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_11_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_alarmstate_0_LC_11_6_3 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_0_LC_11_6_3  (
            .in0(N__17581),
            .in1(_gnd_net_),
            .in2(N__17593),
            .in3(N__18216),
            .lcout(\Lab_UT.dictrl.next_alarmstate_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18086),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_11_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_11_6_4 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_1_1_0__m4_LC_11_6_4  (
            .in0(N__17566),
            .in1(N__18352),
            .in2(N__18260),
            .in3(N__17580),
            .lcout(\Lab_UT.dictrl.next_alarmstate_1_0 ),
            .ltout(\Lab_UT.dictrl.next_alarmstate_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_11_6_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.next_alarmstate_RNI4S8S6_0_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__18215),
            .in2(N__17590),
            .in3(N__18181),
            .lcout(\Lab_UT.dictrl.next_alarmstateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_11_6_6 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI6ASS3_LC_11_6_6  (
            .in0(N__18304),
            .in1(N__18119),
            .in2(_gnd_net_),
            .in3(N__17579),
            .lcout(\Lab_UT.dictrl.next_alarmstate_latmux_0_mb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_11_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_11_6_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_RNI8PIF_0_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(N__18118),
            .in2(_gnd_net_),
            .in3(N__18303),
            .lcout(\Lab_UT.dictrl.idle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_ret_1_LC_11_7_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_1_LC_11_7_0  (
            .in0(N__18188),
            .in1(N__18146),
            .in2(_gnd_net_),
            .in3(N__18363),
            .lcout(\Lab_UT.alarmchar10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18077),
            .ce(),
            .sr(N__17810));
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_11_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_11_7_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_2_LC_11_7_1 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_2_LC_11_7_1  (
            .in0(N__18364),
            .in1(N__18189),
            .in2(_gnd_net_),
            .in3(N__18148),
            .lcout(\Lab_UT.alarmchar10_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18077),
            .ce(),
            .sr(N__17810));
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_0_LC_11_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_0_LC_11_7_4  (
            .in0(N__18218),
            .in1(N__18185),
            .in2(_gnd_net_),
            .in3(N__18145),
            .lcout(\Lab_UT.alarmstate_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18077),
            .ce(),
            .sr(N__17810));
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_11_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.alarmstate_0_1_LC_11_7_6 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_0_1_LC_11_7_6  (
            .in0(N__18187),
            .in1(N__18355),
            .in2(N__18223),
            .in3(N__18331),
            .lcout(\Lab_UT.alarmstate_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18077),
            .ce(),
            .sr(N__17810));
    defparam \Lab_UT.alarmchar_5_LC_11_8_0 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_5_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.alarmchar_5_LC_11_8_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \Lab_UT.alarmchar_5_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__18283),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.alarmcharZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18070),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.bcd2segment4.G_1_LC_12_6_7 .C_ON=1'b0;
    defparam \Lab_UT.bcd2segment4.G_1_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.bcd2segment4.G_1_LC_12_6_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.bcd2segment4.G_1_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__18180),
            .in2(_gnd_net_),
            .in3(N__18253),
            .lcout(\Lab_UT.bcd2segment4.GZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_12_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_12_7_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.alarmstate_ret_LC_12_7_2 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \Lab_UT.dictrl.alarmstate_ret_LC_12_7_2  (
            .in0(N__18222),
            .in1(N__18186),
            .in2(_gnd_net_),
            .in3(N__18147),
            .lcout(\Lab_UT.dictrl.alarmstate_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18087),
            .ce(),
            .sr(N__17811));
endmodule // latticehx1k
