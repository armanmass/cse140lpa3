// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 20 2019 23:36:29

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__23173;
    wire N__23172;
    wire N__23171;
    wire N__23164;
    wire N__23163;
    wire N__23162;
    wire N__23155;
    wire N__23154;
    wire N__23153;
    wire N__23146;
    wire N__23145;
    wire N__23144;
    wire N__23137;
    wire N__23136;
    wire N__23135;
    wire N__23128;
    wire N__23127;
    wire N__23126;
    wire N__23119;
    wire N__23118;
    wire N__23117;
    wire N__23110;
    wire N__23109;
    wire N__23108;
    wire N__23101;
    wire N__23100;
    wire N__23099;
    wire N__23092;
    wire N__23091;
    wire N__23090;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23063;
    wire N__23060;
    wire N__23057;
    wire N__23052;
    wire N__23049;
    wire N__23048;
    wire N__23047;
    wire N__23044;
    wire N__23039;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23021;
    wire N__23020;
    wire N__23017;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22989;
    wire N__22988;
    wire N__22987;
    wire N__22984;
    wire N__22983;
    wire N__22982;
    wire N__22981;
    wire N__22980;
    wire N__22975;
    wire N__22970;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22932;
    wire N__22929;
    wire N__22928;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22914;
    wire N__22911;
    wire N__22908;
    wire N__22907;
    wire N__22904;
    wire N__22901;
    wire N__22900;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22882;
    wire N__22877;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22851;
    wire N__22850;
    wire N__22849;
    wire N__22848;
    wire N__22847;
    wire N__22846;
    wire N__22845;
    wire N__22844;
    wire N__22843;
    wire N__22842;
    wire N__22841;
    wire N__22840;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22836;
    wire N__22835;
    wire N__22834;
    wire N__22833;
    wire N__22832;
    wire N__22831;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22824;
    wire N__22823;
    wire N__22822;
    wire N__22821;
    wire N__22820;
    wire N__22819;
    wire N__22818;
    wire N__22817;
    wire N__22816;
    wire N__22815;
    wire N__22814;
    wire N__22813;
    wire N__22812;
    wire N__22811;
    wire N__22810;
    wire N__22809;
    wire N__22808;
    wire N__22807;
    wire N__22806;
    wire N__22805;
    wire N__22804;
    wire N__22803;
    wire N__22802;
    wire N__22801;
    wire N__22800;
    wire N__22799;
    wire N__22798;
    wire N__22797;
    wire N__22796;
    wire N__22795;
    wire N__22794;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22790;
    wire N__22789;
    wire N__22788;
    wire N__22787;
    wire N__22786;
    wire N__22785;
    wire N__22784;
    wire N__22783;
    wire N__22782;
    wire N__22781;
    wire N__22780;
    wire N__22779;
    wire N__22778;
    wire N__22777;
    wire N__22776;
    wire N__22775;
    wire N__22774;
    wire N__22771;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22567;
    wire N__22560;
    wire N__22559;
    wire N__22558;
    wire N__22557;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22534;
    wire N__22533;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22527;
    wire N__22526;
    wire N__22525;
    wire N__22524;
    wire N__22523;
    wire N__22522;
    wire N__22521;
    wire N__22520;
    wire N__22519;
    wire N__22518;
    wire N__22517;
    wire N__22516;
    wire N__22515;
    wire N__22514;
    wire N__22513;
    wire N__22512;
    wire N__22511;
    wire N__22510;
    wire N__22509;
    wire N__22508;
    wire N__22507;
    wire N__22506;
    wire N__22505;
    wire N__22504;
    wire N__22503;
    wire N__22502;
    wire N__22501;
    wire N__22500;
    wire N__22499;
    wire N__22498;
    wire N__22497;
    wire N__22496;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22484;
    wire N__22483;
    wire N__22482;
    wire N__22481;
    wire N__22480;
    wire N__22479;
    wire N__22478;
    wire N__22477;
    wire N__22476;
    wire N__22475;
    wire N__22474;
    wire N__22473;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22299;
    wire N__22296;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22282;
    wire N__22277;
    wire N__22274;
    wire N__22269;
    wire N__22268;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22237;
    wire N__22234;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22193;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22173;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22137;
    wire N__22134;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22106;
    wire N__22105;
    wire N__22104;
    wire N__22103;
    wire N__22098;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22092;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22065;
    wire N__22062;
    wire N__22057;
    wire N__22056;
    wire N__22049;
    wire N__22044;
    wire N__22041;
    wire N__22040;
    wire N__22039;
    wire N__22038;
    wire N__22033;
    wire N__22024;
    wire N__22021;
    wire N__22020;
    wire N__22017;
    wire N__22012;
    wire N__22009;
    wire N__22004;
    wire N__21997;
    wire N__21994;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21937;
    wire N__21936;
    wire N__21935;
    wire N__21932;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21913;
    wire N__21912;
    wire N__21911;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21903;
    wire N__21900;
    wire N__21899;
    wire N__21898;
    wire N__21897;
    wire N__21890;
    wire N__21887;
    wire N__21886;
    wire N__21885;
    wire N__21882;
    wire N__21881;
    wire N__21880;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21840;
    wire N__21839;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21835;
    wire N__21832;
    wire N__21827;
    wire N__21824;
    wire N__21821;
    wire N__21820;
    wire N__21817;
    wire N__21802;
    wire N__21787;
    wire N__21782;
    wire N__21779;
    wire N__21774;
    wire N__21767;
    wire N__21760;
    wire N__21757;
    wire N__21750;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21728;
    wire N__21725;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21721;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21699;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21664;
    wire N__21657;
    wire N__21656;
    wire N__21653;
    wire N__21652;
    wire N__21651;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21632;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21621;
    wire N__21614;
    wire N__21607;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21589;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21561;
    wire N__21560;
    wire N__21557;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21546;
    wire N__21545;
    wire N__21544;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21532;
    wire N__21531;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21506;
    wire N__21503;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21491;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21475;
    wire N__21466;
    wire N__21459;
    wire N__21456;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21401;
    wire N__21398;
    wire N__21387;
    wire N__21386;
    wire N__21385;
    wire N__21384;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21370;
    wire N__21369;
    wire N__21368;
    wire N__21367;
    wire N__21366;
    wire N__21365;
    wire N__21364;
    wire N__21363;
    wire N__21360;
    wire N__21359;
    wire N__21358;
    wire N__21357;
    wire N__21356;
    wire N__21355;
    wire N__21354;
    wire N__21349;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21317;
    wire N__21308;
    wire N__21303;
    wire N__21300;
    wire N__21299;
    wire N__21298;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21289;
    wire N__21284;
    wire N__21281;
    wire N__21274;
    wire N__21271;
    wire N__21264;
    wire N__21255;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21227;
    wire N__21220;
    wire N__21217;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21167;
    wire N__21164;
    wire N__21159;
    wire N__21158;
    wire N__21157;
    wire N__21154;
    wire N__21153;
    wire N__21150;
    wire N__21149;
    wire N__21148;
    wire N__21147;
    wire N__21146;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21120;
    wire N__21117;
    wire N__21108;
    wire N__21103;
    wire N__21100;
    wire N__21095;
    wire N__21088;
    wire N__21081;
    wire N__21078;
    wire N__21077;
    wire N__21074;
    wire N__21073;
    wire N__21072;
    wire N__21071;
    wire N__21070;
    wire N__21069;
    wire N__21066;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21059;
    wire N__21048;
    wire N__21045;
    wire N__21040;
    wire N__21039;
    wire N__21038;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21021;
    wire N__21018;
    wire N__21013;
    wire N__21006;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20984;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20965;
    wire N__20964;
    wire N__20963;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20938;
    wire N__20927;
    wire N__20924;
    wire N__20921;
    wire N__20916;
    wire N__20905;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20887;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20865;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20857;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20853;
    wire N__20852;
    wire N__20851;
    wire N__20848;
    wire N__20845;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20820;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20801;
    wire N__20800;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20784;
    wire N__20781;
    wire N__20780;
    wire N__20779;
    wire N__20774;
    wire N__20767;
    wire N__20760;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20741;
    wire N__20738;
    wire N__20733;
    wire N__20730;
    wire N__20723;
    wire N__20706;
    wire N__20705;
    wire N__20704;
    wire N__20703;
    wire N__20702;
    wire N__20699;
    wire N__20696;
    wire N__20693;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20677;
    wire N__20672;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20653;
    wire N__20652;
    wire N__20651;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20641;
    wire N__20638;
    wire N__20637;
    wire N__20636;
    wire N__20633;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20620;
    wire N__20617;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20582;
    wire N__20581;
    wire N__20578;
    wire N__20573;
    wire N__20568;
    wire N__20565;
    wire N__20564;
    wire N__20563;
    wire N__20562;
    wire N__20559;
    wire N__20552;
    wire N__20547;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20537;
    wire N__20532;
    wire N__20531;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20510;
    wire N__20509;
    wire N__20506;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20490;
    wire N__20487;
    wire N__20486;
    wire N__20485;
    wire N__20482;
    wire N__20481;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20469;
    wire N__20468;
    wire N__20465;
    wire N__20460;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20414;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20372;
    wire N__20371;
    wire N__20370;
    wire N__20369;
    wire N__20368;
    wire N__20367;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20352;
    wire N__20351;
    wire N__20348;
    wire N__20347;
    wire N__20346;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20305;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20295;
    wire N__20292;
    wire N__20287;
    wire N__20282;
    wire N__20279;
    wire N__20274;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20252;
    wire N__20249;
    wire N__20246;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20230;
    wire N__20221;
    wire N__20218;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20183;
    wire N__20182;
    wire N__20181;
    wire N__20180;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20175;
    wire N__20174;
    wire N__20169;
    wire N__20168;
    wire N__20165;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20118;
    wire N__20113;
    wire N__20104;
    wire N__20099;
    wire N__20096;
    wire N__20095;
    wire N__20092;
    wire N__20089;
    wire N__20078;
    wire N__20073;
    wire N__20066;
    wire N__20063;
    wire N__20054;
    wire N__20051;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19981;
    wire N__19974;
    wire N__19973;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19958;
    wire N__19955;
    wire N__19950;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19943;
    wire N__19942;
    wire N__19939;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19902;
    wire N__19901;
    wire N__19900;
    wire N__19899;
    wire N__19896;
    wire N__19895;
    wire N__19894;
    wire N__19893;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19884;
    wire N__19883;
    wire N__19882;
    wire N__19879;
    wire N__19876;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19838;
    wire N__19835;
    wire N__19832;
    wire N__19829;
    wire N__19822;
    wire N__19817;
    wire N__19814;
    wire N__19807;
    wire N__19800;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19789;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19781;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19771;
    wire N__19766;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19740;
    wire N__19737;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19726;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19714;
    wire N__19711;
    wire N__19704;
    wire N__19703;
    wire N__19702;
    wire N__19701;
    wire N__19700;
    wire N__19693;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19677;
    wire N__19676;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19650;
    wire N__19647;
    wire N__19646;
    wire N__19645;
    wire N__19644;
    wire N__19641;
    wire N__19640;
    wire N__19639;
    wire N__19638;
    wire N__19635;
    wire N__19630;
    wire N__19627;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19600;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19575;
    wire N__19572;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19547;
    wire N__19546;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19502;
    wire N__19499;
    wire N__19498;
    wire N__19491;
    wire N__19488;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19473;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19463;
    wire N__19456;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19438;
    wire N__19433;
    wire N__19430;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19418;
    wire N__19417;
    wire N__19416;
    wire N__19407;
    wire N__19404;
    wire N__19403;
    wire N__19402;
    wire N__19401;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19385;
    wire N__19380;
    wire N__19377;
    wire N__19376;
    wire N__19373;
    wire N__19372;
    wire N__19371;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19357;
    wire N__19350;
    wire N__19349;
    wire N__19346;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19292;
    wire N__19291;
    wire N__19290;
    wire N__19285;
    wire N__19280;
    wire N__19279;
    wire N__19274;
    wire N__19271;
    wire N__19268;
    wire N__19265;
    wire N__19260;
    wire N__19259;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19247;
    wire N__19244;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19197;
    wire N__19194;
    wire N__19187;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19172;
    wire N__19167;
    wire N__19166;
    wire N__19165;
    wire N__19162;
    wire N__19161;
    wire N__19158;
    wire N__19151;
    wire N__19148;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19128;
    wire N__19127;
    wire N__19126;
    wire N__19123;
    wire N__19122;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19079;
    wire N__19078;
    wire N__19077;
    wire N__19072;
    wire N__19069;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19057;
    wire N__19054;
    wire N__19047;
    wire N__19046;
    wire N__19045;
    wire N__19044;
    wire N__19041;
    wire N__19036;
    wire N__19033;
    wire N__19026;
    wire N__19025;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19017;
    wire N__19016;
    wire N__19013;
    wire N__19010;
    wire N__19003;
    wire N__19000;
    wire N__18995;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18981;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18960;
    wire N__18959;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18899;
    wire N__18898;
    wire N__18897;
    wire N__18894;
    wire N__18893;
    wire N__18890;
    wire N__18889;
    wire N__18888;
    wire N__18887;
    wire N__18884;
    wire N__18883;
    wire N__18882;
    wire N__18877;
    wire N__18874;
    wire N__18871;
    wire N__18868;
    wire N__18865;
    wire N__18860;
    wire N__18855;
    wire N__18854;
    wire N__18845;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18826;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18767;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18740;
    wire N__18739;
    wire N__18738;
    wire N__18733;
    wire N__18730;
    wire N__18729;
    wire N__18726;
    wire N__18721;
    wire N__18720;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18716;
    wire N__18715;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18707;
    wire N__18704;
    wire N__18701;
    wire N__18696;
    wire N__18695;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18669;
    wire N__18668;
    wire N__18667;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18655;
    wire N__18652;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18632;
    wire N__18625;
    wire N__18620;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18537;
    wire N__18536;
    wire N__18533;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18521;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18505;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18482;
    wire N__18481;
    wire N__18480;
    wire N__18479;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18455;
    wire N__18454;
    wire N__18453;
    wire N__18444;
    wire N__18441;
    wire N__18440;
    wire N__18437;
    wire N__18434;
    wire N__18433;
    wire N__18432;
    wire N__18423;
    wire N__18420;
    wire N__18419;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18405;
    wire N__18402;
    wire N__18401;
    wire N__18398;
    wire N__18395;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18287;
    wire N__18286;
    wire N__18283;
    wire N__18282;
    wire N__18281;
    wire N__18276;
    wire N__18273;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18257;
    wire N__18252;
    wire N__18251;
    wire N__18250;
    wire N__18249;
    wire N__18248;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18225;
    wire N__18224;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18216;
    wire N__18215;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18195;
    wire N__18192;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18169;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18154;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18137;
    wire N__18136;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18116;
    wire N__18113;
    wire N__18108;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18077;
    wire N__18076;
    wire N__18073;
    wire N__18068;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17993;
    wire N__17990;
    wire N__17989;
    wire N__17988;
    wire N__17985;
    wire N__17978;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17957;
    wire N__17954;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17931;
    wire N__17928;
    wire N__17927;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17921;
    wire N__17920;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17904;
    wire N__17895;
    wire N__17894;
    wire N__17891;
    wire N__17890;
    wire N__17887;
    wire N__17886;
    wire N__17883;
    wire N__17876;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17858;
    wire N__17853;
    wire N__17852;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17835;
    wire N__17834;
    wire N__17833;
    wire N__17830;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17816;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17806;
    wire N__17799;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17787;
    wire N__17782;
    wire N__17779;
    wire N__17772;
    wire N__17767;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17747;
    wire N__17746;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17722;
    wire N__17717;
    wire N__17714;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17677;
    wire N__17676;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17636;
    wire N__17635;
    wire N__17634;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17620;
    wire N__17617;
    wire N__17616;
    wire N__17615;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17600;
    wire N__17597;
    wire N__17596;
    wire N__17591;
    wire N__17588;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17567;
    wire N__17566;
    wire N__17565;
    wire N__17564;
    wire N__17563;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17540;
    wire N__17537;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17516;
    wire N__17515;
    wire N__17514;
    wire N__17511;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17472;
    wire N__17471;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17463;
    wire N__17462;
    wire N__17461;
    wire N__17460;
    wire N__17457;
    wire N__17452;
    wire N__17447;
    wire N__17442;
    wire N__17437;
    wire N__17430;
    wire N__17429;
    wire N__17428;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17409;
    wire N__17402;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17380;
    wire N__17379;
    wire N__17378;
    wire N__17377;
    wire N__17376;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17362;
    wire N__17355;
    wire N__17346;
    wire N__17343;
    wire N__17342;
    wire N__17339;
    wire N__17338;
    wire N__17337;
    wire N__17336;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17320;
    wire N__17313;
    wire N__17312;
    wire N__17311;
    wire N__17308;
    wire N__17307;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17277;
    wire N__17276;
    wire N__17275;
    wire N__17272;
    wire N__17271;
    wire N__17270;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17256;
    wire N__17251;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17234;
    wire N__17233;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17210;
    wire N__17207;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17195;
    wire N__17194;
    wire N__17193;
    wire N__17192;
    wire N__17185;
    wire N__17180;
    wire N__17177;
    wire N__17176;
    wire N__17171;
    wire N__17168;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17104;
    wire N__17101;
    wire N__17096;
    wire N__17091;
    wire N__17088;
    wire N__17087;
    wire N__17086;
    wire N__17083;
    wire N__17082;
    wire N__17079;
    wire N__17078;
    wire N__17075;
    wire N__17068;
    wire N__17065;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17036;
    wire N__17035;
    wire N__17034;
    wire N__17031;
    wire N__17030;
    wire N__17027;
    wire N__17026;
    wire N__17025;
    wire N__17022;
    wire N__17021;
    wire N__17018;
    wire N__17007;
    wire N__17006;
    wire N__16999;
    wire N__16998;
    wire N__16995;
    wire N__16994;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16975;
    wire N__16972;
    wire N__16967;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16866;
    wire N__16865;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16847;
    wire N__16846;
    wire N__16843;
    wire N__16838;
    wire N__16837;
    wire N__16832;
    wire N__16829;
    wire N__16828;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16769;
    wire N__16768;
    wire N__16767;
    wire N__16766;
    wire N__16765;
    wire N__16764;
    wire N__16763;
    wire N__16762;
    wire N__16761;
    wire N__16750;
    wire N__16745;
    wire N__16738;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16722;
    wire N__16719;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16641;
    wire N__16638;
    wire N__16637;
    wire N__16636;
    wire N__16635;
    wire N__16634;
    wire N__16633;
    wire N__16630;
    wire N__16627;
    wire N__16624;
    wire N__16623;
    wire N__16622;
    wire N__16621;
    wire N__16620;
    wire N__16619;
    wire N__16618;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16595;
    wire N__16590;
    wire N__16587;
    wire N__16582;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16550;
    wire N__16549;
    wire N__16548;
    wire N__16547;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16499;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16481;
    wire N__16480;
    wire N__16479;
    wire N__16478;
    wire N__16475;
    wire N__16474;
    wire N__16471;
    wire N__16460;
    wire N__16457;
    wire N__16452;
    wire N__16451;
    wire N__16450;
    wire N__16449;
    wire N__16446;
    wire N__16445;
    wire N__16444;
    wire N__16441;
    wire N__16440;
    wire N__16437;
    wire N__16436;
    wire N__16433;
    wire N__16418;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16383;
    wire N__16382;
    wire N__16381;
    wire N__16376;
    wire N__16373;
    wire N__16368;
    wire N__16367;
    wire N__16364;
    wire N__16363;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16351;
    wire N__16348;
    wire N__16341;
    wire N__16340;
    wire N__16339;
    wire N__16336;
    wire N__16331;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16316;
    wire N__16313;
    wire N__16310;
    wire N__16307;
    wire N__16304;
    wire N__16301;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16280;
    wire N__16277;
    wire N__16274;
    wire N__16271;
    wire N__16270;
    wire N__16269;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16241;
    wire N__16238;
    wire N__16235;
    wire N__16230;
    wire N__16229;
    wire N__16228;
    wire N__16225;
    wire N__16220;
    wire N__16215;
    wire N__16214;
    wire N__16213;
    wire N__16210;
    wire N__16209;
    wire N__16206;
    wire N__16205;
    wire N__16202;
    wire N__16197;
    wire N__16190;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16175;
    wire N__16172;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16164;
    wire N__16163;
    wire N__16160;
    wire N__16159;
    wire N__16154;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16134;
    wire N__16131;
    wire N__16130;
    wire N__16129;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16109;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16093;
    wire N__16086;
    wire N__16083;
    wire N__16082;
    wire N__16081;
    wire N__16080;
    wire N__16077;
    wire N__16070;
    wire N__16065;
    wire N__16062;
    wire N__16061;
    wire N__16060;
    wire N__16059;
    wire N__16058;
    wire N__16057;
    wire N__16056;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16034;
    wire N__16033;
    wire N__16032;
    wire N__16031;
    wire N__16030;
    wire N__16029;
    wire N__16014;
    wire N__16013;
    wire N__16012;
    wire N__16009;
    wire N__16008;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15977;
    wire N__15972;
    wire N__15969;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15953;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15930;
    wire N__15929;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15919;
    wire N__15914;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15900;
    wire N__15897;
    wire N__15896;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15878;
    wire N__15867;
    wire N__15866;
    wire N__15861;
    wire N__15860;
    wire N__15859;
    wire N__15858;
    wire N__15857;
    wire N__15854;
    wire N__15851;
    wire N__15844;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15824;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15820;
    wire N__15817;
    wire N__15814;
    wire N__15811;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15789;
    wire N__15788;
    wire N__15787;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15776;
    wire N__15773;
    wire N__15772;
    wire N__15765;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15734;
    wire N__15729;
    wire N__15726;
    wire N__15725;
    wire N__15724;
    wire N__15723;
    wire N__15722;
    wire N__15719;
    wire N__15716;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15696;
    wire N__15695;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15680;
    wire N__15679;
    wire N__15678;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15663;
    wire N__15658;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15641;
    wire N__15640;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15629;
    wire N__15626;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15606;
    wire N__15605;
    wire N__15604;
    wire N__15603;
    wire N__15602;
    wire N__15601;
    wire N__15600;
    wire N__15599;
    wire N__15598;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15528;
    wire N__15525;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15517;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15487;
    wire N__15484;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15464;
    wire N__15463;
    wire N__15462;
    wire N__15461;
    wire N__15458;
    wire N__15457;
    wire N__15454;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15429;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15410;
    wire N__15405;
    wire N__15396;
    wire N__15395;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15378;
    wire N__15377;
    wire N__15372;
    wire N__15369;
    wire N__15364;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15350;
    wire N__15345;
    wire N__15344;
    wire N__15343;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15311;
    wire N__15310;
    wire N__15307;
    wire N__15302;
    wire N__15299;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15227;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15215;
    wire N__15214;
    wire N__15211;
    wire N__15206;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15173;
    wire N__15172;
    wire N__15171;
    wire N__15170;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15154;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15140;
    wire N__15139;
    wire N__15136;
    wire N__15131;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15080;
    wire N__15079;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15067;
    wire N__15060;
    wire N__15059;
    wire N__15056;
    wire N__15055;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15048;
    wire N__15039;
    wire N__15036;
    wire N__15035;
    wire N__15032;
    wire N__15031;
    wire N__15030;
    wire N__15027;
    wire N__15026;
    wire N__15025;
    wire N__15024;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15010;
    wire N__15003;
    wire N__14990;
    wire N__14987;
    wire N__14976;
    wire N__14975;
    wire N__14974;
    wire N__14973;
    wire N__14970;
    wire N__14963;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14955;
    wire N__14954;
    wire N__14953;
    wire N__14952;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14945;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14930;
    wire N__14917;
    wire N__14914;
    wire N__14901;
    wire N__14900;
    wire N__14899;
    wire N__14896;
    wire N__14893;
    wire N__14890;
    wire N__14889;
    wire N__14888;
    wire N__14887;
    wire N__14876;
    wire N__14875;
    wire N__14872;
    wire N__14869;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14834;
    wire N__14833;
    wire N__14830;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14798;
    wire N__14795;
    wire N__14794;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14772;
    wire N__14771;
    wire N__14770;
    wire N__14767;
    wire N__14766;
    wire N__14765;
    wire N__14764;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14745;
    wire N__14740;
    wire N__14733;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14716;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14694;
    wire N__14691;
    wire N__14690;
    wire N__14685;
    wire N__14682;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14664;
    wire N__14661;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14636;
    wire N__14635;
    wire N__14632;
    wire N__14627;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14612;
    wire N__14607;
    wire N__14604;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14590;
    wire N__14585;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14568;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14562;
    wire N__14557;
    wire N__14546;
    wire N__14543;
    wire N__14538;
    wire N__14537;
    wire N__14536;
    wire N__14535;
    wire N__14534;
    wire N__14533;
    wire N__14532;
    wire N__14527;
    wire N__14516;
    wire N__14513;
    wire N__14508;
    wire N__14507;
    wire N__14504;
    wire N__14503;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14472;
    wire N__14463;
    wire N__14460;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14448;
    wire N__14445;
    wire N__14444;
    wire N__14443;
    wire N__14438;
    wire N__14435;
    wire N__14430;
    wire N__14427;
    wire N__14424;
    wire N__14423;
    wire N__14422;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14404;
    wire N__14395;
    wire N__14388;
    wire N__14387;
    wire N__14384;
    wire N__14383;
    wire N__14380;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14361;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14273;
    wire N__14272;
    wire N__14271;
    wire N__14268;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14231;
    wire N__14226;
    wire N__14223;
    wire N__14222;
    wire N__14221;
    wire N__14220;
    wire N__14219;
    wire N__14218;
    wire N__14215;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14197;
    wire N__14190;
    wire N__14189;
    wire N__14188;
    wire N__14187;
    wire N__14186;
    wire N__14185;
    wire N__14184;
    wire N__14181;
    wire N__14178;
    wire N__14167;
    wire N__14160;
    wire N__14159;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14147;
    wire N__14146;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14084;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14048;
    wire N__14047;
    wire N__14044;
    wire N__14039;
    wire N__14034;
    wire N__14033;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14023;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14005;
    wire N__14002;
    wire N__13995;
    wire N__13992;
    wire N__13991;
    wire N__13988;
    wire N__13987;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13957;
    wire N__13954;
    wire N__13947;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13937;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13922;
    wire N__13917;
    wire N__13914;
    wire N__13913;
    wire N__13912;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13872;
    wire N__13871;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13863;
    wire N__13862;
    wire N__13861;
    wire N__13858;
    wire N__13857;
    wire N__13846;
    wire N__13841;
    wire N__13838;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13823;
    wire N__13820;
    wire N__13819;
    wire N__13818;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13814;
    wire N__13813;
    wire N__13812;
    wire N__13811;
    wire N__13810;
    wire N__13809;
    wire N__13806;
    wire N__13805;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13791;
    wire N__13784;
    wire N__13775;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13707;
    wire N__13706;
    wire N__13705;
    wire N__13704;
    wire N__13703;
    wire N__13702;
    wire N__13701;
    wire N__13700;
    wire N__13699;
    wire N__13698;
    wire N__13697;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13677;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13657;
    wire N__13650;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13589;
    wire N__13588;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13575;
    wire N__13572;
    wire N__13569;
    wire N__13564;
    wire N__13559;
    wire N__13556;
    wire N__13551;
    wire N__13548;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13495;
    wire N__13494;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13482;
    wire N__13479;
    wire N__13478;
    wire N__13477;
    wire N__13476;
    wire N__13475;
    wire N__13468;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13452;
    wire N__13443;
    wire N__13442;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13432;
    wire N__13431;
    wire N__13428;
    wire N__13425;
    wire N__13424;
    wire N__13421;
    wire N__13420;
    wire N__13417;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13401;
    wire N__13398;
    wire N__13389;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13381;
    wire N__13380;
    wire N__13379;
    wire N__13378;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13359;
    wire N__13350;
    wire N__13347;
    wire N__13346;
    wire N__13343;
    wire N__13342;
    wire N__13339;
    wire N__13338;
    wire N__13337;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13323;
    wire N__13322;
    wire N__13321;
    wire N__13320;
    wire N__13319;
    wire N__13314;
    wire N__13313;
    wire N__13312;
    wire N__13311;
    wire N__13308;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13287;
    wire N__13284;
    wire N__13277;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13250;
    wire N__13247;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13226;
    wire N__13221;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13172;
    wire N__13171;
    wire N__13170;
    wire N__13169;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13155;
    wire N__13152;
    wire N__13151;
    wire N__13150;
    wire N__13145;
    wire N__13140;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13120;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13113;
    wire N__13110;
    wire N__13101;
    wire N__13096;
    wire N__13093;
    wire N__13088;
    wire N__13079;
    wire N__13074;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13043;
    wire N__13038;
    wire N__13037;
    wire N__13036;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13030;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13008;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12987;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12962;
    wire N__12961;
    wire N__12960;
    wire N__12957;
    wire N__12950;
    wire N__12947;
    wire N__12942;
    wire N__12941;
    wire N__12940;
    wire N__12939;
    wire N__12936;
    wire N__12929;
    wire N__12924;
    wire N__12921;
    wire N__12920;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12880;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12864;
    wire N__12861;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12843;
    wire N__12842;
    wire N__12841;
    wire N__12838;
    wire N__12833;
    wire N__12830;
    wire N__12825;
    wire N__12822;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12791;
    wire N__12788;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12776;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12764;
    wire N__12759;
    wire N__12756;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12728;
    wire N__12727;
    wire N__12726;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12712;
    wire N__12709;
    wire N__12704;
    wire N__12699;
    wire N__12698;
    wire N__12697;
    wire N__12696;
    wire N__12695;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12687;
    wire N__12686;
    wire N__12685;
    wire N__12682;
    wire N__12681;
    wire N__12676;
    wire N__12669;
    wire N__12668;
    wire N__12667;
    wire N__12666;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12648;
    wire N__12641;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12615;
    wire N__12608;
    wire N__12603;
    wire N__12602;
    wire N__12601;
    wire N__12600;
    wire N__12599;
    wire N__12598;
    wire N__12597;
    wire N__12596;
    wire N__12591;
    wire N__12586;
    wire N__12579;
    wire N__12576;
    wire N__12575;
    wire N__12574;
    wire N__12573;
    wire N__12572;
    wire N__12571;
    wire N__12570;
    wire N__12569;
    wire N__12568;
    wire N__12561;
    wire N__12558;
    wire N__12549;
    wire N__12540;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12522;
    wire N__12521;
    wire N__12520;
    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12514;
    wire N__12513;
    wire N__12512;
    wire N__12511;
    wire N__12508;
    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12504;
    wire N__12503;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12493;
    wire N__12492;
    wire N__12485;
    wire N__12482;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12442;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12407;
    wire N__12400;
    wire N__12395;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12377;
    wire N__12376;
    wire N__12373;
    wire N__12368;
    wire N__12365;
    wire N__12360;
    wire N__12357;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12337;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12321;
    wire N__12320;
    wire N__12319;
    wire N__12318;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12312;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12292;
    wire N__12285;
    wire N__12284;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12280;
    wire N__12277;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12243;
    wire N__12240;
    wire N__12239;
    wire N__12238;
    wire N__12235;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12199;
    wire N__12198;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12170;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12128;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12120;
    wire N__12119;
    wire N__12116;
    wire N__12107;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12017;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__12000;
    wire N__11999;
    wire N__11998;
    wire N__11997;
    wire N__11996;
    wire N__11993;
    wire N__11992;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11968;
    wire N__11959;
    wire N__11954;
    wire N__11951;
    wire N__11946;
    wire N__11931;
    wire N__11930;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11921;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11905;
    wire N__11902;
    wire N__11895;
    wire N__11894;
    wire N__11893;
    wire N__11890;
    wire N__11889;
    wire N__11888;
    wire N__11887;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11870;
    wire N__11861;
    wire N__11860;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11839;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11814;
    wire N__11813;
    wire N__11812;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11793;
    wire N__11788;
    wire N__11781;
    wire N__11780;
    wire N__11779;
    wire N__11776;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11768;
    wire N__11765;
    wire N__11758;
    wire N__11755;
    wire N__11754;
    wire N__11749;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11733;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11718;
    wire N__11717;
    wire N__11714;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11710;
    wire N__11709;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11704;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11690;
    wire N__11685;
    wire N__11680;
    wire N__11675;
    wire N__11670;
    wire N__11667;
    wire N__11662;
    wire N__11653;
    wire N__11650;
    wire N__11645;
    wire N__11640;
    wire N__11635;
    wire N__11632;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11603;
    wire N__11600;
    wire N__11599;
    wire N__11594;
    wire N__11591;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11576;
    wire N__11575;
    wire N__11572;
    wire N__11567;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11433;
    wire N__11430;
    wire N__11417;
    wire N__11412;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11406;
    wire N__11403;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11392;
    wire N__11391;
    wire N__11388;
    wire N__11375;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11354;
    wire N__11353;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11330;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11318;
    wire N__11317;
    wire N__11316;
    wire N__11315;
    wire N__11314;
    wire N__11313;
    wire N__11310;
    wire N__11297;
    wire N__11292;
    wire N__11291;
    wire N__11290;
    wire N__11289;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11277;
    wire N__11274;
    wire N__11269;
    wire N__11258;
    wire N__11253;
    wire N__11252;
    wire N__11251;
    wire N__11248;
    wire N__11247;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11230;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11216;
    wire N__11215;
    wire N__11214;
    wire N__11213;
    wire N__11212;
    wire N__11209;
    wire N__11208;
    wire N__11197;
    wire N__11192;
    wire N__11189;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11168;
    wire N__11167;
    wire N__11166;
    wire N__11165;
    wire N__11164;
    wire N__11151;
    wire N__11148;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11136;
    wire N__11135;
    wire N__11134;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11081;
    wire N__11080;
    wire N__11077;
    wire N__11072;
    wire N__11067;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11057;
    wire N__11056;
    wire N__11051;
    wire N__11046;
    wire N__11041;
    wire N__11036;
    wire N__11031;
    wire N__11028;
    wire N__11027;
    wire N__11026;
    wire N__11019;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11008;
    wire N__11007;
    wire N__11004;
    wire N__10993;
    wire N__10990;
    wire N__10985;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10968;
    wire N__10959;
    wire N__10956;
    wire N__10953;
    wire N__10948;
    wire N__10941;
    wire N__10940;
    wire N__10937;
    wire N__10936;
    wire N__10935;
    wire N__10934;
    wire N__10929;
    wire N__10924;
    wire N__10921;
    wire N__10916;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10908;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10845;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10825;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10802;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10784;
    wire N__10779;
    wire N__10778;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10755;
    wire N__10752;
    wire N__10751;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10739;
    wire N__10738;
    wire N__10737;
    wire N__10736;
    wire N__10735;
    wire N__10730;
    wire N__10727;
    wire N__10720;
    wire N__10717;
    wire N__10710;
    wire N__10709;
    wire N__10708;
    wire N__10705;
    wire N__10704;
    wire N__10701;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10652;
    wire N__10651;
    wire N__10648;
    wire N__10643;
    wire N__10638;
    wire N__10635;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10586;
    wire N__10585;
    wire N__10584;
    wire N__10583;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10554;
    wire N__10553;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10535;
    wire N__10532;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10512;
    wire N__10509;
    wire N__10506;
    wire N__10503;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10479;
    wire N__10476;
    wire N__10473;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10458;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10421;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10389;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10184;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10172;
    wire N__10169;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10146;
    wire N__10145;
    wire N__10144;
    wire N__10141;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10131;
    wire N__10128;
    wire N__10123;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9941;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9912;
    wire N__9903;
    wire N__9900;
    wire N__9899;
    wire N__9898;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9886;
    wire N__9879;
    wire N__9876;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9872;
    wire N__9869;
    wire N__9860;
    wire N__9855;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9837;
    wire N__9834;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9794;
    wire N__9793;
    wire N__9792;
    wire N__9791;
    wire N__9788;
    wire N__9779;
    wire N__9774;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9768;
    wire N__9765;
    wire N__9764;
    wire N__9761;
    wire N__9756;
    wire N__9753;
    wire N__9748;
    wire N__9741;
    wire N__9738;
    wire N__9735;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9704;
    wire N__9701;
    wire N__9700;
    wire N__9699;
    wire N__9696;
    wire N__9689;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9608;
    wire N__9605;
    wire N__9604;
    wire N__9603;
    wire N__9600;
    wire N__9595;
    wire N__9592;
    wire N__9585;
    wire N__9584;
    wire N__9581;
    wire N__9580;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9486;
    wire N__9485;
    wire N__9484;
    wire N__9481;
    wire N__9476;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9464;
    wire N__9461;
    wire N__9460;
    wire N__9457;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9445;
    wire N__9438;
    wire N__9435;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9412;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9392;
    wire N__9387;
    wire N__9382;
    wire N__9375;
    wire N__9372;
    wire N__9371;
    wire N__9368;
    wire N__9367;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9361;
    wire N__9358;
    wire N__9351;
    wire N__9346;
    wire N__9339;
    wire N__9338;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9320;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9288;
    wire N__9287;
    wire N__9286;
    wire N__9285;
    wire N__9282;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9262;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9254;
    wire N__9245;
    wire N__9236;
    wire N__9231;
    wire N__9230;
    wire N__9229;
    wire N__9228;
    wire N__9227;
    wire N__9226;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9203;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9171;
    wire N__9170;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9146;
    wire N__9143;
    wire N__9140;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9129;
    wire N__9122;
    wire N__9117;
    wire N__9116;
    wire N__9115;
    wire N__9114;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9098;
    wire N__9097;
    wire N__9096;
    wire N__9093;
    wire N__9088;
    wire N__9085;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9065;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9050;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9042;
    wire N__9039;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9021;
    wire N__9020;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9004;
    wire N__8997;
    wire N__8994;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8986;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8970;
    wire N__8967;
    wire N__8966;
    wire N__8965;
    wire N__8964;
    wire N__8963;
    wire N__8958;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8925;
    wire N__8922;
    wire N__8915;
    wire N__8912;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8894;
    wire N__8893;
    wire N__8892;
    wire N__8889;
    wire N__8884;
    wire N__8881;
    wire N__8874;
    wire N__8873;
    wire N__8872;
    wire N__8869;
    wire N__8864;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8842;
    wire N__8837;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8821;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8809;
    wire N__8806;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8792;
    wire N__8789;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8746;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8732;
    wire N__8731;
    wire N__8730;
    wire N__8729;
    wire N__8720;
    wire N__8717;
    wire N__8712;
    wire N__8711;
    wire N__8710;
    wire N__8707;
    wire N__8706;
    wire N__8699;
    wire N__8696;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8662;
    wire N__8655;
    wire N__8652;
    wire N__8651;
    wire N__8650;
    wire N__8647;
    wire N__8644;
    wire N__8637;
    wire N__8634;
    wire N__8633;
    wire N__8632;
    wire N__8631;
    wire N__8630;
    wire N__8619;
    wire N__8616;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8594;
    wire N__8593;
    wire N__8592;
    wire N__8591;
    wire N__8590;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8561;
    wire N__8560;
    wire N__8557;
    wire N__8556;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8539;
    wire N__8532;
    wire N__8531;
    wire N__8530;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8519;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8507;
    wire N__8502;
    wire N__8493;
    wire N__8490;
    wire N__8489;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8474;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8464;
    wire N__8457;
    wire N__8456;
    wire N__8455;
    wire N__8452;
    wire N__8447;
    wire N__8444;
    wire N__8439;
    wire N__8438;
    wire N__8437;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8416;
    wire N__8415;
    wire N__8414;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8370;
    wire N__8367;
    wire N__8366;
    wire N__8365;
    wire N__8364;
    wire N__8363;
    wire N__8358;
    wire N__8351;
    wire N__8346;
    wire N__8345;
    wire N__8344;
    wire N__8343;
    wire N__8342;
    wire N__8337;
    wire N__8330;
    wire N__8325;
    wire N__8324;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8312;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8294;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8280;
    wire N__8277;
    wire N__8276;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8238;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.vbuf_count.un328_ci_3_cascade_ ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.un350_ci ;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_2_2 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_5 ;
    wire uart_RXD;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.un284_ci ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un44_ci_cascade_ ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.un88_ci_3 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un44_ci ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un220_ci ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un4_l_count_11 ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.un4_l_count_16_cascade_ ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.un143_ci_0 ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un66_ci ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.un110_ci ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu2.trig_rd_is_det_cascade_ ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.un404_ci_cascade_ ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.mem0.N_76_i ;
    wire \uu2.mem0.N_73_i ;
    wire \uu2.mem0.N_79_i ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu0.sec_clkDZ0 ;
    wire oneSecStrb_cascade_;
    wire \uu2.N_118_cascade_ ;
    wire \uu2.N_117 ;
    wire \uu2.N_117_cascade_ ;
    wire \INVuu2.w_addr_user_nesr_7C_net ;
    wire \uu2.mem0.N_75_i ;
    wire \uu2.mem0.N_74_i ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.N_186 ;
    wire \uu2.w_addr_user_3_i_a2_2_6 ;
    wire \uu2.N_150_cascade_ ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.N_115_cascade_ ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.un28_w_addr_user_i_0_0 ;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.mem0.N_78_i ;
    wire \uu2.mem0.N_77_i ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire vbuf_tx_data_5;
    wire \uu2.r_data_wire_6 ;
    wire vbuf_tx_data_6;
    wire \uu2.r_data_wire_7 ;
    wire vbuf_tx_data_7;
    wire \INVuu2.r_data_reg_0C_net ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.un165_ci_0 ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmap_RNIAE522Z0Z_93_cascade_ ;
    wire \INVuu2.bitmap_215C_net ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.bitmap_RNIKL222Z0Z_212_cascade_ ;
    wire \uu2.bitmap_pmux_27_ns_1 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \Lab_UT.sec1_3 ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmap_pmux_24_i_m2_am_1 ;
    wire \uu2.un51_w_data_displaying_cascade_ ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.w_addr_displaying_4_1 ;
    wire \uu2.un51_w_data_displaying ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i5_mux_cascade_ ;
    wire \uu2.N_404 ;
    wire \uu2.bitmap_pmux_29_0_cascade_ ;
    wire \uu2.bitmap_pmux ;
    wire \INVuu2.bitmap_40C_net ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmap_RNI1PH82Z0Z_40_cascade_ ;
    wire \uu2.N_401_cascade_ ;
    wire \uu2.N_406 ;
    wire \uu2.un31_w_data_displaying_1 ;
    wire \uu2.un49_w_data_displaying_1 ;
    wire \uu2.mem0.N_81_i ;
    wire \uu2.mem0.N_80_i ;
    wire \uu2.mem0.N_72_i ;
    wire \uu2.N_111_cascade_ ;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.mem0.w_data_i_a2_1_0_cascade_ ;
    wire \uu2.mem0.N_82_i ;
    wire \uu2.mem0.N_110 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.N_225 ;
    wire \uu2.N_144_cascade_ ;
    wire \uu2.N_361 ;
    wire \uu2.mem0.w_data_0_a2_0_4_cascade_ ;
    wire \uu2.mem0.w_data_4 ;
    wire L3_tx_data_5;
    wire L3_tx_data_4;
    wire \uu2.N_109 ;
    wire \uu2.N_111 ;
    wire \uu2.N_109_cascade_ ;
    wire L3_tx_data_rdy;
    wire \Lab_UT.dispString.N_61 ;
    wire \Lab_UT.dispString.un46_dOutP_i_m_3 ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_3_cascade_ ;
    wire \Lab_UT.dispString.dOutP_6 ;
    wire L3_tx_data_3;
    wire \Lab_UT.dispString.N_50 ;
    wire \Lab_UT.dispString.N_28_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_3 ;
    wire \buart.Z_tx.un1_bitcount_c3_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.un1_bitcount_c2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire vbuf_tx_data_rdy;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.bitmap_pmux_25_bm_1 ;
    wire \Lab_UT.sec2_3 ;
    wire \Lab_UT.sec2_2 ;
    wire \Lab_UT.sec2_1 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \uu2.N_216_cascade_ ;
    wire \Lab_UT.sec1_1 ;
    wire \Lab_UT.sec1_2 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.bitmap_pmux_24_i_m2_bm_1_cascade_ ;
    wire \uu2.bitmap_RNI1UT12Z0Z_75 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \Lab_UT.min2_2 ;
    wire \Lab_UT.min2_1 ;
    wire \Lab_UT.min2_3 ;
    wire \Lab_UT.min2_0 ;
    wire \INVuu2.bitmap_296C_net ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.un437_ci_0_cascade_ ;
    wire \INVuu2.bitmap_69C_net ;
    wire L3_tx_data_6;
    wire \uu2.mem0.w_data_6 ;
    wire \INVuu2.w_addr_displaying_8C_net ;
    wire \uu2.un31_w_data_displaying_2 ;
    wire \uu2.un33_w_data_displaying ;
    wire \uu2.w_addr_i_0_tzZ0Z_0 ;
    wire \uu2.un21_w_addr_displaying_i_cascade_ ;
    wire \INVuu2.w_addr_displaying_nesr_3C_net ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.bitmap_pmux_sn_N_65 ;
    wire \uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.bitmap_pmux_sn_i7_mux_0 ;
    wire \uu2.un15_w_data_displaying_2 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.N_383_cascade_ ;
    wire \uu2.N_215 ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_ ;
    wire \uu2.bitmap_RNIS4UH1Z0Z_314 ;
    wire \uu2.N_397 ;
    wire \uu2.bitmap_pmux_sn_N_15 ;
    wire \uu2.bitmap_pmux_sn_N_54_mux_cascade_ ;
    wire \uu2.bitmap_RNIELSJ2Z0Z_111 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.un21_w_addr_displaying_i ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.N_115 ;
    wire \uu2.N_144 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire o_One_Sec_Pulse;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_2C_net ;
    wire \Lab_UT.dispString.dOutP_1_iv_0_4 ;
    wire \Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ;
    wire L3_tx_data_1;
    wire \Lab_UT.dispString.dOutP_0_iv_0_5 ;
    wire \Lab_UT.dispString.N_41_cascade_ ;
    wire \Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_ ;
    wire \Lab_UT.dispString.dOut_RNO_0Z0Z_0 ;
    wire L3_tx_data_0;
    wire \Lab_UT.alarmchar_1 ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_ ;
    wire \Lab_UT.dispString.dOut_RNO_0Z0Z_2 ;
    wire L3_tx_data_2;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.N_32 ;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire \Lab_UT.dispString.dOut_RNO_0Z0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_5_14_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_3_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_2_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.didp.un2_did_alarmMatch_0_cascade_ ;
    wire \Lab_UT.sec2_0 ;
    wire \Lab_UT.loadalarm_0_0_cascade_ ;
    wire \Lab_UT.sec1_0 ;
    wire \Lab_UT.didp.did_alarmMatch_7 ;
    wire \uu2.un15_w_data_displaying_5 ;
    wire \uu2.o_adder_vbuf_w_addr_displaying_6_cascade_ ;
    wire \INVuu2.w_addr_displaying_ness_6C_net ;
    wire \uu2.un21_w_addr_displaying_i_0 ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.un15_w_data_displaying_6 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.bitmap_pmux_sn_N_36 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmap_pmux_25_am_1 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.bitmap_RNIV8902Z0Z_66 ;
    wire \Lab_UT.min1_2 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmap_pmux_26_bm_1 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \uu2.N_217 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_11 ;
    wire \Lab_UT.didp.countrce4.q_5_2_cascade_ ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_ ;
    wire \Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i ;
    wire \Lab_UT.dictrl.alarmstate_0_sqmuxa_1 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_0_i_0 ;
    wire \Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_0 ;
    wire \Lab_UT.dictrl.N_127_0_0 ;
    wire \Lab_UT.trig ;
    wire \Lab_UT.dictrl.N_127_0_0_cascade_ ;
    wire \Lab_UT.dictrl.justentered_0 ;
    wire \Lab_UT.shifter_ret_3_RNIK5FS8_0 ;
    wire \Lab_UT.shifter_ret_3_RNIQBH29_0 ;
    wire \Lab_UT.armed ;
    wire \Lab_UT.armed_cascade_ ;
    wire \Lab_UT.alarmMatch ;
    wire G_203;
    wire \Lab_UT.dictrl.alarmstate8_2_reti ;
    wire \Lab_UT.dictrl.alarmstate8_10_3_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate8 ;
    wire bu_rx_data_7;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_6 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_0_7 ;
    wire bu_rx_data_i_4_fast_3;
    wire buart__rx_shifter_ret_5_fast;
    wire \Lab_UT.dictrl.g1_1Z0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.N_98_mux_1 ;
    wire \Lab_UT.dictrl.N_98_mux_0_0 ;
    wire \Lab_UT.dictrl.g0_3_1_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_1_cascade_ ;
    wire \Lab_UT.didp.countrce1.un13_qPone ;
    wire \Lab_UT.didp.un1_dicLdSones_0 ;
    wire \Lab_UT.didp.un1_dicLdSones_0_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_2 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.didp.did_alarmMatch_5 ;
    wire \Lab_UT.didp.un1_dicLdMones_0_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_1 ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.min1_0 ;
    wire \Lab_UT.min1_1 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.didp.did_alarmMatch_3 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_ ;
    wire \Lab_UT.didp.did_alarmMatch_1 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_12 ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.loadalarm_1 ;
    wire \Lab_UT.loadalarm_0_0 ;
    wire \Lab_UT.min1_3 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.dicRun_2 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.didp.countrce4.un13_qPone ;
    wire \Lab_UT.didp.countrce4.q_5_0_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_0 ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.didp.countrce4.un20_qPone ;
    wire \Lab_UT.didp.countrce4.q_5_3_cascade_ ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.un1_dicLdMtens_0 ;
    wire \Lab_UT.dictrl.N_116_mux_0_cascade_ ;
    wire \Lab_UT.dictrl.N_116_mux_0_0_0 ;
    wire \Lab_UT.dictrl.N_1304_0_1_0_cascade_ ;
    wire \Lab_UT.dictrl.N_1304_0 ;
    wire \Lab_UT.dictrl.N_1304_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_88_0_0 ;
    wire \Lab_UT.dictrl.g1_1_1_cascade_ ;
    wire \Lab_UT.dictrl.g1_0 ;
    wire \Lab_UT.dictrl.m25_xZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.N_116_mux_cascade_ ;
    wire \Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_0_a3_4 ;
    wire \Lab_UT.dictrl.N_98_mux_4_cascade_ ;
    wire \Lab_UT.dictrl.g1_1_1_0 ;
    wire bu_rx_data_fast_4;
    wire \Lab_UT.dictrl.N_98_mux_0 ;
    wire \Lab_UT.dictrl.g0_3_1_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_4Z0Z_1 ;
    wire buart__rx_shifter_ret_1_fast;
    wire \Lab_UT.dictrl.N_20_0 ;
    wire \Lab_UT.dictrl.g0_5_2 ;
    wire bu_rx_data_i_4_fast_7;
    wire buart__rx_sample_g;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.didp.did_alarmMatch_2 ;
    wire \Lab_UT.didp.di_Sones_1 ;
    wire \Lab_UT.didp.di_Sones_3 ;
    wire \Lab_UT.didp.di_Sones_2 ;
    wire \Lab_UT.didp.di_Mones_1 ;
    wire \Lab_UT.didp.di_Mones_0 ;
    wire \Lab_UT.didp.countrce3.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_2_cascade_ ;
    wire \Lab_UT.didp.countrce3.un13_qPone ;
    wire \Lab_UT.didp.di_Mones_2 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_3_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdMones_0 ;
    wire \Lab_UT.didp.di_Mones_3 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.ce_12_2_3 ;
    wire \Lab_UT.didp.un24_ce_2 ;
    wire \Lab_UT.didp.reset_12_1_3 ;
    wire \Lab_UT.didp.di_Mtens_1 ;
    wire \Lab_UT.didp.ce_12_3_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_3 ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.un18_ce ;
    wire oneSecStrb;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \resetGen.un241_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_count_2_0_4_cascade_ ;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \Lab_UT.dicRun_1 ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.un252_ci ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un11_l_count_i ;
    wire \Lab_UT.dicLdASones_0 ;
    wire \Lab_UT.dictrl.g3_1 ;
    wire \Lab_UT.dictrl.i9_mux_0_cascade_ ;
    wire \Lab_UT.dictrl.N_2000_0_cascade_ ;
    wire \Lab_UT.dictrl.state_i_4_2 ;
    wire \Lab_UT.dicLdAMones_2 ;
    wire \Lab_UT.dictrl.N_94_0 ;
    wire \Lab_UT.dictrl.N_2000_0 ;
    wire \Lab_UT.dictrl.g1 ;
    wire \Lab_UT.dictrl.g1_3_1 ;
    wire \Lab_UT.dictrl.N_88_0 ;
    wire \Lab_UT.dictrl.g1Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.i9_mux_0_1_0_cascade_ ;
    wire \Lab_UT.dictrl.N_94_0_1_0 ;
    wire \Lab_UT.dictrl.N_2000_0_1_0_cascade_ ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_ ;
    wire \Lab_UT.dictrl.N_96_1_cascade_ ;
    wire \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3 ;
    wire \Lab_UT.dictrl.m36_0 ;
    wire \Lab_UT.dictrl.g1_5_0 ;
    wire \Lab_UT.dictrl.m45_1 ;
    wire \Lab_UT.dictrl.m25Z0Z_0 ;
    wire \Lab_UT.dictrl.N_6_0 ;
    wire \Lab_UT.dictrl.N_5 ;
    wire \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ;
    wire \Lab_UT.dictrl.state_fast_0 ;
    wire bu_rx_data_i_4_0;
    wire \Lab_UT.dictrl.g1_5 ;
    wire \Lab_UT.dictrl.g0_5_4 ;
    wire \Lab_UT.dicLdMones_1 ;
    wire \Lab_UT.dictrl.N_1300_0_cascade_ ;
    wire \Lab_UT.dictrl.g1_2_0 ;
    wire \Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_ ;
    wire buart__rx_shifter_0_fast_2;
    wire \Lab_UT.dictrl.g0_5_5 ;
    wire \Lab_UT.dictrl.N_7 ;
    wire \Lab_UT.dictrl.g0_4_a4_4 ;
    wire \Lab_UT.dictrl.N_5_2 ;
    wire buart__rx_shifter_0_fast_3;
    wire bu_rx_data_5_rep1;
    wire bu_rx_data_4_rep1;
    wire bu_rx_data_fast_5;
    wire bu_rx_data_i_4_7_rep1;
    wire \Lab_UT.dictrl.g0_28_1Z0Z_0 ;
    wire bu_rx_data_fast_6;
    wire \Lab_UT.dictrl.m31_xZ0Z0 ;
    wire bu_rx_data_6_rep1;
    wire \Lab_UT.dictrl.g0_43_xZ0 ;
    wire \Lab_UT.dictrl.N_84_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate8_2 ;
    wire \Lab_UT.dictrl.g1_0_0_0_0 ;
    wire \Lab_UT.dictrl.g0_4_a4Z0Z_5 ;
    wire \Lab_UT.didp.countrce2.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce2.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce2.q_5_3_cascade_ ;
    wire \Lab_UT.didp.di_Stens_3 ;
    wire \Lab_UT.didp.countrce2.q_5_0 ;
    wire bu_rx_data_2;
    wire \Lab_UT.didp.countrce2.un13_qPone ;
    wire \Lab_UT.didp.countrce2.q_5_2_cascade_ ;
    wire \Lab_UT.didp.di_Stens_2 ;
    wire \Lab_UT.didp.di_Stens_0 ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.didp.countrce2.q_5_1_cascade_ ;
    wire \Lab_UT.didp.di_Stens_1 ;
    wire \Lab_UT.LdStens ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.LdStens_i_4 ;
    wire \Lab_UT.didp.un1_dicLdStens_0 ;
    wire \Lab_UT.LdSones ;
    wire \Lab_UT.didp.di_Sones_0 ;
    wire \Lab_UT.didp.countrce1.q_5_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2 ;
    wire \Lab_UT.LdSones_i_4 ;
    wire bfn_9_5_0_;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \Lab_UT.dictrl.state_i_4_0 ;
    wire \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.state_i_4_1 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2 ;
    wire \Lab_UT.dictrl.dicLdStens_1 ;
    wire \Lab_UT.dictrl.N_101_cascade_ ;
    wire \Lab_UT.dictrl.N_5_0 ;
    wire \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.state_fast_3 ;
    wire \Lab_UT.dictrl.state_3_rep1 ;
    wire bu_rx_data_rdy_0_g;
    wire bu_rx_data_0;
    wire \Lab_UT.dictrl.g0_9Z0Z_1 ;
    wire \Lab_UT.dictrl.m25Z0Z_4 ;
    wire \Lab_UT.dictrl.N_116_mux_1_cascade_ ;
    wire \Lab_UT.dictrl.N_120_0_cascade_ ;
    wire \Lab_UT.dictrl.N_1302_0 ;
    wire \Lab_UT.dictrl.N_119_0 ;
    wire \Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0 ;
    wire \Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0 ;
    wire \Lab_UT.dictrl.N_120 ;
    wire \Lab_UT.dictrl.N_99 ;
    wire \Lab_UT.dictrl.N_96 ;
    wire \Lab_UT.dictrl.N_99_cascade_ ;
    wire \Lab_UT.dictrl.N_101 ;
    wire \Lab_UT.dictrl.N_100_cascade_ ;
    wire \Lab_UT.dictrl.next_state_0_1 ;
    wire \Lab_UT.dictrl.N_104_cascade_ ;
    wire \Lab_UT.dictrl.N_99_0_cascade_ ;
    wire \Lab_UT.dictrl.N_96_0_0 ;
    wire \Lab_UT.dictrl.g2 ;
    wire \Lab_UT.dictrl.g0_0_0_a3_5 ;
    wire \Lab_UT.dictrl.N_98_mux_2 ;
    wire bu_rx_data_i_4_5;
    wire \resetGen.escKeyZ0Z_4 ;
    wire \resetGen.escKeyZ0Z_5_cascade_ ;
    wire \resetGen.escKeyZ0 ;
    wire \Lab_UT.dictrl.g1_0_0_0 ;
    wire \Lab_UT.dictrl.N_88_2 ;
    wire bu_rx_data_i_4_3;
    wire \Lab_UT.dictrl.N_95_0_cascade_ ;
    wire \Lab_UT.dictrl.N_103_0 ;
    wire \Lab_UT.dictrl.g1_2_1_0 ;
    wire \Lab_UT.dictrl.g1_3 ;
    wire \Lab_UT.dictrl.N_88 ;
    wire \Lab_UT.dictrl.N_95 ;
    wire \Lab_UT.dictrl.N_103 ;
    wire bu_rx_data_3;
    wire \Lab_UT.dictrl.m63_0Z0Z_1 ;
    wire \Lab_UT.dictrl.N_95_0_0_1 ;
    wire \Lab_UT.dictrl.N_98_mux ;
    wire \Lab_UT.dictrl.N_84 ;
    wire \Lab_UT.dictrl.N_89 ;
    wire \Lab_UT.dictrl.m68_1 ;
    wire \Lab_UT.dictrl.N_89_cascade_ ;
    wire \Lab_UT.dictrl.N_99_mux ;
    wire \Lab_UT.dictrl.N_102 ;
    wire \Lab_UT.dictrl.g1_1Z0Z_0 ;
    wire \Lab_UT.dictrl.g1_2Z0Z_1 ;
    wire \Lab_UT.dictrl.N_102_0 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire buart__rx_ser_clk_cascade_;
    wire \Lab_UT.dictrl.N_83 ;
    wire \Lab_UT.dictrl.N_194_cascade_ ;
    wire buart__rx_sample;
    wire buart__rx_bitcount_2;
    wire buart__rx_bitcount_1;
    wire buart__rx_bitcount_4;
    wire m89_bm;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire buart__rx_N_27_0_i_cascade_;
    wire \Lab_UT.dictrl.N_107_mux_cascade_ ;
    wire m89_am;
    wire buart__rx_hh_0;
    wire buart__rx_hh_1;
    wire \Lab_UT.dictrl.N_102_mux ;
    wire buart__rx_N_27_0_i;
    wire buart__rx_startbit_cascade_;
    wire buart__rx_bitcount_0;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \Lab_UT.dictrl.i9_mux_0_0 ;
    wire \Lab_UT.dictrl.N_94_0_0 ;
    wire \Lab_UT.dictrl.N_2000_0_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3 ;
    wire \Lab_UT.dictrl.N_121_mux ;
    wire Lab_UT_dictrl_next_state_3_cascade_;
    wire \Lab_UT.dictrl.state_ret_12_RNOZ0Z_3 ;
    wire \Lab_UT.dictrl.next_state_0_0_2 ;
    wire \Lab_UT.dictrl.state_ret_12_RNOZ0Z_4 ;
    wire \Lab_UT.dictrl.state_ret_12and_a0_1 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0 ;
    wire \Lab_UT.dictrl.state_ret_12and_0_0_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1 ;
    wire \Lab_UT.dictrl.state_3_rep2 ;
    wire buart__rx_bitcount_3;
    wire buart__rx_valid_3;
    wire Lab_UT_dictrl_next_state_3;
    wire bu_rx_data_rdy_cascade_;
    wire rst;
    wire \Lab_UT.dictrl.N_119_mux ;
    wire \Lab_UT.dictrl.i9_mux_cascade_ ;
    wire \Lab_UT.dictrl.N_94 ;
    wire \Lab_UT.dictrl.next_state_0_2 ;
    wire \Lab_UT.dictrl.N_90 ;
    wire \Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.N_119 ;
    wire \Lab_UT.dictrl.N_139_cascade_ ;
    wire \Lab_UT.dictrl.N_116_mux ;
    wire \Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ;
    wire \Lab_UT.dictrl.g2_2 ;
    wire \Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1 ;
    wire \Lab_UT.dictrl.N_5_1 ;
    wire \Lab_UT.dictrl.g2_0_0_0_0 ;
    wire \Lab_UT.dictrl.stateZ0Z_3 ;
    wire \Lab_UT.dictrl.N_103_0_0_0 ;
    wire \Lab_UT.dictrl.N_1302_1_0_0 ;
    wire \Lab_UT.dictrl.N_119_0_0_0_cascade_ ;
    wire \Lab_UT.dictrl.stateZ0Z_2 ;
    wire \Lab_UT.dictrl.g1Z0Z_4 ;
    wire \Lab_UT.dictrl.stateZ0Z_0 ;
    wire \Lab_UT.dictrl.m46_i_0_a5_1 ;
    wire \Lab_UT.dictrl.N_86 ;
    wire \Lab_UT.dictrl.N_8 ;
    wire \Lab_UT.dictrl.next_state_0_0 ;
    wire Lab_UT_dictrl_un1_next_state66_0;
    wire \Lab_UT.dictrl.m46_i_0_0_0 ;
    wire bu_rx_data_i_3_1;
    wire bu_rx_data_i_4_7;
    wire bu_rx_data_6;
    wire bu_rx_data_i_4_4;
    wire \Lab_UT.dictrl.stateZ0Z_1 ;
    wire g0_3_4_cascade_;
    wire g0_3_5;
    wire \Lab_UT.dictrl.g1Z0Z_2 ;
    wire N_12;
    wire \Lab_UT.dictrl.state_0_rep1 ;
    wire bu_rx_data_4;
    wire \Lab_UT.dictrl.N_13 ;
    wire bu_rx_data_5;
    wire bu_rx_data_1;
    wire bu_rx_data_i_4_3_rep1;
    wire bu_rx_data_i_4_2;
    wire m46_i_0_a3_2;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_12_3_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire buart__rx_ser_clk;
    wire buart__rx_startbit;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.dictrl.next_state_0_3 ;
    wire clk_g;
    wire bu_rx_data_rdy;
    wire rst_g;
    wire bu_rx_data_rdy_0;
    wire \resetGen.r_m3_i_a3_0_2 ;
    wire N_6;
    wire Lab_UT_dictrl_next_state_0_1_2;
    wire Lab_UT_dictrl_next_state_0_0_0;
    wire rst_RNIAL6V33;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__8217),
            .RESETB(N__22914),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__9186,N__9489,N__9465,N__9855,N__9942,N__9339,N__9438,N__9405,N__9375}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__9300,N__9624,N__9639,N__9309,N__9666,N__9684,N__9549,N__10467,N__10479}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__11514,dangling_wire_31,N__10341,dangling_wire_32,N__10815,dangling_wire_33,N__10311,dangling_wire_34,N__10452,dangling_wire_35,N__10305,dangling_wire_36,N__10608}),
            .RCLKE(),
            .RCLK(N__22829),
            .RE(N__22907),
            .WCLKE(N__10634),
            .WCLK(N__22828),
            .WE(N__10635));
    IO_PAD led_obuft_3_iopad (
            .OE(N__23173),
            .DIN(N__23172),
            .DOUT(N__23171),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__23173),
            .PADOUT(N__23172),
            .PADIN(N__23171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__23164),
            .DIN(N__23163),
            .DOUT(N__23162),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__23164),
            .PADOUT(N__23163),
            .PADIN(N__23162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__23155),
            .DIN(N__23154),
            .DOUT(N__23153),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__23155),
            .PADOUT(N__23154),
            .PADIN(N__23153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__23146),
            .DIN(N__23145),
            .DOUT(N__23144),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__23146),
            .PADOUT(N__23145),
            .PADIN(N__23144),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__22807),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__23137),
            .DIN(N__23136),
            .DOUT(N__23135),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__23137),
            .PADOUT(N__23136),
            .PADIN(N__23135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__23128),
            .DIN(N__23127),
            .DOUT(N__23126),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__23128),
            .PADOUT(N__23127),
            .PADIN(N__23126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__23119),
            .DIN(N__23118),
            .DOUT(N__23117),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__23119),
            .PADOUT(N__23118),
            .PADIN(N__23117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__23110),
            .DIN(N__23109),
            .DOUT(N__23108),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__23110),
            .PADOUT(N__23109),
            .PADIN(N__23108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__23101),
            .DIN(N__23100),
            .DOUT(N__23099),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__23101),
            .PADOUT(N__23100),
            .PADIN(N__23099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10086),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__23092),
            .DIN(N__23091),
            .DOUT(N__23090),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__23092),
            .PADOUT(N__23091),
            .PADIN(N__23090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5648 (
            .O(N__23073),
            .I(N__23070));
    LocalMux I__5647 (
            .O(N__23070),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__5646 (
            .O(N__23067),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__5645 (
            .O(N__23064),
            .I(N__23060));
    InMux I__5644 (
            .O(N__23063),
            .I(N__23057));
    LocalMux I__5643 (
            .O(N__23060),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__5642 (
            .O(N__23057),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__5641 (
            .O(N__23052),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__5640 (
            .O(N__23049),
            .I(N__23044));
    InMux I__5639 (
            .O(N__23048),
            .I(N__23039));
    InMux I__5638 (
            .O(N__23047),
            .I(N__23039));
    LocalMux I__5637 (
            .O(N__23044),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__5636 (
            .O(N__23039),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__5635 (
            .O(N__23034),
            .I(N__23031));
    InMux I__5634 (
            .O(N__23031),
            .I(N__23028));
    LocalMux I__5633 (
            .O(N__23028),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__5632 (
            .O(N__23025),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__5631 (
            .O(N__23022),
            .I(N__23017));
    InMux I__5630 (
            .O(N__23021),
            .I(N__23013));
    InMux I__5629 (
            .O(N__23020),
            .I(N__23010));
    LocalMux I__5628 (
            .O(N__23017),
            .I(N__23007));
    InMux I__5627 (
            .O(N__23016),
            .I(N__23004));
    LocalMux I__5626 (
            .O(N__23013),
            .I(buart__rx_ser_clk));
    LocalMux I__5625 (
            .O(N__23010),
            .I(buart__rx_ser_clk));
    Odrv4 I__5624 (
            .O(N__23007),
            .I(buart__rx_ser_clk));
    LocalMux I__5623 (
            .O(N__23004),
            .I(buart__rx_ser_clk));
    CascadeMux I__5622 (
            .O(N__22995),
            .I(N__22991));
    CascadeMux I__5621 (
            .O(N__22994),
            .I(N__22984));
    InMux I__5620 (
            .O(N__22991),
            .I(N__22975));
    InMux I__5619 (
            .O(N__22990),
            .I(N__22975));
    InMux I__5618 (
            .O(N__22989),
            .I(N__22970));
    InMux I__5617 (
            .O(N__22988),
            .I(N__22970));
    InMux I__5616 (
            .O(N__22987),
            .I(N__22961));
    InMux I__5615 (
            .O(N__22984),
            .I(N__22961));
    InMux I__5614 (
            .O(N__22983),
            .I(N__22961));
    InMux I__5613 (
            .O(N__22982),
            .I(N__22961));
    InMux I__5612 (
            .O(N__22981),
            .I(N__22958));
    InMux I__5611 (
            .O(N__22980),
            .I(N__22955));
    LocalMux I__5610 (
            .O(N__22975),
            .I(N__22952));
    LocalMux I__5609 (
            .O(N__22970),
            .I(N__22949));
    LocalMux I__5608 (
            .O(N__22961),
            .I(N__22946));
    LocalMux I__5607 (
            .O(N__22958),
            .I(N__22943));
    LocalMux I__5606 (
            .O(N__22955),
            .I(buart__rx_startbit));
    Odrv4 I__5605 (
            .O(N__22952),
            .I(buart__rx_startbit));
    Odrv4 I__5604 (
            .O(N__22949),
            .I(buart__rx_startbit));
    Odrv4 I__5603 (
            .O(N__22946),
            .I(buart__rx_startbit));
    Odrv4 I__5602 (
            .O(N__22943),
            .I(buart__rx_startbit));
    InMux I__5601 (
            .O(N__22932),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__5600 (
            .O(N__22929),
            .I(N__22925));
    InMux I__5599 (
            .O(N__22928),
            .I(N__22922));
    InMux I__5598 (
            .O(N__22925),
            .I(N__22919));
    LocalMux I__5597 (
            .O(N__22922),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__5596 (
            .O(N__22919),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    IoInMux I__5595 (
            .O(N__22914),
            .I(N__22911));
    LocalMux I__5594 (
            .O(N__22911),
            .I(N__22908));
    IoSpan4Mux I__5593 (
            .O(N__22908),
            .I(N__22904));
    SRMux I__5592 (
            .O(N__22907),
            .I(N__22901));
    IoSpan4Mux I__5591 (
            .O(N__22904),
            .I(N__22896));
    LocalMux I__5590 (
            .O(N__22901),
            .I(N__22893));
    InMux I__5589 (
            .O(N__22900),
            .I(N__22890));
    InMux I__5588 (
            .O(N__22899),
            .I(N__22887));
    Span4Mux_s2_h I__5587 (
            .O(N__22896),
            .I(N__22882));
    Span4Mux_v I__5586 (
            .O(N__22893),
            .I(N__22882));
    LocalMux I__5585 (
            .O(N__22890),
            .I(N__22877));
    LocalMux I__5584 (
            .O(N__22887),
            .I(N__22877));
    Span4Mux_h I__5583 (
            .O(N__22882),
            .I(N__22872));
    Span4Mux_s1_h I__5582 (
            .O(N__22877),
            .I(N__22872));
    Odrv4 I__5581 (
            .O(N__22872),
            .I(CONSTANT_ONE_NET));
    InMux I__5580 (
            .O(N__22869),
            .I(N__22866));
    LocalMux I__5579 (
            .O(N__22866),
            .I(N__22863));
    Odrv4 I__5578 (
            .O(N__22863),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    InMux I__5577 (
            .O(N__22860),
            .I(N__22857));
    LocalMux I__5576 (
            .O(N__22857),
            .I(N__22771));
    ClkMux I__5575 (
            .O(N__22856),
            .I(N__22602));
    ClkMux I__5574 (
            .O(N__22855),
            .I(N__22602));
    ClkMux I__5573 (
            .O(N__22854),
            .I(N__22602));
    ClkMux I__5572 (
            .O(N__22853),
            .I(N__22602));
    ClkMux I__5571 (
            .O(N__22852),
            .I(N__22602));
    ClkMux I__5570 (
            .O(N__22851),
            .I(N__22602));
    ClkMux I__5569 (
            .O(N__22850),
            .I(N__22602));
    ClkMux I__5568 (
            .O(N__22849),
            .I(N__22602));
    ClkMux I__5567 (
            .O(N__22848),
            .I(N__22602));
    ClkMux I__5566 (
            .O(N__22847),
            .I(N__22602));
    ClkMux I__5565 (
            .O(N__22846),
            .I(N__22602));
    ClkMux I__5564 (
            .O(N__22845),
            .I(N__22602));
    ClkMux I__5563 (
            .O(N__22844),
            .I(N__22602));
    ClkMux I__5562 (
            .O(N__22843),
            .I(N__22602));
    ClkMux I__5561 (
            .O(N__22842),
            .I(N__22602));
    ClkMux I__5560 (
            .O(N__22841),
            .I(N__22602));
    ClkMux I__5559 (
            .O(N__22840),
            .I(N__22602));
    ClkMux I__5558 (
            .O(N__22839),
            .I(N__22602));
    ClkMux I__5557 (
            .O(N__22838),
            .I(N__22602));
    ClkMux I__5556 (
            .O(N__22837),
            .I(N__22602));
    ClkMux I__5555 (
            .O(N__22836),
            .I(N__22602));
    ClkMux I__5554 (
            .O(N__22835),
            .I(N__22602));
    ClkMux I__5553 (
            .O(N__22834),
            .I(N__22602));
    ClkMux I__5552 (
            .O(N__22833),
            .I(N__22602));
    ClkMux I__5551 (
            .O(N__22832),
            .I(N__22602));
    ClkMux I__5550 (
            .O(N__22831),
            .I(N__22602));
    ClkMux I__5549 (
            .O(N__22830),
            .I(N__22602));
    ClkMux I__5548 (
            .O(N__22829),
            .I(N__22602));
    ClkMux I__5547 (
            .O(N__22828),
            .I(N__22602));
    ClkMux I__5546 (
            .O(N__22827),
            .I(N__22602));
    ClkMux I__5545 (
            .O(N__22826),
            .I(N__22602));
    ClkMux I__5544 (
            .O(N__22825),
            .I(N__22602));
    ClkMux I__5543 (
            .O(N__22824),
            .I(N__22602));
    ClkMux I__5542 (
            .O(N__22823),
            .I(N__22602));
    ClkMux I__5541 (
            .O(N__22822),
            .I(N__22602));
    ClkMux I__5540 (
            .O(N__22821),
            .I(N__22602));
    ClkMux I__5539 (
            .O(N__22820),
            .I(N__22602));
    ClkMux I__5538 (
            .O(N__22819),
            .I(N__22602));
    ClkMux I__5537 (
            .O(N__22818),
            .I(N__22602));
    ClkMux I__5536 (
            .O(N__22817),
            .I(N__22602));
    ClkMux I__5535 (
            .O(N__22816),
            .I(N__22602));
    ClkMux I__5534 (
            .O(N__22815),
            .I(N__22602));
    ClkMux I__5533 (
            .O(N__22814),
            .I(N__22602));
    ClkMux I__5532 (
            .O(N__22813),
            .I(N__22602));
    ClkMux I__5531 (
            .O(N__22812),
            .I(N__22602));
    ClkMux I__5530 (
            .O(N__22811),
            .I(N__22602));
    ClkMux I__5529 (
            .O(N__22810),
            .I(N__22602));
    ClkMux I__5528 (
            .O(N__22809),
            .I(N__22602));
    ClkMux I__5527 (
            .O(N__22808),
            .I(N__22602));
    ClkMux I__5526 (
            .O(N__22807),
            .I(N__22602));
    ClkMux I__5525 (
            .O(N__22806),
            .I(N__22602));
    ClkMux I__5524 (
            .O(N__22805),
            .I(N__22602));
    ClkMux I__5523 (
            .O(N__22804),
            .I(N__22602));
    ClkMux I__5522 (
            .O(N__22803),
            .I(N__22602));
    ClkMux I__5521 (
            .O(N__22802),
            .I(N__22602));
    ClkMux I__5520 (
            .O(N__22801),
            .I(N__22602));
    ClkMux I__5519 (
            .O(N__22800),
            .I(N__22602));
    ClkMux I__5518 (
            .O(N__22799),
            .I(N__22602));
    ClkMux I__5517 (
            .O(N__22798),
            .I(N__22602));
    ClkMux I__5516 (
            .O(N__22797),
            .I(N__22602));
    ClkMux I__5515 (
            .O(N__22796),
            .I(N__22602));
    ClkMux I__5514 (
            .O(N__22795),
            .I(N__22602));
    ClkMux I__5513 (
            .O(N__22794),
            .I(N__22602));
    ClkMux I__5512 (
            .O(N__22793),
            .I(N__22602));
    ClkMux I__5511 (
            .O(N__22792),
            .I(N__22602));
    ClkMux I__5510 (
            .O(N__22791),
            .I(N__22602));
    ClkMux I__5509 (
            .O(N__22790),
            .I(N__22602));
    ClkMux I__5508 (
            .O(N__22789),
            .I(N__22602));
    ClkMux I__5507 (
            .O(N__22788),
            .I(N__22602));
    ClkMux I__5506 (
            .O(N__22787),
            .I(N__22602));
    ClkMux I__5505 (
            .O(N__22786),
            .I(N__22602));
    ClkMux I__5504 (
            .O(N__22785),
            .I(N__22602));
    ClkMux I__5503 (
            .O(N__22784),
            .I(N__22602));
    ClkMux I__5502 (
            .O(N__22783),
            .I(N__22602));
    ClkMux I__5501 (
            .O(N__22782),
            .I(N__22602));
    ClkMux I__5500 (
            .O(N__22781),
            .I(N__22602));
    ClkMux I__5499 (
            .O(N__22780),
            .I(N__22602));
    ClkMux I__5498 (
            .O(N__22779),
            .I(N__22602));
    ClkMux I__5497 (
            .O(N__22778),
            .I(N__22602));
    ClkMux I__5496 (
            .O(N__22777),
            .I(N__22602));
    ClkMux I__5495 (
            .O(N__22776),
            .I(N__22602));
    ClkMux I__5494 (
            .O(N__22775),
            .I(N__22602));
    ClkMux I__5493 (
            .O(N__22774),
            .I(N__22602));
    Glb2LocalMux I__5492 (
            .O(N__22771),
            .I(N__22602));
    GlobalMux I__5491 (
            .O(N__22602),
            .I(N__22599));
    gio2CtrlBuf I__5490 (
            .O(N__22599),
            .I(clk_g));
    CascadeMux I__5489 (
            .O(N__22596),
            .I(N__22593));
    InMux I__5488 (
            .O(N__22593),
            .I(N__22590));
    LocalMux I__5487 (
            .O(N__22590),
            .I(N__22587));
    Span4Mux_v I__5486 (
            .O(N__22587),
            .I(N__22584));
    Span4Mux_h I__5485 (
            .O(N__22584),
            .I(N__22577));
    InMux I__5484 (
            .O(N__22583),
            .I(N__22574));
    InMux I__5483 (
            .O(N__22582),
            .I(N__22567));
    InMux I__5482 (
            .O(N__22581),
            .I(N__22567));
    InMux I__5481 (
            .O(N__22580),
            .I(N__22567));
    Odrv4 I__5480 (
            .O(N__22577),
            .I(bu_rx_data_rdy));
    LocalMux I__5479 (
            .O(N__22574),
            .I(bu_rx_data_rdy));
    LocalMux I__5478 (
            .O(N__22567),
            .I(bu_rx_data_rdy));
    InMux I__5477 (
            .O(N__22560),
            .I(N__22551));
    InMux I__5476 (
            .O(N__22559),
            .I(N__22548));
    InMux I__5475 (
            .O(N__22558),
            .I(N__22545));
    InMux I__5474 (
            .O(N__22557),
            .I(N__22542));
    InMux I__5473 (
            .O(N__22556),
            .I(N__22539));
    SRMux I__5472 (
            .O(N__22555),
            .I(N__22534));
    InMux I__5471 (
            .O(N__22554),
            .I(N__22534));
    LocalMux I__5470 (
            .O(N__22551),
            .I(N__22492));
    LocalMux I__5469 (
            .O(N__22548),
            .I(N__22489));
    LocalMux I__5468 (
            .O(N__22545),
            .I(N__22486));
    LocalMux I__5467 (
            .O(N__22542),
            .I(N__22469));
    LocalMux I__5466 (
            .O(N__22539),
            .I(N__22466));
    LocalMux I__5465 (
            .O(N__22534),
            .I(N__22463));
    SRMux I__5464 (
            .O(N__22533),
            .I(N__22344));
    SRMux I__5463 (
            .O(N__22532),
            .I(N__22344));
    SRMux I__5462 (
            .O(N__22531),
            .I(N__22344));
    SRMux I__5461 (
            .O(N__22530),
            .I(N__22344));
    SRMux I__5460 (
            .O(N__22529),
            .I(N__22344));
    SRMux I__5459 (
            .O(N__22528),
            .I(N__22344));
    SRMux I__5458 (
            .O(N__22527),
            .I(N__22344));
    SRMux I__5457 (
            .O(N__22526),
            .I(N__22344));
    SRMux I__5456 (
            .O(N__22525),
            .I(N__22344));
    SRMux I__5455 (
            .O(N__22524),
            .I(N__22344));
    SRMux I__5454 (
            .O(N__22523),
            .I(N__22344));
    SRMux I__5453 (
            .O(N__22522),
            .I(N__22344));
    SRMux I__5452 (
            .O(N__22521),
            .I(N__22344));
    SRMux I__5451 (
            .O(N__22520),
            .I(N__22344));
    SRMux I__5450 (
            .O(N__22519),
            .I(N__22344));
    SRMux I__5449 (
            .O(N__22518),
            .I(N__22344));
    SRMux I__5448 (
            .O(N__22517),
            .I(N__22344));
    SRMux I__5447 (
            .O(N__22516),
            .I(N__22344));
    SRMux I__5446 (
            .O(N__22515),
            .I(N__22344));
    SRMux I__5445 (
            .O(N__22514),
            .I(N__22344));
    SRMux I__5444 (
            .O(N__22513),
            .I(N__22344));
    SRMux I__5443 (
            .O(N__22512),
            .I(N__22344));
    SRMux I__5442 (
            .O(N__22511),
            .I(N__22344));
    SRMux I__5441 (
            .O(N__22510),
            .I(N__22344));
    SRMux I__5440 (
            .O(N__22509),
            .I(N__22344));
    SRMux I__5439 (
            .O(N__22508),
            .I(N__22344));
    SRMux I__5438 (
            .O(N__22507),
            .I(N__22344));
    SRMux I__5437 (
            .O(N__22506),
            .I(N__22344));
    SRMux I__5436 (
            .O(N__22505),
            .I(N__22344));
    SRMux I__5435 (
            .O(N__22504),
            .I(N__22344));
    SRMux I__5434 (
            .O(N__22503),
            .I(N__22344));
    SRMux I__5433 (
            .O(N__22502),
            .I(N__22344));
    SRMux I__5432 (
            .O(N__22501),
            .I(N__22344));
    SRMux I__5431 (
            .O(N__22500),
            .I(N__22344));
    SRMux I__5430 (
            .O(N__22499),
            .I(N__22344));
    SRMux I__5429 (
            .O(N__22498),
            .I(N__22344));
    SRMux I__5428 (
            .O(N__22497),
            .I(N__22344));
    SRMux I__5427 (
            .O(N__22496),
            .I(N__22344));
    SRMux I__5426 (
            .O(N__22495),
            .I(N__22344));
    Glb2LocalMux I__5425 (
            .O(N__22492),
            .I(N__22344));
    Glb2LocalMux I__5424 (
            .O(N__22489),
            .I(N__22344));
    Glb2LocalMux I__5423 (
            .O(N__22486),
            .I(N__22344));
    SRMux I__5422 (
            .O(N__22485),
            .I(N__22344));
    SRMux I__5421 (
            .O(N__22484),
            .I(N__22344));
    SRMux I__5420 (
            .O(N__22483),
            .I(N__22344));
    SRMux I__5419 (
            .O(N__22482),
            .I(N__22344));
    SRMux I__5418 (
            .O(N__22481),
            .I(N__22344));
    SRMux I__5417 (
            .O(N__22480),
            .I(N__22344));
    SRMux I__5416 (
            .O(N__22479),
            .I(N__22344));
    SRMux I__5415 (
            .O(N__22478),
            .I(N__22344));
    SRMux I__5414 (
            .O(N__22477),
            .I(N__22344));
    SRMux I__5413 (
            .O(N__22476),
            .I(N__22344));
    SRMux I__5412 (
            .O(N__22475),
            .I(N__22344));
    SRMux I__5411 (
            .O(N__22474),
            .I(N__22344));
    SRMux I__5410 (
            .O(N__22473),
            .I(N__22344));
    SRMux I__5409 (
            .O(N__22472),
            .I(N__22344));
    Glb2LocalMux I__5408 (
            .O(N__22469),
            .I(N__22344));
    Glb2LocalMux I__5407 (
            .O(N__22466),
            .I(N__22344));
    Glb2LocalMux I__5406 (
            .O(N__22463),
            .I(N__22344));
    GlobalMux I__5405 (
            .O(N__22344),
            .I(N__22341));
    gio2CtrlBuf I__5404 (
            .O(N__22341),
            .I(rst_g));
    IoInMux I__5403 (
            .O(N__22338),
            .I(N__22335));
    LocalMux I__5402 (
            .O(N__22335),
            .I(bu_rx_data_rdy_0));
    InMux I__5401 (
            .O(N__22332),
            .I(N__22329));
    LocalMux I__5400 (
            .O(N__22329),
            .I(\resetGen.r_m3_i_a3_0_2 ));
    InMux I__5399 (
            .O(N__22326),
            .I(N__22323));
    LocalMux I__5398 (
            .O(N__22323),
            .I(N_6));
    CascadeMux I__5397 (
            .O(N__22320),
            .I(N__22317));
    InMux I__5396 (
            .O(N__22317),
            .I(N__22314));
    LocalMux I__5395 (
            .O(N__22314),
            .I(N__22311));
    Span4Mux_v I__5394 (
            .O(N__22311),
            .I(N__22308));
    Odrv4 I__5393 (
            .O(N__22308),
            .I(Lab_UT_dictrl_next_state_0_1_2));
    InMux I__5392 (
            .O(N__22305),
            .I(N__22302));
    LocalMux I__5391 (
            .O(N__22302),
            .I(Lab_UT_dictrl_next_state_0_0_0));
    CEMux I__5390 (
            .O(N__22299),
            .I(N__22296));
    LocalMux I__5389 (
            .O(N__22296),
            .I(N__22292));
    CEMux I__5388 (
            .O(N__22295),
            .I(N__22289));
    Span4Mux_s0_h I__5387 (
            .O(N__22292),
            .I(N__22286));
    LocalMux I__5386 (
            .O(N__22289),
            .I(N__22283));
    Span4Mux_v I__5385 (
            .O(N__22286),
            .I(N__22277));
    Span4Mux_h I__5384 (
            .O(N__22283),
            .I(N__22277));
    CEMux I__5383 (
            .O(N__22282),
            .I(N__22274));
    Odrv4 I__5382 (
            .O(N__22277),
            .I(rst_RNIAL6V33));
    LocalMux I__5381 (
            .O(N__22274),
            .I(rst_RNIAL6V33));
    CascadeMux I__5380 (
            .O(N__22269),
            .I(N__22265));
    CascadeMux I__5379 (
            .O(N__22268),
            .I(N__22259));
    InMux I__5378 (
            .O(N__22265),
            .I(N__22256));
    CascadeMux I__5377 (
            .O(N__22264),
            .I(N__22253));
    CascadeMux I__5376 (
            .O(N__22263),
            .I(N__22244));
    InMux I__5375 (
            .O(N__22262),
            .I(N__22237));
    InMux I__5374 (
            .O(N__22259),
            .I(N__22237));
    LocalMux I__5373 (
            .O(N__22256),
            .I(N__22234));
    InMux I__5372 (
            .O(N__22253),
            .I(N__22227));
    InMux I__5371 (
            .O(N__22252),
            .I(N__22227));
    InMux I__5370 (
            .O(N__22251),
            .I(N__22227));
    InMux I__5369 (
            .O(N__22250),
            .I(N__22224));
    CascadeMux I__5368 (
            .O(N__22249),
            .I(N__22221));
    InMux I__5367 (
            .O(N__22248),
            .I(N__22209));
    InMux I__5366 (
            .O(N__22247),
            .I(N__22209));
    InMux I__5365 (
            .O(N__22244),
            .I(N__22209));
    InMux I__5364 (
            .O(N__22243),
            .I(N__22206));
    InMux I__5363 (
            .O(N__22242),
            .I(N__22203));
    LocalMux I__5362 (
            .O(N__22237),
            .I(N__22193));
    Span4Mux_v I__5361 (
            .O(N__22234),
            .I(N__22193));
    LocalMux I__5360 (
            .O(N__22227),
            .I(N__22188));
    LocalMux I__5359 (
            .O(N__22224),
            .I(N__22188));
    InMux I__5358 (
            .O(N__22221),
            .I(N__22185));
    InMux I__5357 (
            .O(N__22220),
            .I(N__22182));
    InMux I__5356 (
            .O(N__22219),
            .I(N__22173));
    InMux I__5355 (
            .O(N__22218),
            .I(N__22173));
    InMux I__5354 (
            .O(N__22217),
            .I(N__22173));
    InMux I__5353 (
            .O(N__22216),
            .I(N__22173));
    LocalMux I__5352 (
            .O(N__22209),
            .I(N__22168));
    LocalMux I__5351 (
            .O(N__22206),
            .I(N__22168));
    LocalMux I__5350 (
            .O(N__22203),
            .I(N__22165));
    InMux I__5349 (
            .O(N__22202),
            .I(N__22162));
    InMux I__5348 (
            .O(N__22201),
            .I(N__22159));
    InMux I__5347 (
            .O(N__22200),
            .I(N__22154));
    InMux I__5346 (
            .O(N__22199),
            .I(N__22154));
    InMux I__5345 (
            .O(N__22198),
            .I(N__22151));
    Span4Mux_v I__5344 (
            .O(N__22193),
            .I(N__22146));
    Span4Mux_v I__5343 (
            .O(N__22188),
            .I(N__22146));
    LocalMux I__5342 (
            .O(N__22185),
            .I(N__22137));
    LocalMux I__5341 (
            .O(N__22182),
            .I(N__22137));
    LocalMux I__5340 (
            .O(N__22173),
            .I(N__22137));
    Span4Mux_v I__5339 (
            .O(N__22168),
            .I(N__22137));
    Span4Mux_h I__5338 (
            .O(N__22165),
            .I(N__22134));
    LocalMux I__5337 (
            .O(N__22162),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    LocalMux I__5336 (
            .O(N__22159),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    LocalMux I__5335 (
            .O(N__22154),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    LocalMux I__5334 (
            .O(N__22151),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5333 (
            .O(N__22146),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5332 (
            .O(N__22137),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    Odrv4 I__5331 (
            .O(N__22134),
            .I(\Lab_UT.dictrl.stateZ0Z_0 ));
    CascadeMux I__5330 (
            .O(N__22119),
            .I(N__22116));
    InMux I__5329 (
            .O(N__22116),
            .I(N__22113));
    LocalMux I__5328 (
            .O(N__22113),
            .I(N__22110));
    Odrv12 I__5327 (
            .O(N__22110),
            .I(\Lab_UT.dictrl.m46_i_0_a5_1 ));
    InMux I__5326 (
            .O(N__22107),
            .I(N__22098));
    InMux I__5325 (
            .O(N__22106),
            .I(N__22098));
    InMux I__5324 (
            .O(N__22105),
            .I(N__22085));
    InMux I__5323 (
            .O(N__22104),
            .I(N__22082));
    InMux I__5322 (
            .O(N__22103),
            .I(N__22079));
    LocalMux I__5321 (
            .O(N__22098),
            .I(N__22076));
    InMux I__5320 (
            .O(N__22097),
            .I(N__22073));
    InMux I__5319 (
            .O(N__22096),
            .I(N__22068));
    InMux I__5318 (
            .O(N__22095),
            .I(N__22068));
    InMux I__5317 (
            .O(N__22094),
            .I(N__22065));
    InMux I__5316 (
            .O(N__22093),
            .I(N__22062));
    InMux I__5315 (
            .O(N__22092),
            .I(N__22057));
    InMux I__5314 (
            .O(N__22091),
            .I(N__22057));
    InMux I__5313 (
            .O(N__22090),
            .I(N__22049));
    InMux I__5312 (
            .O(N__22089),
            .I(N__22049));
    InMux I__5311 (
            .O(N__22088),
            .I(N__22049));
    LocalMux I__5310 (
            .O(N__22085),
            .I(N__22044));
    LocalMux I__5309 (
            .O(N__22082),
            .I(N__22044));
    LocalMux I__5308 (
            .O(N__22079),
            .I(N__22041));
    Span4Mux_v I__5307 (
            .O(N__22076),
            .I(N__22033));
    LocalMux I__5306 (
            .O(N__22073),
            .I(N__22033));
    LocalMux I__5305 (
            .O(N__22068),
            .I(N__22024));
    LocalMux I__5304 (
            .O(N__22065),
            .I(N__22024));
    LocalMux I__5303 (
            .O(N__22062),
            .I(N__22024));
    LocalMux I__5302 (
            .O(N__22057),
            .I(N__22024));
    InMux I__5301 (
            .O(N__22056),
            .I(N__22021));
    LocalMux I__5300 (
            .O(N__22049),
            .I(N__22017));
    Span4Mux_v I__5299 (
            .O(N__22044),
            .I(N__22012));
    Span4Mux_s3_h I__5298 (
            .O(N__22041),
            .I(N__22012));
    InMux I__5297 (
            .O(N__22040),
            .I(N__22009));
    InMux I__5296 (
            .O(N__22039),
            .I(N__22004));
    InMux I__5295 (
            .O(N__22038),
            .I(N__22004));
    Span4Mux_h I__5294 (
            .O(N__22033),
            .I(N__21997));
    Span4Mux_v I__5293 (
            .O(N__22024),
            .I(N__21997));
    LocalMux I__5292 (
            .O(N__22021),
            .I(N__21997));
    InMux I__5291 (
            .O(N__22020),
            .I(N__21994));
    Odrv4 I__5290 (
            .O(N__22017),
            .I(\Lab_UT.dictrl.N_86 ));
    Odrv4 I__5289 (
            .O(N__22012),
            .I(\Lab_UT.dictrl.N_86 ));
    LocalMux I__5288 (
            .O(N__22009),
            .I(\Lab_UT.dictrl.N_86 ));
    LocalMux I__5287 (
            .O(N__22004),
            .I(\Lab_UT.dictrl.N_86 ));
    Odrv4 I__5286 (
            .O(N__21997),
            .I(\Lab_UT.dictrl.N_86 ));
    LocalMux I__5285 (
            .O(N__21994),
            .I(\Lab_UT.dictrl.N_86 ));
    InMux I__5284 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__5283 (
            .O(N__21978),
            .I(\Lab_UT.dictrl.N_8 ));
    CascadeMux I__5282 (
            .O(N__21975),
            .I(N__21972));
    InMux I__5281 (
            .O(N__21972),
            .I(N__21969));
    LocalMux I__5280 (
            .O(N__21969),
            .I(N__21965));
    InMux I__5279 (
            .O(N__21968),
            .I(N__21962));
    Span4Mux_h I__5278 (
            .O(N__21965),
            .I(N__21959));
    LocalMux I__5277 (
            .O(N__21962),
            .I(N__21956));
    Odrv4 I__5276 (
            .O(N__21959),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    Odrv12 I__5275 (
            .O(N__21956),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    CascadeMux I__5274 (
            .O(N__21951),
            .I(N__21938));
    CascadeMux I__5273 (
            .O(N__21950),
            .I(N__21932));
    InMux I__5272 (
            .O(N__21949),
            .I(N__21926));
    CascadeMux I__5271 (
            .O(N__21948),
            .I(N__21923));
    InMux I__5270 (
            .O(N__21947),
            .I(N__21920));
    CascadeMux I__5269 (
            .O(N__21946),
            .I(N__21917));
    InMux I__5268 (
            .O(N__21945),
            .I(N__21914));
    CascadeMux I__5267 (
            .O(N__21944),
            .I(N__21907));
    CascadeMux I__5266 (
            .O(N__21943),
            .I(N__21904));
    CascadeMux I__5265 (
            .O(N__21942),
            .I(N__21900));
    InMux I__5264 (
            .O(N__21941),
            .I(N__21890));
    InMux I__5263 (
            .O(N__21938),
            .I(N__21890));
    InMux I__5262 (
            .O(N__21937),
            .I(N__21890));
    CascadeMux I__5261 (
            .O(N__21936),
            .I(N__21887));
    CascadeMux I__5260 (
            .O(N__21935),
            .I(N__21882));
    InMux I__5259 (
            .O(N__21932),
            .I(N__21876));
    InMux I__5258 (
            .O(N__21931),
            .I(N__21873));
    InMux I__5257 (
            .O(N__21930),
            .I(N__21868));
    InMux I__5256 (
            .O(N__21929),
            .I(N__21868));
    LocalMux I__5255 (
            .O(N__21926),
            .I(N__21865));
    InMux I__5254 (
            .O(N__21923),
            .I(N__21862));
    LocalMux I__5253 (
            .O(N__21920),
            .I(N__21859));
    InMux I__5252 (
            .O(N__21917),
            .I(N__21856));
    LocalMux I__5251 (
            .O(N__21914),
            .I(N__21853));
    InMux I__5250 (
            .O(N__21913),
            .I(N__21840));
    InMux I__5249 (
            .O(N__21912),
            .I(N__21840));
    InMux I__5248 (
            .O(N__21911),
            .I(N__21840));
    InMux I__5247 (
            .O(N__21910),
            .I(N__21840));
    InMux I__5246 (
            .O(N__21907),
            .I(N__21840));
    InMux I__5245 (
            .O(N__21904),
            .I(N__21840));
    CascadeMux I__5244 (
            .O(N__21903),
            .I(N__21832));
    InMux I__5243 (
            .O(N__21900),
            .I(N__21827));
    InMux I__5242 (
            .O(N__21899),
            .I(N__21827));
    InMux I__5241 (
            .O(N__21898),
            .I(N__21824));
    InMux I__5240 (
            .O(N__21897),
            .I(N__21821));
    LocalMux I__5239 (
            .O(N__21890),
            .I(N__21817));
    InMux I__5238 (
            .O(N__21887),
            .I(N__21802));
    InMux I__5237 (
            .O(N__21886),
            .I(N__21802));
    InMux I__5236 (
            .O(N__21885),
            .I(N__21802));
    InMux I__5235 (
            .O(N__21882),
            .I(N__21802));
    InMux I__5234 (
            .O(N__21881),
            .I(N__21802));
    InMux I__5233 (
            .O(N__21880),
            .I(N__21802));
    InMux I__5232 (
            .O(N__21879),
            .I(N__21802));
    LocalMux I__5231 (
            .O(N__21876),
            .I(N__21787));
    LocalMux I__5230 (
            .O(N__21873),
            .I(N__21787));
    LocalMux I__5229 (
            .O(N__21868),
            .I(N__21787));
    Span4Mux_h I__5228 (
            .O(N__21865),
            .I(N__21787));
    LocalMux I__5227 (
            .O(N__21862),
            .I(N__21787));
    Span4Mux_v I__5226 (
            .O(N__21859),
            .I(N__21787));
    LocalMux I__5225 (
            .O(N__21856),
            .I(N__21787));
    Span12Mux_s9_v I__5224 (
            .O(N__21853),
            .I(N__21782));
    LocalMux I__5223 (
            .O(N__21840),
            .I(N__21782));
    InMux I__5222 (
            .O(N__21839),
            .I(N__21779));
    InMux I__5221 (
            .O(N__21838),
            .I(N__21774));
    InMux I__5220 (
            .O(N__21837),
            .I(N__21774));
    InMux I__5219 (
            .O(N__21836),
            .I(N__21767));
    InMux I__5218 (
            .O(N__21835),
            .I(N__21767));
    InMux I__5217 (
            .O(N__21832),
            .I(N__21767));
    LocalMux I__5216 (
            .O(N__21827),
            .I(N__21760));
    LocalMux I__5215 (
            .O(N__21824),
            .I(N__21760));
    LocalMux I__5214 (
            .O(N__21821),
            .I(N__21760));
    InMux I__5213 (
            .O(N__21820),
            .I(N__21757));
    Span4Mux_v I__5212 (
            .O(N__21817),
            .I(N__21750));
    LocalMux I__5211 (
            .O(N__21802),
            .I(N__21750));
    Span4Mux_v I__5210 (
            .O(N__21787),
            .I(N__21750));
    Odrv12 I__5209 (
            .O(N__21782),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    LocalMux I__5208 (
            .O(N__21779),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    LocalMux I__5207 (
            .O(N__21774),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    LocalMux I__5206 (
            .O(N__21767),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    Odrv12 I__5205 (
            .O(N__21760),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    LocalMux I__5204 (
            .O(N__21757),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    Odrv4 I__5203 (
            .O(N__21750),
            .I(Lab_UT_dictrl_un1_next_state66_0));
    InMux I__5202 (
            .O(N__21735),
            .I(N__21732));
    LocalMux I__5201 (
            .O(N__21732),
            .I(\Lab_UT.dictrl.m46_i_0_0_0 ));
    InMux I__5200 (
            .O(N__21729),
            .I(N__21725));
    InMux I__5199 (
            .O(N__21728),
            .I(N__21717));
    LocalMux I__5198 (
            .O(N__21725),
            .I(N__21714));
    InMux I__5197 (
            .O(N__21724),
            .I(N__21709));
    InMux I__5196 (
            .O(N__21723),
            .I(N__21709));
    InMux I__5195 (
            .O(N__21722),
            .I(N__21706));
    InMux I__5194 (
            .O(N__21721),
            .I(N__21703));
    InMux I__5193 (
            .O(N__21720),
            .I(N__21700));
    LocalMux I__5192 (
            .O(N__21717),
            .I(N__21695));
    Span4Mux_v I__5191 (
            .O(N__21714),
            .I(N__21692));
    LocalMux I__5190 (
            .O(N__21709),
            .I(N__21687));
    LocalMux I__5189 (
            .O(N__21706),
            .I(N__21687));
    LocalMux I__5188 (
            .O(N__21703),
            .I(N__21682));
    LocalMux I__5187 (
            .O(N__21700),
            .I(N__21682));
    InMux I__5186 (
            .O(N__21699),
            .I(N__21679));
    InMux I__5185 (
            .O(N__21698),
            .I(N__21676));
    Span4Mux_h I__5184 (
            .O(N__21695),
            .I(N__21673));
    Span4Mux_h I__5183 (
            .O(N__21692),
            .I(N__21664));
    Span4Mux_v I__5182 (
            .O(N__21687),
            .I(N__21664));
    Span4Mux_v I__5181 (
            .O(N__21682),
            .I(N__21664));
    LocalMux I__5180 (
            .O(N__21679),
            .I(N__21664));
    LocalMux I__5179 (
            .O(N__21676),
            .I(bu_rx_data_i_3_1));
    Odrv4 I__5178 (
            .O(N__21673),
            .I(bu_rx_data_i_3_1));
    Odrv4 I__5177 (
            .O(N__21664),
            .I(bu_rx_data_i_3_1));
    InMux I__5176 (
            .O(N__21657),
            .I(N__21653));
    InMux I__5175 (
            .O(N__21656),
            .I(N__21645));
    LocalMux I__5174 (
            .O(N__21653),
            .I(N__21642));
    InMux I__5173 (
            .O(N__21652),
            .I(N__21639));
    InMux I__5172 (
            .O(N__21651),
            .I(N__21632));
    InMux I__5171 (
            .O(N__21650),
            .I(N__21632));
    InMux I__5170 (
            .O(N__21649),
            .I(N__21632));
    CascadeMux I__5169 (
            .O(N__21648),
            .I(N__21625));
    LocalMux I__5168 (
            .O(N__21645),
            .I(N__21622));
    Span4Mux_v I__5167 (
            .O(N__21642),
            .I(N__21614));
    LocalMux I__5166 (
            .O(N__21639),
            .I(N__21614));
    LocalMux I__5165 (
            .O(N__21632),
            .I(N__21614));
    InMux I__5164 (
            .O(N__21631),
            .I(N__21607));
    InMux I__5163 (
            .O(N__21630),
            .I(N__21607));
    InMux I__5162 (
            .O(N__21629),
            .I(N__21607));
    InMux I__5161 (
            .O(N__21628),
            .I(N__21602));
    InMux I__5160 (
            .O(N__21625),
            .I(N__21602));
    Span4Mux_h I__5159 (
            .O(N__21622),
            .I(N__21599));
    InMux I__5158 (
            .O(N__21621),
            .I(N__21596));
    Span4Mux_h I__5157 (
            .O(N__21614),
            .I(N__21589));
    LocalMux I__5156 (
            .O(N__21607),
            .I(N__21589));
    LocalMux I__5155 (
            .O(N__21602),
            .I(N__21589));
    Odrv4 I__5154 (
            .O(N__21599),
            .I(bu_rx_data_i_4_7));
    LocalMux I__5153 (
            .O(N__21596),
            .I(bu_rx_data_i_4_7));
    Odrv4 I__5152 (
            .O(N__21589),
            .I(bu_rx_data_i_4_7));
    CascadeMux I__5151 (
            .O(N__21582),
            .I(N__21576));
    CascadeMux I__5150 (
            .O(N__21581),
            .I(N__21573));
    CascadeMux I__5149 (
            .O(N__21580),
            .I(N__21568));
    CascadeMux I__5148 (
            .O(N__21579),
            .I(N__21565));
    InMux I__5147 (
            .O(N__21576),
            .I(N__21562));
    InMux I__5146 (
            .O(N__21573),
            .I(N__21557));
    CascadeMux I__5145 (
            .O(N__21572),
            .I(N__21553));
    InMux I__5144 (
            .O(N__21571),
            .I(N__21550));
    InMux I__5143 (
            .O(N__21568),
            .I(N__21547));
    InMux I__5142 (
            .O(N__21565),
            .I(N__21541));
    LocalMux I__5141 (
            .O(N__21562),
            .I(N__21536));
    InMux I__5140 (
            .O(N__21561),
            .I(N__21533));
    CascadeMux I__5139 (
            .O(N__21560),
            .I(N__21527));
    LocalMux I__5138 (
            .O(N__21557),
            .I(N__21524));
    InMux I__5137 (
            .O(N__21556),
            .I(N__21519));
    InMux I__5136 (
            .O(N__21553),
            .I(N__21519));
    LocalMux I__5135 (
            .O(N__21550),
            .I(N__21516));
    LocalMux I__5134 (
            .O(N__21547),
            .I(N__21513));
    InMux I__5133 (
            .O(N__21546),
            .I(N__21506));
    InMux I__5132 (
            .O(N__21545),
            .I(N__21506));
    InMux I__5131 (
            .O(N__21544),
            .I(N__21506));
    LocalMux I__5130 (
            .O(N__21541),
            .I(N__21503));
    CascadeMux I__5129 (
            .O(N__21540),
            .I(N__21499));
    CascadeMux I__5128 (
            .O(N__21539),
            .I(N__21496));
    Span4Mux_s2_h I__5127 (
            .O(N__21536),
            .I(N__21491));
    LocalMux I__5126 (
            .O(N__21533),
            .I(N__21491));
    InMux I__5125 (
            .O(N__21532),
            .I(N__21486));
    InMux I__5124 (
            .O(N__21531),
            .I(N__21486));
    InMux I__5123 (
            .O(N__21530),
            .I(N__21483));
    InMux I__5122 (
            .O(N__21527),
            .I(N__21480));
    Span4Mux_s2_h I__5121 (
            .O(N__21524),
            .I(N__21475));
    LocalMux I__5120 (
            .O(N__21519),
            .I(N__21475));
    Span4Mux_s2_v I__5119 (
            .O(N__21516),
            .I(N__21466));
    Span4Mux_h I__5118 (
            .O(N__21513),
            .I(N__21466));
    LocalMux I__5117 (
            .O(N__21506),
            .I(N__21466));
    Span4Mux_h I__5116 (
            .O(N__21503),
            .I(N__21466));
    InMux I__5115 (
            .O(N__21502),
            .I(N__21459));
    InMux I__5114 (
            .O(N__21499),
            .I(N__21459));
    InMux I__5113 (
            .O(N__21496),
            .I(N__21459));
    Span4Mux_h I__5112 (
            .O(N__21491),
            .I(N__21456));
    LocalMux I__5111 (
            .O(N__21486),
            .I(bu_rx_data_6));
    LocalMux I__5110 (
            .O(N__21483),
            .I(bu_rx_data_6));
    LocalMux I__5109 (
            .O(N__21480),
            .I(bu_rx_data_6));
    Odrv4 I__5108 (
            .O(N__21475),
            .I(bu_rx_data_6));
    Odrv4 I__5107 (
            .O(N__21466),
            .I(bu_rx_data_6));
    LocalMux I__5106 (
            .O(N__21459),
            .I(bu_rx_data_6));
    Odrv4 I__5105 (
            .O(N__21456),
            .I(bu_rx_data_6));
    InMux I__5104 (
            .O(N__21441),
            .I(N__21437));
    InMux I__5103 (
            .O(N__21440),
            .I(N__21433));
    LocalMux I__5102 (
            .O(N__21437),
            .I(N__21427));
    InMux I__5101 (
            .O(N__21436),
            .I(N__21424));
    LocalMux I__5100 (
            .O(N__21433),
            .I(N__21421));
    InMux I__5099 (
            .O(N__21432),
            .I(N__21418));
    CascadeMux I__5098 (
            .O(N__21431),
            .I(N__21415));
    InMux I__5097 (
            .O(N__21430),
            .I(N__21412));
    Span12Mux_s6_h I__5096 (
            .O(N__21427),
            .I(N__21409));
    LocalMux I__5095 (
            .O(N__21424),
            .I(N__21406));
    Span4Mux_s3_h I__5094 (
            .O(N__21421),
            .I(N__21401));
    LocalMux I__5093 (
            .O(N__21418),
            .I(N__21401));
    InMux I__5092 (
            .O(N__21415),
            .I(N__21398));
    LocalMux I__5091 (
            .O(N__21412),
            .I(bu_rx_data_i_4_4));
    Odrv12 I__5090 (
            .O(N__21409),
            .I(bu_rx_data_i_4_4));
    Odrv4 I__5089 (
            .O(N__21406),
            .I(bu_rx_data_i_4_4));
    Odrv4 I__5088 (
            .O(N__21401),
            .I(bu_rx_data_i_4_4));
    LocalMux I__5087 (
            .O(N__21398),
            .I(bu_rx_data_i_4_4));
    InMux I__5086 (
            .O(N__21387),
            .I(N__21380));
    InMux I__5085 (
            .O(N__21386),
            .I(N__21377));
    InMux I__5084 (
            .O(N__21385),
            .I(N__21374));
    InMux I__5083 (
            .O(N__21384),
            .I(N__21371));
    CascadeMux I__5082 (
            .O(N__21383),
            .I(N__21360));
    LocalMux I__5081 (
            .O(N__21380),
            .I(N__21349));
    LocalMux I__5080 (
            .O(N__21377),
            .I(N__21349));
    LocalMux I__5079 (
            .O(N__21374),
            .I(N__21346));
    LocalMux I__5078 (
            .O(N__21371),
            .I(N__21337));
    InMux I__5077 (
            .O(N__21370),
            .I(N__21332));
    InMux I__5076 (
            .O(N__21369),
            .I(N__21332));
    InMux I__5075 (
            .O(N__21368),
            .I(N__21329));
    InMux I__5074 (
            .O(N__21367),
            .I(N__21326));
    InMux I__5073 (
            .O(N__21366),
            .I(N__21317));
    InMux I__5072 (
            .O(N__21365),
            .I(N__21317));
    InMux I__5071 (
            .O(N__21364),
            .I(N__21317));
    InMux I__5070 (
            .O(N__21363),
            .I(N__21317));
    InMux I__5069 (
            .O(N__21360),
            .I(N__21308));
    InMux I__5068 (
            .O(N__21359),
            .I(N__21308));
    InMux I__5067 (
            .O(N__21358),
            .I(N__21308));
    InMux I__5066 (
            .O(N__21357),
            .I(N__21308));
    InMux I__5065 (
            .O(N__21356),
            .I(N__21303));
    InMux I__5064 (
            .O(N__21355),
            .I(N__21303));
    InMux I__5063 (
            .O(N__21354),
            .I(N__21300));
    Span4Mux_v I__5062 (
            .O(N__21349),
            .I(N__21289));
    Span4Mux_v I__5061 (
            .O(N__21346),
            .I(N__21289));
    InMux I__5060 (
            .O(N__21345),
            .I(N__21284));
    InMux I__5059 (
            .O(N__21344),
            .I(N__21284));
    InMux I__5058 (
            .O(N__21343),
            .I(N__21281));
    InMux I__5057 (
            .O(N__21342),
            .I(N__21274));
    InMux I__5056 (
            .O(N__21341),
            .I(N__21274));
    InMux I__5055 (
            .O(N__21340),
            .I(N__21274));
    Span4Mux_v I__5054 (
            .O(N__21337),
            .I(N__21271));
    LocalMux I__5053 (
            .O(N__21332),
            .I(N__21264));
    LocalMux I__5052 (
            .O(N__21329),
            .I(N__21264));
    LocalMux I__5051 (
            .O(N__21326),
            .I(N__21264));
    LocalMux I__5050 (
            .O(N__21317),
            .I(N__21255));
    LocalMux I__5049 (
            .O(N__21308),
            .I(N__21255));
    LocalMux I__5048 (
            .O(N__21303),
            .I(N__21255));
    LocalMux I__5047 (
            .O(N__21300),
            .I(N__21255));
    InMux I__5046 (
            .O(N__21299),
            .I(N__21251));
    InMux I__5045 (
            .O(N__21298),
            .I(N__21248));
    InMux I__5044 (
            .O(N__21297),
            .I(N__21243));
    InMux I__5043 (
            .O(N__21296),
            .I(N__21243));
    InMux I__5042 (
            .O(N__21295),
            .I(N__21240));
    InMux I__5041 (
            .O(N__21294),
            .I(N__21237));
    Span4Mux_h I__5040 (
            .O(N__21289),
            .I(N__21234));
    LocalMux I__5039 (
            .O(N__21284),
            .I(N__21227));
    LocalMux I__5038 (
            .O(N__21281),
            .I(N__21227));
    LocalMux I__5037 (
            .O(N__21274),
            .I(N__21227));
    Span4Mux_v I__5036 (
            .O(N__21271),
            .I(N__21220));
    Span4Mux_v I__5035 (
            .O(N__21264),
            .I(N__21220));
    Span4Mux_v I__5034 (
            .O(N__21255),
            .I(N__21220));
    InMux I__5033 (
            .O(N__21254),
            .I(N__21217));
    LocalMux I__5032 (
            .O(N__21251),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5031 (
            .O(N__21248),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5030 (
            .O(N__21243),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5029 (
            .O(N__21240),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5028 (
            .O(N__21237),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5027 (
            .O(N__21234),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5026 (
            .O(N__21227),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__5025 (
            .O(N__21220),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__5024 (
            .O(N__21217),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    CascadeMux I__5023 (
            .O(N__21198),
            .I(g0_3_4_cascade_));
    InMux I__5022 (
            .O(N__21195),
            .I(N__21192));
    LocalMux I__5021 (
            .O(N__21192),
            .I(N__21189));
    Span4Mux_h I__5020 (
            .O(N__21189),
            .I(N__21186));
    Odrv4 I__5019 (
            .O(N__21186),
            .I(g0_3_5));
    InMux I__5018 (
            .O(N__21183),
            .I(N__21180));
    LocalMux I__5017 (
            .O(N__21180),
            .I(\Lab_UT.dictrl.g1Z0Z_2 ));
    InMux I__5016 (
            .O(N__21177),
            .I(N__21174));
    LocalMux I__5015 (
            .O(N__21174),
            .I(N__21171));
    Odrv12 I__5014 (
            .O(N__21171),
            .I(N_12));
    CascadeMux I__5013 (
            .O(N__21168),
            .I(N__21164));
    InMux I__5012 (
            .O(N__21167),
            .I(N__21159));
    InMux I__5011 (
            .O(N__21164),
            .I(N__21159));
    LocalMux I__5010 (
            .O(N__21159),
            .I(N__21154));
    CascadeMux I__5009 (
            .O(N__21158),
            .I(N__21150));
    InMux I__5008 (
            .O(N__21157),
            .I(N__21142));
    Span4Mux_v I__5007 (
            .O(N__21154),
            .I(N__21139));
    InMux I__5006 (
            .O(N__21153),
            .I(N__21132));
    InMux I__5005 (
            .O(N__21150),
            .I(N__21132));
    InMux I__5004 (
            .O(N__21149),
            .I(N__21132));
    InMux I__5003 (
            .O(N__21148),
            .I(N__21129));
    CascadeMux I__5002 (
            .O(N__21147),
            .I(N__21126));
    CascadeMux I__5001 (
            .O(N__21146),
            .I(N__21122));
    InMux I__5000 (
            .O(N__21145),
            .I(N__21117));
    LocalMux I__4999 (
            .O(N__21142),
            .I(N__21108));
    Span4Mux_h I__4998 (
            .O(N__21139),
            .I(N__21108));
    LocalMux I__4997 (
            .O(N__21132),
            .I(N__21108));
    LocalMux I__4996 (
            .O(N__21129),
            .I(N__21108));
    InMux I__4995 (
            .O(N__21126),
            .I(N__21103));
    InMux I__4994 (
            .O(N__21125),
            .I(N__21103));
    InMux I__4993 (
            .O(N__21122),
            .I(N__21100));
    InMux I__4992 (
            .O(N__21121),
            .I(N__21095));
    InMux I__4991 (
            .O(N__21120),
            .I(N__21095));
    LocalMux I__4990 (
            .O(N__21117),
            .I(N__21088));
    Sp12to4 I__4989 (
            .O(N__21108),
            .I(N__21088));
    LocalMux I__4988 (
            .O(N__21103),
            .I(N__21088));
    LocalMux I__4987 (
            .O(N__21100),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    LocalMux I__4986 (
            .O(N__21095),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv12 I__4985 (
            .O(N__21088),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    InMux I__4984 (
            .O(N__21081),
            .I(N__21078));
    LocalMux I__4983 (
            .O(N__21078),
            .I(N__21074));
    InMux I__4982 (
            .O(N__21077),
            .I(N__21066));
    Span4Mux_v I__4981 (
            .O(N__21074),
            .I(N__21059));
    InMux I__4980 (
            .O(N__21073),
            .I(N__21048));
    InMux I__4979 (
            .O(N__21072),
            .I(N__21048));
    InMux I__4978 (
            .O(N__21071),
            .I(N__21048));
    InMux I__4977 (
            .O(N__21070),
            .I(N__21048));
    InMux I__4976 (
            .O(N__21069),
            .I(N__21048));
    LocalMux I__4975 (
            .O(N__21066),
            .I(N__21045));
    InMux I__4974 (
            .O(N__21065),
            .I(N__21040));
    InMux I__4973 (
            .O(N__21064),
            .I(N__21040));
    InMux I__4972 (
            .O(N__21063),
            .I(N__21032));
    InMux I__4971 (
            .O(N__21062),
            .I(N__21029));
    Span4Mux_h I__4970 (
            .O(N__21059),
            .I(N__21026));
    LocalMux I__4969 (
            .O(N__21048),
            .I(N__21021));
    Span4Mux_h I__4968 (
            .O(N__21045),
            .I(N__21021));
    LocalMux I__4967 (
            .O(N__21040),
            .I(N__21018));
    InMux I__4966 (
            .O(N__21039),
            .I(N__21013));
    InMux I__4965 (
            .O(N__21038),
            .I(N__21013));
    InMux I__4964 (
            .O(N__21037),
            .I(N__21006));
    InMux I__4963 (
            .O(N__21036),
            .I(N__21006));
    InMux I__4962 (
            .O(N__21035),
            .I(N__21006));
    LocalMux I__4961 (
            .O(N__21032),
            .I(bu_rx_data_4));
    LocalMux I__4960 (
            .O(N__21029),
            .I(bu_rx_data_4));
    Odrv4 I__4959 (
            .O(N__21026),
            .I(bu_rx_data_4));
    Odrv4 I__4958 (
            .O(N__21021),
            .I(bu_rx_data_4));
    Odrv4 I__4957 (
            .O(N__21018),
            .I(bu_rx_data_4));
    LocalMux I__4956 (
            .O(N__21013),
            .I(bu_rx_data_4));
    LocalMux I__4955 (
            .O(N__21006),
            .I(bu_rx_data_4));
    InMux I__4954 (
            .O(N__20991),
            .I(N__20988));
    LocalMux I__4953 (
            .O(N__20988),
            .I(\Lab_UT.dictrl.N_13 ));
    InMux I__4952 (
            .O(N__20985),
            .I(N__20981));
    InMux I__4951 (
            .O(N__20984),
            .I(N__20977));
    LocalMux I__4950 (
            .O(N__20981),
            .I(N__20974));
    InMux I__4949 (
            .O(N__20980),
            .I(N__20971));
    LocalMux I__4948 (
            .O(N__20977),
            .I(N__20959));
    Span4Mux_s1_h I__4947 (
            .O(N__20974),
            .I(N__20956));
    LocalMux I__4946 (
            .O(N__20971),
            .I(N__20953));
    InMux I__4945 (
            .O(N__20970),
            .I(N__20948));
    InMux I__4944 (
            .O(N__20969),
            .I(N__20948));
    InMux I__4943 (
            .O(N__20968),
            .I(N__20938));
    InMux I__4942 (
            .O(N__20967),
            .I(N__20938));
    InMux I__4941 (
            .O(N__20966),
            .I(N__20927));
    InMux I__4940 (
            .O(N__20965),
            .I(N__20927));
    InMux I__4939 (
            .O(N__20964),
            .I(N__20927));
    InMux I__4938 (
            .O(N__20963),
            .I(N__20927));
    InMux I__4937 (
            .O(N__20962),
            .I(N__20927));
    Span4Mux_v I__4936 (
            .O(N__20959),
            .I(N__20924));
    Span4Mux_h I__4935 (
            .O(N__20956),
            .I(N__20921));
    Span4Mux_s2_h I__4934 (
            .O(N__20953),
            .I(N__20916));
    LocalMux I__4933 (
            .O(N__20948),
            .I(N__20916));
    InMux I__4932 (
            .O(N__20947),
            .I(N__20905));
    InMux I__4931 (
            .O(N__20946),
            .I(N__20905));
    InMux I__4930 (
            .O(N__20945),
            .I(N__20905));
    InMux I__4929 (
            .O(N__20944),
            .I(N__20905));
    InMux I__4928 (
            .O(N__20943),
            .I(N__20905));
    LocalMux I__4927 (
            .O(N__20938),
            .I(bu_rx_data_5));
    LocalMux I__4926 (
            .O(N__20927),
            .I(bu_rx_data_5));
    Odrv4 I__4925 (
            .O(N__20924),
            .I(bu_rx_data_5));
    Odrv4 I__4924 (
            .O(N__20921),
            .I(bu_rx_data_5));
    Odrv4 I__4923 (
            .O(N__20916),
            .I(bu_rx_data_5));
    LocalMux I__4922 (
            .O(N__20905),
            .I(bu_rx_data_5));
    InMux I__4921 (
            .O(N__20892),
            .I(N__20889));
    LocalMux I__4920 (
            .O(N__20889),
            .I(N__20883));
    InMux I__4919 (
            .O(N__20888),
            .I(N__20880));
    InMux I__4918 (
            .O(N__20887),
            .I(N__20872));
    InMux I__4917 (
            .O(N__20886),
            .I(N__20869));
    Span4Mux_s3_v I__4916 (
            .O(N__20883),
            .I(N__20866));
    LocalMux I__4915 (
            .O(N__20880),
            .I(N__20861));
    InMux I__4914 (
            .O(N__20879),
            .I(N__20858));
    InMux I__4913 (
            .O(N__20878),
            .I(N__20848));
    InMux I__4912 (
            .O(N__20877),
            .I(N__20845));
    InMux I__4911 (
            .O(N__20876),
            .I(N__20840));
    InMux I__4910 (
            .O(N__20875),
            .I(N__20840));
    LocalMux I__4909 (
            .O(N__20872),
            .I(N__20837));
    LocalMux I__4908 (
            .O(N__20869),
            .I(N__20834));
    Span4Mux_v I__4907 (
            .O(N__20866),
            .I(N__20830));
    InMux I__4906 (
            .O(N__20865),
            .I(N__20825));
    InMux I__4905 (
            .O(N__20864),
            .I(N__20825));
    Span4Mux_v I__4904 (
            .O(N__20861),
            .I(N__20820));
    LocalMux I__4903 (
            .O(N__20858),
            .I(N__20820));
    InMux I__4902 (
            .O(N__20857),
            .I(N__20815));
    InMux I__4901 (
            .O(N__20856),
            .I(N__20815));
    InMux I__4900 (
            .O(N__20855),
            .I(N__20812));
    InMux I__4899 (
            .O(N__20854),
            .I(N__20809));
    InMux I__4898 (
            .O(N__20853),
            .I(N__20806));
    InMux I__4897 (
            .O(N__20852),
            .I(N__20803));
    InMux I__4896 (
            .O(N__20851),
            .I(N__20796));
    LocalMux I__4895 (
            .O(N__20848),
            .I(N__20793));
    LocalMux I__4894 (
            .O(N__20845),
            .I(N__20784));
    LocalMux I__4893 (
            .O(N__20840),
            .I(N__20784));
    Span12Mux_s0_v I__4892 (
            .O(N__20837),
            .I(N__20784));
    Sp12to4 I__4891 (
            .O(N__20834),
            .I(N__20784));
    CascadeMux I__4890 (
            .O(N__20833),
            .I(N__20781));
    Span4Mux_v I__4889 (
            .O(N__20830),
            .I(N__20774));
    LocalMux I__4888 (
            .O(N__20825),
            .I(N__20774));
    Span4Mux_h I__4887 (
            .O(N__20820),
            .I(N__20767));
    LocalMux I__4886 (
            .O(N__20815),
            .I(N__20767));
    LocalMux I__4885 (
            .O(N__20812),
            .I(N__20767));
    LocalMux I__4884 (
            .O(N__20809),
            .I(N__20760));
    LocalMux I__4883 (
            .O(N__20806),
            .I(N__20760));
    LocalMux I__4882 (
            .O(N__20803),
            .I(N__20760));
    InMux I__4881 (
            .O(N__20802),
            .I(N__20755));
    InMux I__4880 (
            .O(N__20801),
            .I(N__20755));
    InMux I__4879 (
            .O(N__20800),
            .I(N__20752));
    InMux I__4878 (
            .O(N__20799),
            .I(N__20749));
    LocalMux I__4877 (
            .O(N__20796),
            .I(N__20744));
    Span4Mux_v I__4876 (
            .O(N__20793),
            .I(N__20744));
    Span12Mux_v I__4875 (
            .O(N__20784),
            .I(N__20741));
    InMux I__4874 (
            .O(N__20781),
            .I(N__20738));
    InMux I__4873 (
            .O(N__20780),
            .I(N__20733));
    InMux I__4872 (
            .O(N__20779),
            .I(N__20733));
    Span4Mux_h I__4871 (
            .O(N__20774),
            .I(N__20730));
    Span4Mux_v I__4870 (
            .O(N__20767),
            .I(N__20723));
    Span4Mux_h I__4869 (
            .O(N__20760),
            .I(N__20723));
    LocalMux I__4868 (
            .O(N__20755),
            .I(N__20723));
    LocalMux I__4867 (
            .O(N__20752),
            .I(bu_rx_data_1));
    LocalMux I__4866 (
            .O(N__20749),
            .I(bu_rx_data_1));
    Odrv4 I__4865 (
            .O(N__20744),
            .I(bu_rx_data_1));
    Odrv12 I__4864 (
            .O(N__20741),
            .I(bu_rx_data_1));
    LocalMux I__4863 (
            .O(N__20738),
            .I(bu_rx_data_1));
    LocalMux I__4862 (
            .O(N__20733),
            .I(bu_rx_data_1));
    Odrv4 I__4861 (
            .O(N__20730),
            .I(bu_rx_data_1));
    Odrv4 I__4860 (
            .O(N__20723),
            .I(bu_rx_data_1));
    CascadeMux I__4859 (
            .O(N__20706),
            .I(N__20699));
    CascadeMux I__4858 (
            .O(N__20705),
            .I(N__20696));
    InMux I__4857 (
            .O(N__20704),
            .I(N__20693));
    InMux I__4856 (
            .O(N__20703),
            .I(N__20688));
    InMux I__4855 (
            .O(N__20702),
            .I(N__20688));
    InMux I__4854 (
            .O(N__20699),
            .I(N__20685));
    InMux I__4853 (
            .O(N__20696),
            .I(N__20682));
    LocalMux I__4852 (
            .O(N__20693),
            .I(N__20677));
    LocalMux I__4851 (
            .O(N__20688),
            .I(N__20677));
    LocalMux I__4850 (
            .O(N__20685),
            .I(N__20672));
    LocalMux I__4849 (
            .O(N__20682),
            .I(N__20672));
    Span4Mux_s3_v I__4848 (
            .O(N__20677),
            .I(N__20667));
    Span4Mux_s3_h I__4847 (
            .O(N__20672),
            .I(N__20667));
    Odrv4 I__4846 (
            .O(N__20667),
            .I(bu_rx_data_i_4_3_rep1));
    CascadeMux I__4845 (
            .O(N__20664),
            .I(N__20661));
    InMux I__4844 (
            .O(N__20661),
            .I(N__20657));
    InMux I__4843 (
            .O(N__20660),
            .I(N__20653));
    LocalMux I__4842 (
            .O(N__20657),
            .I(N__20648));
    InMux I__4841 (
            .O(N__20656),
            .I(N__20645));
    LocalMux I__4840 (
            .O(N__20653),
            .I(N__20642));
    InMux I__4839 (
            .O(N__20652),
            .I(N__20638));
    InMux I__4838 (
            .O(N__20651),
            .I(N__20633));
    Span4Mux_h I__4837 (
            .O(N__20648),
            .I(N__20629));
    LocalMux I__4836 (
            .O(N__20645),
            .I(N__20626));
    Span4Mux_h I__4835 (
            .O(N__20642),
            .I(N__20623));
    InMux I__4834 (
            .O(N__20641),
            .I(N__20620));
    LocalMux I__4833 (
            .O(N__20638),
            .I(N__20617));
    InMux I__4832 (
            .O(N__20637),
            .I(N__20612));
    InMux I__4831 (
            .O(N__20636),
            .I(N__20612));
    LocalMux I__4830 (
            .O(N__20633),
            .I(N__20609));
    InMux I__4829 (
            .O(N__20632),
            .I(N__20606));
    Odrv4 I__4828 (
            .O(N__20629),
            .I(bu_rx_data_i_4_2));
    Odrv12 I__4827 (
            .O(N__20626),
            .I(bu_rx_data_i_4_2));
    Odrv4 I__4826 (
            .O(N__20623),
            .I(bu_rx_data_i_4_2));
    LocalMux I__4825 (
            .O(N__20620),
            .I(bu_rx_data_i_4_2));
    Odrv4 I__4824 (
            .O(N__20617),
            .I(bu_rx_data_i_4_2));
    LocalMux I__4823 (
            .O(N__20612),
            .I(bu_rx_data_i_4_2));
    Odrv12 I__4822 (
            .O(N__20609),
            .I(bu_rx_data_i_4_2));
    LocalMux I__4821 (
            .O(N__20606),
            .I(bu_rx_data_i_4_2));
    InMux I__4820 (
            .O(N__20589),
            .I(N__20586));
    LocalMux I__4819 (
            .O(N__20586),
            .I(m46_i_0_a3_2));
    InMux I__4818 (
            .O(N__20583),
            .I(N__20578));
    InMux I__4817 (
            .O(N__20582),
            .I(N__20573));
    InMux I__4816 (
            .O(N__20581),
            .I(N__20573));
    LocalMux I__4815 (
            .O(N__20578),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__4814 (
            .O(N__20573),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__4813 (
            .O(N__20568),
            .I(N__20565));
    InMux I__4812 (
            .O(N__20565),
            .I(N__20559));
    InMux I__4811 (
            .O(N__20564),
            .I(N__20552));
    InMux I__4810 (
            .O(N__20563),
            .I(N__20552));
    InMux I__4809 (
            .O(N__20562),
            .I(N__20552));
    LocalMux I__4808 (
            .O(N__20559),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__4807 (
            .O(N__20552),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    InMux I__4806 (
            .O(N__20547),
            .I(N__20542));
    InMux I__4805 (
            .O(N__20546),
            .I(N__20537));
    InMux I__4804 (
            .O(N__20545),
            .I(N__20537));
    LocalMux I__4803 (
            .O(N__20542),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__4802 (
            .O(N__20537),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__4801 (
            .O(N__20532),
            .I(N__20526));
    InMux I__4800 (
            .O(N__20531),
            .I(N__20526));
    LocalMux I__4799 (
            .O(N__20526),
            .I(N__20523));
    Span4Mux_s2_h I__4798 (
            .O(N__20523),
            .I(N__20520));
    Odrv4 I__4797 (
            .O(N__20520),
            .I(\Lab_UT.dictrl.N_90 ));
    CascadeMux I__4796 (
            .O(N__20517),
            .I(\Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_ ));
    InMux I__4795 (
            .O(N__20514),
            .I(N__20511));
    LocalMux I__4794 (
            .O(N__20511),
            .I(N__20506));
    InMux I__4793 (
            .O(N__20510),
            .I(N__20501));
    InMux I__4792 (
            .O(N__20509),
            .I(N__20501));
    Span4Mux_v I__4791 (
            .O(N__20506),
            .I(N__20498));
    LocalMux I__4790 (
            .O(N__20501),
            .I(N__20495));
    Odrv4 I__4789 (
            .O(N__20498),
            .I(\Lab_UT.dictrl.N_119 ));
    Odrv12 I__4788 (
            .O(N__20495),
            .I(\Lab_UT.dictrl.N_119 ));
    CascadeMux I__4787 (
            .O(N__20490),
            .I(\Lab_UT.dictrl.N_139_cascade_ ));
    InMux I__4786 (
            .O(N__20487),
            .I(N__20482));
    InMux I__4785 (
            .O(N__20486),
            .I(N__20476));
    InMux I__4784 (
            .O(N__20485),
            .I(N__20476));
    LocalMux I__4783 (
            .O(N__20482),
            .I(N__20473));
    InMux I__4782 (
            .O(N__20481),
            .I(N__20470));
    LocalMux I__4781 (
            .O(N__20476),
            .I(N__20465));
    Span4Mux_v I__4780 (
            .O(N__20473),
            .I(N__20460));
    LocalMux I__4779 (
            .O(N__20470),
            .I(N__20460));
    InMux I__4778 (
            .O(N__20469),
            .I(N__20455));
    InMux I__4777 (
            .O(N__20468),
            .I(N__20455));
    Span4Mux_h I__4776 (
            .O(N__20465),
            .I(N__20452));
    Span4Mux_h I__4775 (
            .O(N__20460),
            .I(N__20449));
    LocalMux I__4774 (
            .O(N__20455),
            .I(N__20446));
    Odrv4 I__4773 (
            .O(N__20452),
            .I(\Lab_UT.dictrl.N_116_mux ));
    Odrv4 I__4772 (
            .O(N__20449),
            .I(\Lab_UT.dictrl.N_116_mux ));
    Odrv4 I__4771 (
            .O(N__20446),
            .I(\Lab_UT.dictrl.N_116_mux ));
    InMux I__4770 (
            .O(N__20439),
            .I(N__20436));
    LocalMux I__4769 (
            .O(N__20436),
            .I(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ));
    CascadeMux I__4768 (
            .O(N__20433),
            .I(N__20430));
    InMux I__4767 (
            .O(N__20430),
            .I(N__20427));
    LocalMux I__4766 (
            .O(N__20427),
            .I(N__20424));
    Span4Mux_s2_h I__4765 (
            .O(N__20424),
            .I(N__20421));
    Odrv4 I__4764 (
            .O(N__20421),
            .I(\Lab_UT.dictrl.g2_2 ));
    InMux I__4763 (
            .O(N__20418),
            .I(N__20415));
    LocalMux I__4762 (
            .O(N__20415),
            .I(N__20410));
    InMux I__4761 (
            .O(N__20414),
            .I(N__20407));
    InMux I__4760 (
            .O(N__20413),
            .I(N__20404));
    Span4Mux_s2_h I__4759 (
            .O(N__20410),
            .I(N__20401));
    LocalMux I__4758 (
            .O(N__20407),
            .I(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1 ));
    LocalMux I__4757 (
            .O(N__20404),
            .I(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1 ));
    Odrv4 I__4756 (
            .O(N__20401),
            .I(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1 ));
    InMux I__4755 (
            .O(N__20394),
            .I(N__20391));
    LocalMux I__4754 (
            .O(N__20391),
            .I(N__20388));
    Odrv4 I__4753 (
            .O(N__20388),
            .I(\Lab_UT.dictrl.N_5_1 ));
    InMux I__4752 (
            .O(N__20385),
            .I(N__20382));
    LocalMux I__4751 (
            .O(N__20382),
            .I(N__20379));
    Span4Mux_s2_h I__4750 (
            .O(N__20379),
            .I(N__20376));
    Odrv4 I__4749 (
            .O(N__20376),
            .I(\Lab_UT.dictrl.g2_0_0_0_0 ));
    CascadeMux I__4748 (
            .O(N__20373),
            .I(N__20363));
    CascadeMux I__4747 (
            .O(N__20372),
            .I(N__20360));
    InMux I__4746 (
            .O(N__20371),
            .I(N__20356));
    CascadeMux I__4745 (
            .O(N__20370),
            .I(N__20353));
    CascadeMux I__4744 (
            .O(N__20369),
            .I(N__20348));
    CascadeMux I__4743 (
            .O(N__20368),
            .I(N__20342));
    CascadeMux I__4742 (
            .O(N__20367),
            .I(N__20338));
    CascadeMux I__4741 (
            .O(N__20366),
            .I(N__20333));
    InMux I__4740 (
            .O(N__20363),
            .I(N__20329));
    InMux I__4739 (
            .O(N__20360),
            .I(N__20326));
    InMux I__4738 (
            .O(N__20359),
            .I(N__20323));
    LocalMux I__4737 (
            .O(N__20356),
            .I(N__20320));
    InMux I__4736 (
            .O(N__20353),
            .I(N__20317));
    InMux I__4735 (
            .O(N__20352),
            .I(N__20312));
    InMux I__4734 (
            .O(N__20351),
            .I(N__20312));
    InMux I__4733 (
            .O(N__20348),
            .I(N__20309));
    InMux I__4732 (
            .O(N__20347),
            .I(N__20306));
    CascadeMux I__4731 (
            .O(N__20346),
            .I(N__20301));
    InMux I__4730 (
            .O(N__20345),
            .I(N__20295));
    InMux I__4729 (
            .O(N__20342),
            .I(N__20295));
    InMux I__4728 (
            .O(N__20341),
            .I(N__20292));
    InMux I__4727 (
            .O(N__20338),
            .I(N__20287));
    InMux I__4726 (
            .O(N__20337),
            .I(N__20287));
    InMux I__4725 (
            .O(N__20336),
            .I(N__20282));
    InMux I__4724 (
            .O(N__20333),
            .I(N__20282));
    CascadeMux I__4723 (
            .O(N__20332),
            .I(N__20279));
    LocalMux I__4722 (
            .O(N__20329),
            .I(N__20274));
    LocalMux I__4721 (
            .O(N__20326),
            .I(N__20274));
    LocalMux I__4720 (
            .O(N__20323),
            .I(N__20265));
    Span4Mux_v I__4719 (
            .O(N__20320),
            .I(N__20265));
    LocalMux I__4718 (
            .O(N__20317),
            .I(N__20265));
    LocalMux I__4717 (
            .O(N__20312),
            .I(N__20265));
    LocalMux I__4716 (
            .O(N__20309),
            .I(N__20262));
    LocalMux I__4715 (
            .O(N__20306),
            .I(N__20259));
    InMux I__4714 (
            .O(N__20305),
            .I(N__20252));
    InMux I__4713 (
            .O(N__20304),
            .I(N__20252));
    InMux I__4712 (
            .O(N__20301),
            .I(N__20252));
    InMux I__4711 (
            .O(N__20300),
            .I(N__20249));
    LocalMux I__4710 (
            .O(N__20295),
            .I(N__20246));
    LocalMux I__4709 (
            .O(N__20292),
            .I(N__20241));
    LocalMux I__4708 (
            .O(N__20287),
            .I(N__20241));
    LocalMux I__4707 (
            .O(N__20282),
            .I(N__20238));
    InMux I__4706 (
            .O(N__20279),
            .I(N__20235));
    Span4Mux_v I__4705 (
            .O(N__20274),
            .I(N__20230));
    Span4Mux_v I__4704 (
            .O(N__20265),
            .I(N__20230));
    Span4Mux_s3_h I__4703 (
            .O(N__20262),
            .I(N__20221));
    Span4Mux_v I__4702 (
            .O(N__20259),
            .I(N__20221));
    LocalMux I__4701 (
            .O(N__20252),
            .I(N__20221));
    LocalMux I__4700 (
            .O(N__20249),
            .I(N__20221));
    Span4Mux_h I__4699 (
            .O(N__20246),
            .I(N__20218));
    Odrv12 I__4698 (
            .O(N__20241),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4697 (
            .O(N__20238),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4696 (
            .O(N__20235),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4695 (
            .O(N__20230),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4694 (
            .O(N__20221),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4693 (
            .O(N__20218),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    InMux I__4692 (
            .O(N__20205),
            .I(N__20202));
    LocalMux I__4691 (
            .O(N__20202),
            .I(N__20199));
    Span4Mux_s2_h I__4690 (
            .O(N__20199),
            .I(N__20196));
    Odrv4 I__4689 (
            .O(N__20196),
            .I(\Lab_UT.dictrl.N_103_0_0_0 ));
    InMux I__4688 (
            .O(N__20193),
            .I(N__20190));
    LocalMux I__4687 (
            .O(N__20190),
            .I(\Lab_UT.dictrl.N_1302_1_0_0 ));
    CascadeMux I__4686 (
            .O(N__20187),
            .I(\Lab_UT.dictrl.N_119_0_0_0_cascade_ ));
    InMux I__4685 (
            .O(N__20184),
            .I(N__20169));
    InMux I__4684 (
            .O(N__20183),
            .I(N__20169));
    InMux I__4683 (
            .O(N__20182),
            .I(N__20165));
    InMux I__4682 (
            .O(N__20181),
            .I(N__20160));
    InMux I__4681 (
            .O(N__20180),
            .I(N__20160));
    CascadeMux I__4680 (
            .O(N__20179),
            .I(N__20155));
    CascadeMux I__4679 (
            .O(N__20178),
            .I(N__20152));
    CascadeMux I__4678 (
            .O(N__20177),
            .I(N__20148));
    InMux I__4677 (
            .O(N__20176),
            .I(N__20145));
    InMux I__4676 (
            .O(N__20175),
            .I(N__20142));
    CascadeMux I__4675 (
            .O(N__20174),
            .I(N__20138));
    LocalMux I__4674 (
            .O(N__20169),
            .I(N__20135));
    InMux I__4673 (
            .O(N__20168),
            .I(N__20125));
    LocalMux I__4672 (
            .O(N__20165),
            .I(N__20122));
    LocalMux I__4671 (
            .O(N__20160),
            .I(N__20119));
    InMux I__4670 (
            .O(N__20159),
            .I(N__20113));
    InMux I__4669 (
            .O(N__20158),
            .I(N__20113));
    InMux I__4668 (
            .O(N__20155),
            .I(N__20104));
    InMux I__4667 (
            .O(N__20152),
            .I(N__20104));
    InMux I__4666 (
            .O(N__20151),
            .I(N__20104));
    InMux I__4665 (
            .O(N__20148),
            .I(N__20104));
    LocalMux I__4664 (
            .O(N__20145),
            .I(N__20099));
    LocalMux I__4663 (
            .O(N__20142),
            .I(N__20099));
    InMux I__4662 (
            .O(N__20141),
            .I(N__20096));
    InMux I__4661 (
            .O(N__20138),
            .I(N__20092));
    Span4Mux_s3_h I__4660 (
            .O(N__20135),
            .I(N__20089));
    InMux I__4659 (
            .O(N__20134),
            .I(N__20078));
    InMux I__4658 (
            .O(N__20133),
            .I(N__20078));
    InMux I__4657 (
            .O(N__20132),
            .I(N__20078));
    InMux I__4656 (
            .O(N__20131),
            .I(N__20078));
    InMux I__4655 (
            .O(N__20130),
            .I(N__20078));
    InMux I__4654 (
            .O(N__20129),
            .I(N__20073));
    InMux I__4653 (
            .O(N__20128),
            .I(N__20073));
    LocalMux I__4652 (
            .O(N__20125),
            .I(N__20066));
    Span4Mux_s3_h I__4651 (
            .O(N__20122),
            .I(N__20066));
    Span4Mux_s3_h I__4650 (
            .O(N__20119),
            .I(N__20066));
    InMux I__4649 (
            .O(N__20118),
            .I(N__20063));
    LocalMux I__4648 (
            .O(N__20113),
            .I(N__20054));
    LocalMux I__4647 (
            .O(N__20104),
            .I(N__20054));
    Span12Mux_s9_v I__4646 (
            .O(N__20099),
            .I(N__20054));
    LocalMux I__4645 (
            .O(N__20096),
            .I(N__20054));
    InMux I__4644 (
            .O(N__20095),
            .I(N__20051));
    LocalMux I__4643 (
            .O(N__20092),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__4642 (
            .O(N__20089),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4641 (
            .O(N__20078),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4640 (
            .O(N__20073),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__4639 (
            .O(N__20066),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4638 (
            .O(N__20063),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv12 I__4637 (
            .O(N__20054),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4636 (
            .O(N__20051),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    CascadeMux I__4635 (
            .O(N__20034),
            .I(N__20031));
    InMux I__4634 (
            .O(N__20031),
            .I(N__20025));
    InMux I__4633 (
            .O(N__20030),
            .I(N__20025));
    LocalMux I__4632 (
            .O(N__20025),
            .I(N__20022));
    Span4Mux_h I__4631 (
            .O(N__20022),
            .I(N__20019));
    Odrv4 I__4630 (
            .O(N__20019),
            .I(\Lab_UT.dictrl.g1Z0Z_4 ));
    CascadeMux I__4629 (
            .O(N__20016),
            .I(Lab_UT_dictrl_next_state_3_cascade_));
    InMux I__4628 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__4627 (
            .O(N__20010),
            .I(\Lab_UT.dictrl.state_ret_12_RNOZ0Z_3 ));
    InMux I__4626 (
            .O(N__20007),
            .I(N__20004));
    LocalMux I__4625 (
            .O(N__20004),
            .I(\Lab_UT.dictrl.next_state_0_0_2 ));
    InMux I__4624 (
            .O(N__20001),
            .I(N__19998));
    LocalMux I__4623 (
            .O(N__19998),
            .I(\Lab_UT.dictrl.state_ret_12_RNOZ0Z_4 ));
    InMux I__4622 (
            .O(N__19995),
            .I(N__19992));
    LocalMux I__4621 (
            .O(N__19992),
            .I(\Lab_UT.dictrl.state_ret_12and_a0_1 ));
    CascadeMux I__4620 (
            .O(N__19989),
            .I(N__19985));
    CascadeMux I__4619 (
            .O(N__19988),
            .I(N__19982));
    InMux I__4618 (
            .O(N__19985),
            .I(N__19974));
    InMux I__4617 (
            .O(N__19982),
            .I(N__19974));
    InMux I__4616 (
            .O(N__19981),
            .I(N__19974));
    LocalMux I__4615 (
            .O(N__19974),
            .I(N__19969));
    InMux I__4614 (
            .O(N__19973),
            .I(N__19966));
    InMux I__4613 (
            .O(N__19972),
            .I(N__19963));
    Span4Mux_s3_h I__4612 (
            .O(N__19969),
            .I(N__19958));
    LocalMux I__4611 (
            .O(N__19966),
            .I(N__19958));
    LocalMux I__4610 (
            .O(N__19963),
            .I(N__19955));
    Odrv4 I__4609 (
            .O(N__19958),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    Odrv4 I__4608 (
            .O(N__19955),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    CascadeMux I__4607 (
            .O(N__19950),
            .I(\Lab_UT.dictrl.state_ret_12and_0_0_cascade_ ));
    InMux I__4606 (
            .O(N__19947),
            .I(N__19939));
    InMux I__4605 (
            .O(N__19946),
            .I(N__19932));
    InMux I__4604 (
            .O(N__19945),
            .I(N__19932));
    InMux I__4603 (
            .O(N__19944),
            .I(N__19932));
    InMux I__4602 (
            .O(N__19943),
            .I(N__19929));
    InMux I__4601 (
            .O(N__19942),
            .I(N__19926));
    LocalMux I__4600 (
            .O(N__19939),
            .I(N__19923));
    LocalMux I__4599 (
            .O(N__19932),
            .I(N__19920));
    LocalMux I__4598 (
            .O(N__19929),
            .I(N__19917));
    LocalMux I__4597 (
            .O(N__19926),
            .I(N__19914));
    Span4Mux_h I__4596 (
            .O(N__19923),
            .I(N__19911));
    Odrv12 I__4595 (
            .O(N__19920),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    Odrv4 I__4594 (
            .O(N__19917),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    Odrv4 I__4593 (
            .O(N__19914),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    Odrv4 I__4592 (
            .O(N__19911),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    CascadeMux I__4591 (
            .O(N__19902),
            .I(N__19896));
    CascadeMux I__4590 (
            .O(N__19901),
            .I(N__19890));
    InMux I__4589 (
            .O(N__19900),
            .I(N__19884));
    InMux I__4588 (
            .O(N__19899),
            .I(N__19879));
    InMux I__4587 (
            .O(N__19896),
            .I(N__19876));
    InMux I__4586 (
            .O(N__19895),
            .I(N__19873));
    InMux I__4585 (
            .O(N__19894),
            .I(N__19870));
    CascadeMux I__4584 (
            .O(N__19893),
            .I(N__19867));
    InMux I__4583 (
            .O(N__19890),
            .I(N__19860));
    InMux I__4582 (
            .O(N__19889),
            .I(N__19860));
    InMux I__4581 (
            .O(N__19888),
            .I(N__19860));
    InMux I__4580 (
            .O(N__19887),
            .I(N__19857));
    LocalMux I__4579 (
            .O(N__19884),
            .I(N__19854));
    InMux I__4578 (
            .O(N__19883),
            .I(N__19851));
    InMux I__4577 (
            .O(N__19882),
            .I(N__19848));
    LocalMux I__4576 (
            .O(N__19879),
            .I(N__19845));
    LocalMux I__4575 (
            .O(N__19876),
            .I(N__19838));
    LocalMux I__4574 (
            .O(N__19873),
            .I(N__19838));
    LocalMux I__4573 (
            .O(N__19870),
            .I(N__19838));
    InMux I__4572 (
            .O(N__19867),
            .I(N__19835));
    LocalMux I__4571 (
            .O(N__19860),
            .I(N__19832));
    LocalMux I__4570 (
            .O(N__19857),
            .I(N__19829));
    Span4Mux_v I__4569 (
            .O(N__19854),
            .I(N__19822));
    LocalMux I__4568 (
            .O(N__19851),
            .I(N__19822));
    LocalMux I__4567 (
            .O(N__19848),
            .I(N__19822));
    Span4Mux_v I__4566 (
            .O(N__19845),
            .I(N__19817));
    Span4Mux_v I__4565 (
            .O(N__19838),
            .I(N__19817));
    LocalMux I__4564 (
            .O(N__19835),
            .I(N__19814));
    Span4Mux_h I__4563 (
            .O(N__19832),
            .I(N__19807));
    Span4Mux_v I__4562 (
            .O(N__19829),
            .I(N__19807));
    Span4Mux_v I__4561 (
            .O(N__19822),
            .I(N__19807));
    Odrv4 I__4560 (
            .O(N__19817),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv12 I__4559 (
            .O(N__19814),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    Odrv4 I__4558 (
            .O(N__19807),
            .I(\Lab_UT.dictrl.state_3_rep2 ));
    InMux I__4557 (
            .O(N__19800),
            .I(N__19796));
    InMux I__4556 (
            .O(N__19799),
            .I(N__19793));
    LocalMux I__4555 (
            .O(N__19796),
            .I(N__19790));
    LocalMux I__4554 (
            .O(N__19793),
            .I(N__19785));
    Span4Mux_v I__4553 (
            .O(N__19790),
            .I(N__19782));
    CascadeMux I__4552 (
            .O(N__19789),
            .I(N__19778));
    InMux I__4551 (
            .O(N__19788),
            .I(N__19771));
    Span4Mux_h I__4550 (
            .O(N__19785),
            .I(N__19766));
    Span4Mux_v I__4549 (
            .O(N__19782),
            .I(N__19766));
    InMux I__4548 (
            .O(N__19781),
            .I(N__19755));
    InMux I__4547 (
            .O(N__19778),
            .I(N__19755));
    InMux I__4546 (
            .O(N__19777),
            .I(N__19755));
    InMux I__4545 (
            .O(N__19776),
            .I(N__19755));
    InMux I__4544 (
            .O(N__19775),
            .I(N__19755));
    InMux I__4543 (
            .O(N__19774),
            .I(N__19752));
    LocalMux I__4542 (
            .O(N__19771),
            .I(N__19749));
    Odrv4 I__4541 (
            .O(N__19766),
            .I(buart__rx_bitcount_3));
    LocalMux I__4540 (
            .O(N__19755),
            .I(buart__rx_bitcount_3));
    LocalMux I__4539 (
            .O(N__19752),
            .I(buart__rx_bitcount_3));
    Odrv4 I__4538 (
            .O(N__19749),
            .I(buart__rx_bitcount_3));
    InMux I__4537 (
            .O(N__19740),
            .I(N__19737));
    LocalMux I__4536 (
            .O(N__19737),
            .I(N__19733));
    InMux I__4535 (
            .O(N__19736),
            .I(N__19730));
    Span4Mux_h I__4534 (
            .O(N__19733),
            .I(N__19727));
    LocalMux I__4533 (
            .O(N__19730),
            .I(N__19722));
    Span4Mux_v I__4532 (
            .O(N__19727),
            .I(N__19719));
    InMux I__4531 (
            .O(N__19726),
            .I(N__19714));
    InMux I__4530 (
            .O(N__19725),
            .I(N__19714));
    Span4Mux_v I__4529 (
            .O(N__19722),
            .I(N__19711));
    Odrv4 I__4528 (
            .O(N__19719),
            .I(buart__rx_valid_3));
    LocalMux I__4527 (
            .O(N__19714),
            .I(buart__rx_valid_3));
    Odrv4 I__4526 (
            .O(N__19711),
            .I(buart__rx_valid_3));
    InMux I__4525 (
            .O(N__19704),
            .I(N__19693));
    InMux I__4524 (
            .O(N__19703),
            .I(N__19693));
    InMux I__4523 (
            .O(N__19702),
            .I(N__19693));
    InMux I__4522 (
            .O(N__19701),
            .I(N__19690));
    InMux I__4521 (
            .O(N__19700),
            .I(N__19687));
    LocalMux I__4520 (
            .O(N__19693),
            .I(N__19684));
    LocalMux I__4519 (
            .O(N__19690),
            .I(N__19681));
    LocalMux I__4518 (
            .O(N__19687),
            .I(N__19678));
    Span4Mux_h I__4517 (
            .O(N__19684),
            .I(N__19673));
    Span4Mux_h I__4516 (
            .O(N__19681),
            .I(N__19670));
    Span4Mux_h I__4515 (
            .O(N__19678),
            .I(N__19667));
    InMux I__4514 (
            .O(N__19677),
            .I(N__19664));
    InMux I__4513 (
            .O(N__19676),
            .I(N__19661));
    Odrv4 I__4512 (
            .O(N__19673),
            .I(Lab_UT_dictrl_next_state_3));
    Odrv4 I__4511 (
            .O(N__19670),
            .I(Lab_UT_dictrl_next_state_3));
    Odrv4 I__4510 (
            .O(N__19667),
            .I(Lab_UT_dictrl_next_state_3));
    LocalMux I__4509 (
            .O(N__19664),
            .I(Lab_UT_dictrl_next_state_3));
    LocalMux I__4508 (
            .O(N__19661),
            .I(Lab_UT_dictrl_next_state_3));
    CascadeMux I__4507 (
            .O(N__19650),
            .I(bu_rx_data_rdy_cascade_));
    IoInMux I__4506 (
            .O(N__19647),
            .I(N__19641));
    InMux I__4505 (
            .O(N__19646),
            .I(N__19635));
    InMux I__4504 (
            .O(N__19645),
            .I(N__19630));
    InMux I__4503 (
            .O(N__19644),
            .I(N__19630));
    LocalMux I__4502 (
            .O(N__19641),
            .I(N__19627));
    InMux I__4501 (
            .O(N__19640),
            .I(N__19620));
    InMux I__4500 (
            .O(N__19639),
            .I(N__19620));
    InMux I__4499 (
            .O(N__19638),
            .I(N__19620));
    LocalMux I__4498 (
            .O(N__19635),
            .I(N__19617));
    LocalMux I__4497 (
            .O(N__19630),
            .I(N__19614));
    Span4Mux_s2_h I__4496 (
            .O(N__19627),
            .I(N__19611));
    LocalMux I__4495 (
            .O(N__19620),
            .I(N__19608));
    Span4Mux_h I__4494 (
            .O(N__19617),
            .I(N__19605));
    Span4Mux_v I__4493 (
            .O(N__19614),
            .I(N__19600));
    Span4Mux_h I__4492 (
            .O(N__19611),
            .I(N__19600));
    Odrv12 I__4491 (
            .O(N__19608),
            .I(rst));
    Odrv4 I__4490 (
            .O(N__19605),
            .I(rst));
    Odrv4 I__4489 (
            .O(N__19600),
            .I(rst));
    InMux I__4488 (
            .O(N__19593),
            .I(N__19590));
    LocalMux I__4487 (
            .O(N__19590),
            .I(N__19587));
    Span4Mux_v I__4486 (
            .O(N__19587),
            .I(N__19583));
    InMux I__4485 (
            .O(N__19586),
            .I(N__19580));
    Odrv4 I__4484 (
            .O(N__19583),
            .I(\Lab_UT.dictrl.N_119_mux ));
    LocalMux I__4483 (
            .O(N__19580),
            .I(\Lab_UT.dictrl.N_119_mux ));
    CascadeMux I__4482 (
            .O(N__19575),
            .I(\Lab_UT.dictrl.i9_mux_cascade_ ));
    InMux I__4481 (
            .O(N__19572),
            .I(N__19568));
    InMux I__4480 (
            .O(N__19571),
            .I(N__19565));
    LocalMux I__4479 (
            .O(N__19568),
            .I(N__19562));
    LocalMux I__4478 (
            .O(N__19565),
            .I(N__19559));
    Odrv12 I__4477 (
            .O(N__19562),
            .I(\Lab_UT.dictrl.N_94 ));
    Odrv12 I__4476 (
            .O(N__19559),
            .I(\Lab_UT.dictrl.N_94 ));
    CascadeMux I__4475 (
            .O(N__19554),
            .I(N__19551));
    InMux I__4474 (
            .O(N__19551),
            .I(N__19548));
    LocalMux I__4473 (
            .O(N__19548),
            .I(N__19542));
    InMux I__4472 (
            .O(N__19547),
            .I(N__19539));
    InMux I__4471 (
            .O(N__19546),
            .I(N__19536));
    InMux I__4470 (
            .O(N__19545),
            .I(N__19533));
    Span4Mux_v I__4469 (
            .O(N__19542),
            .I(N__19526));
    LocalMux I__4468 (
            .O(N__19539),
            .I(N__19526));
    LocalMux I__4467 (
            .O(N__19536),
            .I(N__19526));
    LocalMux I__4466 (
            .O(N__19533),
            .I(N__19523));
    Span4Mux_v I__4465 (
            .O(N__19526),
            .I(N__19520));
    Span4Mux_s1_h I__4464 (
            .O(N__19523),
            .I(N__19517));
    Odrv4 I__4463 (
            .O(N__19520),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    Odrv4 I__4462 (
            .O(N__19517),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    CascadeMux I__4461 (
            .O(N__19512),
            .I(\Lab_UT.dictrl.N_107_mux_cascade_ ));
    InMux I__4460 (
            .O(N__19509),
            .I(N__19506));
    LocalMux I__4459 (
            .O(N__19506),
            .I(m89_am));
    CascadeMux I__4458 (
            .O(N__19503),
            .I(N__19499));
    InMux I__4457 (
            .O(N__19502),
            .I(N__19491));
    InMux I__4456 (
            .O(N__19499),
            .I(N__19491));
    InMux I__4455 (
            .O(N__19498),
            .I(N__19491));
    LocalMux I__4454 (
            .O(N__19491),
            .I(N__19488));
    Span4Mux_v I__4453 (
            .O(N__19488),
            .I(N__19484));
    InMux I__4452 (
            .O(N__19487),
            .I(N__19481));
    Sp12to4 I__4451 (
            .O(N__19484),
            .I(N__19478));
    LocalMux I__4450 (
            .O(N__19481),
            .I(buart__rx_hh_0));
    Odrv12 I__4449 (
            .O(N__19478),
            .I(buart__rx_hh_0));
    InMux I__4448 (
            .O(N__19473),
            .I(N__19463));
    InMux I__4447 (
            .O(N__19472),
            .I(N__19463));
    InMux I__4446 (
            .O(N__19471),
            .I(N__19456));
    InMux I__4445 (
            .O(N__19470),
            .I(N__19456));
    InMux I__4444 (
            .O(N__19469),
            .I(N__19456));
    CascadeMux I__4443 (
            .O(N__19468),
            .I(N__19453));
    LocalMux I__4442 (
            .O(N__19463),
            .I(N__19448));
    LocalMux I__4441 (
            .O(N__19456),
            .I(N__19445));
    InMux I__4440 (
            .O(N__19453),
            .I(N__19438));
    InMux I__4439 (
            .O(N__19452),
            .I(N__19438));
    InMux I__4438 (
            .O(N__19451),
            .I(N__19438));
    Span4Mux_h I__4437 (
            .O(N__19448),
            .I(N__19433));
    Span4Mux_v I__4436 (
            .O(N__19445),
            .I(N__19433));
    LocalMux I__4435 (
            .O(N__19438),
            .I(N__19430));
    Span4Mux_v I__4434 (
            .O(N__19433),
            .I(N__19425));
    Span4Mux_v I__4433 (
            .O(N__19430),
            .I(N__19425));
    Sp12to4 I__4432 (
            .O(N__19425),
            .I(N__19422));
    Odrv12 I__4431 (
            .O(N__19422),
            .I(buart__rx_hh_1));
    InMux I__4430 (
            .O(N__19419),
            .I(N__19407));
    InMux I__4429 (
            .O(N__19418),
            .I(N__19407));
    InMux I__4428 (
            .O(N__19417),
            .I(N__19407));
    InMux I__4427 (
            .O(N__19416),
            .I(N__19407));
    LocalMux I__4426 (
            .O(N__19407),
            .I(\Lab_UT.dictrl.N_102_mux ));
    InMux I__4425 (
            .O(N__19404),
            .I(N__19396));
    InMux I__4424 (
            .O(N__19403),
            .I(N__19396));
    InMux I__4423 (
            .O(N__19402),
            .I(N__19393));
    InMux I__4422 (
            .O(N__19401),
            .I(N__19390));
    LocalMux I__4421 (
            .O(N__19396),
            .I(N__19385));
    LocalMux I__4420 (
            .O(N__19393),
            .I(N__19385));
    LocalMux I__4419 (
            .O(N__19390),
            .I(buart__rx_N_27_0_i));
    Odrv4 I__4418 (
            .O(N__19385),
            .I(buart__rx_N_27_0_i));
    CascadeMux I__4417 (
            .O(N__19380),
            .I(buart__rx_startbit_cascade_));
    InMux I__4416 (
            .O(N__19377),
            .I(N__19373));
    InMux I__4415 (
            .O(N__19376),
            .I(N__19367));
    LocalMux I__4414 (
            .O(N__19373),
            .I(N__19364));
    InMux I__4413 (
            .O(N__19372),
            .I(N__19357));
    InMux I__4412 (
            .O(N__19371),
            .I(N__19357));
    InMux I__4411 (
            .O(N__19370),
            .I(N__19357));
    LocalMux I__4410 (
            .O(N__19367),
            .I(buart__rx_bitcount_0));
    Odrv4 I__4409 (
            .O(N__19364),
            .I(buart__rx_bitcount_0));
    LocalMux I__4408 (
            .O(N__19357),
            .I(buart__rx_bitcount_0));
    CEMux I__4407 (
            .O(N__19350),
            .I(N__19346));
    CEMux I__4406 (
            .O(N__19349),
            .I(N__19342));
    LocalMux I__4405 (
            .O(N__19346),
            .I(N__19339));
    CEMux I__4404 (
            .O(N__19345),
            .I(N__19336));
    LocalMux I__4403 (
            .O(N__19342),
            .I(N__19333));
    Span4Mux_h I__4402 (
            .O(N__19339),
            .I(N__19330));
    LocalMux I__4401 (
            .O(N__19336),
            .I(N__19327));
    Odrv12 I__4400 (
            .O(N__19333),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__4399 (
            .O(N__19330),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__4398 (
            .O(N__19327),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__4397 (
            .O(N__19320),
            .I(N__19317));
    LocalMux I__4396 (
            .O(N__19317),
            .I(N__19314));
    Span4Mux_h I__4395 (
            .O(N__19314),
            .I(N__19311));
    Odrv4 I__4394 (
            .O(N__19311),
            .I(\Lab_UT.dictrl.i9_mux_0_0 ));
    InMux I__4393 (
            .O(N__19308),
            .I(N__19305));
    LocalMux I__4392 (
            .O(N__19305),
            .I(N__19302));
    Span4Mux_v I__4391 (
            .O(N__19302),
            .I(N__19299));
    Odrv4 I__4390 (
            .O(N__19299),
            .I(\Lab_UT.dictrl.N_94_0_0 ));
    CascadeMux I__4389 (
            .O(N__19296),
            .I(\Lab_UT.dictrl.N_2000_0_0_cascade_ ));
    InMux I__4388 (
            .O(N__19293),
            .I(N__19285));
    InMux I__4387 (
            .O(N__19292),
            .I(N__19285));
    InMux I__4386 (
            .O(N__19291),
            .I(N__19280));
    InMux I__4385 (
            .O(N__19290),
            .I(N__19280));
    LocalMux I__4384 (
            .O(N__19285),
            .I(N__19274));
    LocalMux I__4383 (
            .O(N__19280),
            .I(N__19274));
    InMux I__4382 (
            .O(N__19279),
            .I(N__19271));
    Span4Mux_v I__4381 (
            .O(N__19274),
            .I(N__19268));
    LocalMux I__4380 (
            .O(N__19271),
            .I(N__19265));
    Odrv4 I__4379 (
            .O(N__19268),
            .I(\Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3 ));
    Odrv12 I__4378 (
            .O(N__19265),
            .I(\Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3 ));
    InMux I__4377 (
            .O(N__19260),
            .I(N__19247));
    InMux I__4376 (
            .O(N__19259),
            .I(N__19247));
    InMux I__4375 (
            .O(N__19258),
            .I(N__19247));
    InMux I__4374 (
            .O(N__19257),
            .I(N__19247));
    InMux I__4373 (
            .O(N__19256),
            .I(N__19244));
    LocalMux I__4372 (
            .O(N__19247),
            .I(N__19239));
    LocalMux I__4371 (
            .O(N__19244),
            .I(N__19239));
    Odrv12 I__4370 (
            .O(N__19239),
            .I(\Lab_UT.dictrl.N_121_mux ));
    InMux I__4369 (
            .O(N__19236),
            .I(N__19233));
    LocalMux I__4368 (
            .O(N__19233),
            .I(N__19230));
    Span4Mux_h I__4367 (
            .O(N__19230),
            .I(N__19227));
    Span4Mux_v I__4366 (
            .O(N__19227),
            .I(N__19224));
    Odrv4 I__4365 (
            .O(N__19224),
            .I(\Lab_UT.dictrl.N_83 ));
    CascadeMux I__4364 (
            .O(N__19221),
            .I(\Lab_UT.dictrl.N_194_cascade_ ));
    IoInMux I__4363 (
            .O(N__19218),
            .I(N__19215));
    LocalMux I__4362 (
            .O(N__19215),
            .I(N__19212));
    IoSpan4Mux I__4361 (
            .O(N__19212),
            .I(N__19209));
    Span4Mux_s2_v I__4360 (
            .O(N__19209),
            .I(N__19206));
    Sp12to4 I__4359 (
            .O(N__19206),
            .I(N__19203));
    Odrv12 I__4358 (
            .O(N__19203),
            .I(buart__rx_sample));
    CascadeMux I__4357 (
            .O(N__19200),
            .I(N__19194));
    InMux I__4356 (
            .O(N__19199),
            .I(N__19187));
    InMux I__4355 (
            .O(N__19198),
            .I(N__19187));
    InMux I__4354 (
            .O(N__19197),
            .I(N__19187));
    InMux I__4353 (
            .O(N__19194),
            .I(N__19183));
    LocalMux I__4352 (
            .O(N__19187),
            .I(N__19180));
    InMux I__4351 (
            .O(N__19186),
            .I(N__19177));
    LocalMux I__4350 (
            .O(N__19183),
            .I(N__19172));
    Span4Mux_v I__4349 (
            .O(N__19180),
            .I(N__19172));
    LocalMux I__4348 (
            .O(N__19177),
            .I(buart__rx_bitcount_2));
    Odrv4 I__4347 (
            .O(N__19172),
            .I(buart__rx_bitcount_2));
    CascadeMux I__4346 (
            .O(N__19167),
            .I(N__19162));
    CascadeMux I__4345 (
            .O(N__19166),
            .I(N__19158));
    InMux I__4344 (
            .O(N__19165),
            .I(N__19151));
    InMux I__4343 (
            .O(N__19162),
            .I(N__19151));
    InMux I__4342 (
            .O(N__19161),
            .I(N__19151));
    InMux I__4341 (
            .O(N__19158),
            .I(N__19148));
    LocalMux I__4340 (
            .O(N__19151),
            .I(N__19144));
    LocalMux I__4339 (
            .O(N__19148),
            .I(N__19141));
    InMux I__4338 (
            .O(N__19147),
            .I(N__19138));
    Span4Mux_v I__4337 (
            .O(N__19144),
            .I(N__19135));
    Odrv4 I__4336 (
            .O(N__19141),
            .I(buart__rx_bitcount_1));
    LocalMux I__4335 (
            .O(N__19138),
            .I(buart__rx_bitcount_1));
    Odrv4 I__4334 (
            .O(N__19135),
            .I(buart__rx_bitcount_1));
    CascadeMux I__4333 (
            .O(N__19128),
            .I(N__19123));
    InMux I__4332 (
            .O(N__19127),
            .I(N__19115));
    InMux I__4331 (
            .O(N__19126),
            .I(N__19115));
    InMux I__4330 (
            .O(N__19123),
            .I(N__19115));
    CascadeMux I__4329 (
            .O(N__19122),
            .I(N__19112));
    LocalMux I__4328 (
            .O(N__19115),
            .I(N__19109));
    InMux I__4327 (
            .O(N__19112),
            .I(N__19106));
    Span4Mux_s2_h I__4326 (
            .O(N__19109),
            .I(N__19103));
    LocalMux I__4325 (
            .O(N__19106),
            .I(buart__rx_bitcount_4));
    Odrv4 I__4324 (
            .O(N__19103),
            .I(buart__rx_bitcount_4));
    InMux I__4323 (
            .O(N__19098),
            .I(N__19095));
    LocalMux I__4322 (
            .O(N__19095),
            .I(m89_bm));
    InMux I__4321 (
            .O(N__19092),
            .I(N__19089));
    LocalMux I__4320 (
            .O(N__19089),
            .I(N__19086));
    Odrv4 I__4319 (
            .O(N__19086),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__4318 (
            .O(N__19083),
            .I(buart__rx_N_27_0_i_cascade_));
    InMux I__4317 (
            .O(N__19080),
            .I(N__19072));
    InMux I__4316 (
            .O(N__19079),
            .I(N__19072));
    CascadeMux I__4315 (
            .O(N__19078),
            .I(N__19069));
    CascadeMux I__4314 (
            .O(N__19077),
            .I(N__19065));
    LocalMux I__4313 (
            .O(N__19072),
            .I(N__19062));
    InMux I__4312 (
            .O(N__19069),
            .I(N__19057));
    InMux I__4311 (
            .O(N__19068),
            .I(N__19057));
    InMux I__4310 (
            .O(N__19065),
            .I(N__19054));
    Odrv4 I__4309 (
            .O(N__19062),
            .I(\Lab_UT.dictrl.N_98_mux ));
    LocalMux I__4308 (
            .O(N__19057),
            .I(\Lab_UT.dictrl.N_98_mux ));
    LocalMux I__4307 (
            .O(N__19054),
            .I(\Lab_UT.dictrl.N_98_mux ));
    InMux I__4306 (
            .O(N__19047),
            .I(N__19041));
    InMux I__4305 (
            .O(N__19046),
            .I(N__19036));
    InMux I__4304 (
            .O(N__19045),
            .I(N__19036));
    InMux I__4303 (
            .O(N__19044),
            .I(N__19033));
    LocalMux I__4302 (
            .O(N__19041),
            .I(\Lab_UT.dictrl.N_84 ));
    LocalMux I__4301 (
            .O(N__19036),
            .I(\Lab_UT.dictrl.N_84 ));
    LocalMux I__4300 (
            .O(N__19033),
            .I(\Lab_UT.dictrl.N_84 ));
    InMux I__4299 (
            .O(N__19026),
            .I(N__19021));
    CascadeMux I__4298 (
            .O(N__19025),
            .I(N__19018));
    InMux I__4297 (
            .O(N__19024),
            .I(N__19013));
    LocalMux I__4296 (
            .O(N__19021),
            .I(N__19010));
    InMux I__4295 (
            .O(N__19018),
            .I(N__19003));
    InMux I__4294 (
            .O(N__19017),
            .I(N__19003));
    InMux I__4293 (
            .O(N__19016),
            .I(N__19003));
    LocalMux I__4292 (
            .O(N__19013),
            .I(N__19000));
    Span4Mux_h I__4291 (
            .O(N__19010),
            .I(N__18995));
    LocalMux I__4290 (
            .O(N__19003),
            .I(N__18995));
    Odrv12 I__4289 (
            .O(N__19000),
            .I(\Lab_UT.dictrl.N_89 ));
    Odrv4 I__4288 (
            .O(N__18995),
            .I(\Lab_UT.dictrl.N_89 ));
    InMux I__4287 (
            .O(N__18990),
            .I(N__18987));
    LocalMux I__4286 (
            .O(N__18987),
            .I(\Lab_UT.dictrl.m68_1 ));
    CascadeMux I__4285 (
            .O(N__18984),
            .I(\Lab_UT.dictrl.N_89_cascade_ ));
    InMux I__4284 (
            .O(N__18981),
            .I(N__18977));
    InMux I__4283 (
            .O(N__18980),
            .I(N__18974));
    LocalMux I__4282 (
            .O(N__18977),
            .I(N__18971));
    LocalMux I__4281 (
            .O(N__18974),
            .I(N__18968));
    Span4Mux_h I__4280 (
            .O(N__18971),
            .I(N__18965));
    Odrv12 I__4279 (
            .O(N__18968),
            .I(\Lab_UT.dictrl.N_99_mux ));
    Odrv4 I__4278 (
            .O(N__18965),
            .I(\Lab_UT.dictrl.N_99_mux ));
    InMux I__4277 (
            .O(N__18960),
            .I(N__18954));
    InMux I__4276 (
            .O(N__18959),
            .I(N__18954));
    LocalMux I__4275 (
            .O(N__18954),
            .I(\Lab_UT.dictrl.N_102 ));
    InMux I__4274 (
            .O(N__18951),
            .I(N__18948));
    LocalMux I__4273 (
            .O(N__18948),
            .I(N__18945));
    Span4Mux_s3_v I__4272 (
            .O(N__18945),
            .I(N__18942));
    Odrv4 I__4271 (
            .O(N__18942),
            .I(\Lab_UT.dictrl.g1_1Z0Z_0 ));
    InMux I__4270 (
            .O(N__18939),
            .I(N__18936));
    LocalMux I__4269 (
            .O(N__18936),
            .I(\Lab_UT.dictrl.g1_2Z0Z_1 ));
    InMux I__4268 (
            .O(N__18933),
            .I(N__18930));
    LocalMux I__4267 (
            .O(N__18930),
            .I(\Lab_UT.dictrl.N_102_0 ));
    CascadeMux I__4266 (
            .O(N__18927),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    CascadeMux I__4265 (
            .O(N__18924),
            .I(buart__rx_ser_clk_cascade_));
    InMux I__4264 (
            .O(N__18921),
            .I(N__18918));
    LocalMux I__4263 (
            .O(N__18918),
            .I(N__18915));
    Odrv4 I__4262 (
            .O(N__18915),
            .I(\Lab_UT.dictrl.g1_0_0_0 ));
    InMux I__4261 (
            .O(N__18912),
            .I(N__18909));
    LocalMux I__4260 (
            .O(N__18909),
            .I(N__18906));
    Span4Mux_h I__4259 (
            .O(N__18906),
            .I(N__18903));
    Odrv4 I__4258 (
            .O(N__18903),
            .I(\Lab_UT.dictrl.N_88_2 ));
    CascadeMux I__4257 (
            .O(N__18900),
            .I(N__18894));
    CascadeMux I__4256 (
            .O(N__18899),
            .I(N__18890));
    CascadeMux I__4255 (
            .O(N__18898),
            .I(N__18884));
    InMux I__4254 (
            .O(N__18897),
            .I(N__18877));
    InMux I__4253 (
            .O(N__18894),
            .I(N__18877));
    InMux I__4252 (
            .O(N__18893),
            .I(N__18874));
    InMux I__4251 (
            .O(N__18890),
            .I(N__18871));
    InMux I__4250 (
            .O(N__18889),
            .I(N__18868));
    CascadeMux I__4249 (
            .O(N__18888),
            .I(N__18865));
    InMux I__4248 (
            .O(N__18887),
            .I(N__18860));
    InMux I__4247 (
            .O(N__18884),
            .I(N__18860));
    InMux I__4246 (
            .O(N__18883),
            .I(N__18855));
    InMux I__4245 (
            .O(N__18882),
            .I(N__18855));
    LocalMux I__4244 (
            .O(N__18877),
            .I(N__18845));
    LocalMux I__4243 (
            .O(N__18874),
            .I(N__18845));
    LocalMux I__4242 (
            .O(N__18871),
            .I(N__18845));
    LocalMux I__4241 (
            .O(N__18868),
            .I(N__18845));
    InMux I__4240 (
            .O(N__18865),
            .I(N__18842));
    LocalMux I__4239 (
            .O(N__18860),
            .I(N__18839));
    LocalMux I__4238 (
            .O(N__18855),
            .I(N__18836));
    InMux I__4237 (
            .O(N__18854),
            .I(N__18833));
    Span4Mux_v I__4236 (
            .O(N__18845),
            .I(N__18826));
    LocalMux I__4235 (
            .O(N__18842),
            .I(N__18826));
    Span4Mux_s3_h I__4234 (
            .O(N__18839),
            .I(N__18826));
    Span4Mux_v I__4233 (
            .O(N__18836),
            .I(N__18821));
    LocalMux I__4232 (
            .O(N__18833),
            .I(N__18821));
    Span4Mux_h I__4231 (
            .O(N__18826),
            .I(N__18818));
    Span4Mux_v I__4230 (
            .O(N__18821),
            .I(N__18815));
    Odrv4 I__4229 (
            .O(N__18818),
            .I(bu_rx_data_i_4_3));
    Odrv4 I__4228 (
            .O(N__18815),
            .I(bu_rx_data_i_4_3));
    CascadeMux I__4227 (
            .O(N__18810),
            .I(\Lab_UT.dictrl.N_95_0_cascade_ ));
    InMux I__4226 (
            .O(N__18807),
            .I(N__18804));
    LocalMux I__4225 (
            .O(N__18804),
            .I(N__18801));
    Odrv12 I__4224 (
            .O(N__18801),
            .I(\Lab_UT.dictrl.N_103_0 ));
    CascadeMux I__4223 (
            .O(N__18798),
            .I(N__18795));
    InMux I__4222 (
            .O(N__18795),
            .I(N__18792));
    LocalMux I__4221 (
            .O(N__18792),
            .I(N__18789));
    Odrv4 I__4220 (
            .O(N__18789),
            .I(\Lab_UT.dictrl.g1_2_1_0 ));
    InMux I__4219 (
            .O(N__18786),
            .I(N__18783));
    LocalMux I__4218 (
            .O(N__18783),
            .I(N__18780));
    Odrv4 I__4217 (
            .O(N__18780),
            .I(\Lab_UT.dictrl.g1_3 ));
    InMux I__4216 (
            .O(N__18777),
            .I(N__18773));
    InMux I__4215 (
            .O(N__18776),
            .I(N__18770));
    LocalMux I__4214 (
            .O(N__18773),
            .I(N__18767));
    LocalMux I__4213 (
            .O(N__18770),
            .I(\Lab_UT.dictrl.N_88 ));
    Odrv4 I__4212 (
            .O(N__18767),
            .I(\Lab_UT.dictrl.N_88 ));
    CascadeMux I__4211 (
            .O(N__18762),
            .I(N__18759));
    InMux I__4210 (
            .O(N__18759),
            .I(N__18756));
    LocalMux I__4209 (
            .O(N__18756),
            .I(N__18753));
    Odrv12 I__4208 (
            .O(N__18753),
            .I(\Lab_UT.dictrl.N_95 ));
    InMux I__4207 (
            .O(N__18750),
            .I(N__18747));
    LocalMux I__4206 (
            .O(N__18747),
            .I(N__18744));
    Odrv4 I__4205 (
            .O(N__18744),
            .I(\Lab_UT.dictrl.N_103 ));
    InMux I__4204 (
            .O(N__18741),
            .I(N__18733));
    InMux I__4203 (
            .O(N__18740),
            .I(N__18733));
    InMux I__4202 (
            .O(N__18739),
            .I(N__18730));
    InMux I__4201 (
            .O(N__18738),
            .I(N__18726));
    LocalMux I__4200 (
            .O(N__18733),
            .I(N__18721));
    LocalMux I__4199 (
            .O(N__18730),
            .I(N__18721));
    InMux I__4198 (
            .O(N__18729),
            .I(N__18711));
    LocalMux I__4197 (
            .O(N__18726),
            .I(N__18708));
    Span4Mux_s2_v I__4196 (
            .O(N__18721),
            .I(N__18704));
    InMux I__4195 (
            .O(N__18720),
            .I(N__18701));
    InMux I__4194 (
            .O(N__18719),
            .I(N__18696));
    InMux I__4193 (
            .O(N__18718),
            .I(N__18696));
    InMux I__4192 (
            .O(N__18717),
            .I(N__18688));
    InMux I__4191 (
            .O(N__18716),
            .I(N__18688));
    InMux I__4190 (
            .O(N__18715),
            .I(N__18688));
    InMux I__4189 (
            .O(N__18714),
            .I(N__18685));
    LocalMux I__4188 (
            .O(N__18711),
            .I(N__18682));
    Span4Mux_s3_v I__4187 (
            .O(N__18708),
            .I(N__18679));
    InMux I__4186 (
            .O(N__18707),
            .I(N__18676));
    Span4Mux_v I__4185 (
            .O(N__18704),
            .I(N__18673));
    LocalMux I__4184 (
            .O(N__18701),
            .I(N__18670));
    LocalMux I__4183 (
            .O(N__18696),
            .I(N__18663));
    InMux I__4182 (
            .O(N__18695),
            .I(N__18660));
    LocalMux I__4181 (
            .O(N__18688),
            .I(N__18655));
    LocalMux I__4180 (
            .O(N__18685),
            .I(N__18655));
    Span4Mux_s3_v I__4179 (
            .O(N__18682),
            .I(N__18652));
    Span4Mux_v I__4178 (
            .O(N__18679),
            .I(N__18647));
    LocalMux I__4177 (
            .O(N__18676),
            .I(N__18647));
    Span4Mux_v I__4176 (
            .O(N__18673),
            .I(N__18644));
    Span12Mux_s10_v I__4175 (
            .O(N__18670),
            .I(N__18641));
    InMux I__4174 (
            .O(N__18669),
            .I(N__18632));
    InMux I__4173 (
            .O(N__18668),
            .I(N__18632));
    InMux I__4172 (
            .O(N__18667),
            .I(N__18632));
    InMux I__4171 (
            .O(N__18666),
            .I(N__18632));
    Span4Mux_v I__4170 (
            .O(N__18663),
            .I(N__18625));
    LocalMux I__4169 (
            .O(N__18660),
            .I(N__18625));
    Span4Mux_h I__4168 (
            .O(N__18655),
            .I(N__18625));
    Span4Mux_v I__4167 (
            .O(N__18652),
            .I(N__18620));
    Span4Mux_h I__4166 (
            .O(N__18647),
            .I(N__18620));
    Odrv4 I__4165 (
            .O(N__18644),
            .I(bu_rx_data_3));
    Odrv12 I__4164 (
            .O(N__18641),
            .I(bu_rx_data_3));
    LocalMux I__4163 (
            .O(N__18632),
            .I(bu_rx_data_3));
    Odrv4 I__4162 (
            .O(N__18625),
            .I(bu_rx_data_3));
    Odrv4 I__4161 (
            .O(N__18620),
            .I(bu_rx_data_3));
    InMux I__4160 (
            .O(N__18609),
            .I(N__18606));
    LocalMux I__4159 (
            .O(N__18606),
            .I(N__18603));
    Odrv12 I__4158 (
            .O(N__18603),
            .I(\Lab_UT.dictrl.m63_0Z0Z_1 ));
    InMux I__4157 (
            .O(N__18600),
            .I(N__18597));
    LocalMux I__4156 (
            .O(N__18597),
            .I(\Lab_UT.dictrl.N_95_0_0_1 ));
    CascadeMux I__4155 (
            .O(N__18594),
            .I(\Lab_UT.dictrl.N_99_0_cascade_ ));
    InMux I__4154 (
            .O(N__18591),
            .I(N__18588));
    LocalMux I__4153 (
            .O(N__18588),
            .I(\Lab_UT.dictrl.N_96_0_0 ));
    InMux I__4152 (
            .O(N__18585),
            .I(N__18582));
    LocalMux I__4151 (
            .O(N__18582),
            .I(N__18579));
    Odrv4 I__4150 (
            .O(N__18579),
            .I(\Lab_UT.dictrl.g2 ));
    CascadeMux I__4149 (
            .O(N__18576),
            .I(N__18573));
    InMux I__4148 (
            .O(N__18573),
            .I(N__18570));
    LocalMux I__4147 (
            .O(N__18570),
            .I(N__18567));
    Span4Mux_h I__4146 (
            .O(N__18567),
            .I(N__18564));
    Odrv4 I__4145 (
            .O(N__18564),
            .I(\Lab_UT.dictrl.g0_0_0_a3_5 ));
    InMux I__4144 (
            .O(N__18561),
            .I(N__18558));
    LocalMux I__4143 (
            .O(N__18558),
            .I(N__18555));
    Span4Mux_h I__4142 (
            .O(N__18555),
            .I(N__18552));
    Odrv4 I__4141 (
            .O(N__18552),
            .I(\Lab_UT.dictrl.N_98_mux_2 ));
    InMux I__4140 (
            .O(N__18549),
            .I(N__18545));
    InMux I__4139 (
            .O(N__18548),
            .I(N__18541));
    LocalMux I__4138 (
            .O(N__18545),
            .I(N__18538));
    CascadeMux I__4137 (
            .O(N__18544),
            .I(N__18533));
    LocalMux I__4136 (
            .O(N__18541),
            .I(N__18529));
    Span4Mux_h I__4135 (
            .O(N__18538),
            .I(N__18526));
    InMux I__4134 (
            .O(N__18537),
            .I(N__18521));
    InMux I__4133 (
            .O(N__18536),
            .I(N__18521));
    InMux I__4132 (
            .O(N__18533),
            .I(N__18516));
    InMux I__4131 (
            .O(N__18532),
            .I(N__18516));
    Span4Mux_h I__4130 (
            .O(N__18529),
            .I(N__18513));
    Span4Mux_v I__4129 (
            .O(N__18526),
            .I(N__18510));
    LocalMux I__4128 (
            .O(N__18521),
            .I(N__18505));
    LocalMux I__4127 (
            .O(N__18516),
            .I(N__18505));
    Odrv4 I__4126 (
            .O(N__18513),
            .I(bu_rx_data_i_4_5));
    Odrv4 I__4125 (
            .O(N__18510),
            .I(bu_rx_data_i_4_5));
    Odrv12 I__4124 (
            .O(N__18505),
            .I(bu_rx_data_i_4_5));
    InMux I__4123 (
            .O(N__18498),
            .I(N__18495));
    LocalMux I__4122 (
            .O(N__18495),
            .I(N__18492));
    Span4Mux_h I__4121 (
            .O(N__18492),
            .I(N__18489));
    Odrv4 I__4120 (
            .O(N__18489),
            .I(\resetGen.escKeyZ0Z_4 ));
    CascadeMux I__4119 (
            .O(N__18486),
            .I(\resetGen.escKeyZ0Z_5_cascade_ ));
    InMux I__4118 (
            .O(N__18483),
            .I(N__18468));
    InMux I__4117 (
            .O(N__18482),
            .I(N__18468));
    InMux I__4116 (
            .O(N__18481),
            .I(N__18468));
    InMux I__4115 (
            .O(N__18480),
            .I(N__18468));
    InMux I__4114 (
            .O(N__18479),
            .I(N__18468));
    LocalMux I__4113 (
            .O(N__18468),
            .I(N__18465));
    Span12Mux_s8_h I__4112 (
            .O(N__18465),
            .I(N__18462));
    Odrv12 I__4111 (
            .O(N__18462),
            .I(\resetGen.escKeyZ0 ));
    CascadeMux I__4110 (
            .O(N__18459),
            .I(\Lab_UT.dictrl.N_120_0_cascade_ ));
    InMux I__4109 (
            .O(N__18456),
            .I(N__18444));
    InMux I__4108 (
            .O(N__18455),
            .I(N__18444));
    InMux I__4107 (
            .O(N__18454),
            .I(N__18444));
    InMux I__4106 (
            .O(N__18453),
            .I(N__18444));
    LocalMux I__4105 (
            .O(N__18444),
            .I(\Lab_UT.dictrl.N_1302_0 ));
    CascadeMux I__4104 (
            .O(N__18441),
            .I(N__18437));
    CascadeMux I__4103 (
            .O(N__18440),
            .I(N__18434));
    InMux I__4102 (
            .O(N__18437),
            .I(N__18423));
    InMux I__4101 (
            .O(N__18434),
            .I(N__18423));
    InMux I__4100 (
            .O(N__18433),
            .I(N__18423));
    InMux I__4099 (
            .O(N__18432),
            .I(N__18423));
    LocalMux I__4098 (
            .O(N__18423),
            .I(\Lab_UT.dictrl.N_119_0 ));
    InMux I__4097 (
            .O(N__18420),
            .I(N__18416));
    InMux I__4096 (
            .O(N__18419),
            .I(N__18413));
    LocalMux I__4095 (
            .O(N__18416),
            .I(N__18410));
    LocalMux I__4094 (
            .O(N__18413),
            .I(N__18405));
    Span4Mux_s3_h I__4093 (
            .O(N__18410),
            .I(N__18405));
    Odrv4 I__4092 (
            .O(N__18405),
            .I(\Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0 ));
    InMux I__4091 (
            .O(N__18402),
            .I(N__18398));
    InMux I__4090 (
            .O(N__18401),
            .I(N__18395));
    LocalMux I__4089 (
            .O(N__18398),
            .I(N__18390));
    LocalMux I__4088 (
            .O(N__18395),
            .I(N__18390));
    Odrv4 I__4087 (
            .O(N__18390),
            .I(\Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0 ));
    InMux I__4086 (
            .O(N__18387),
            .I(N__18384));
    LocalMux I__4085 (
            .O(N__18384),
            .I(N__18381));
    Odrv4 I__4084 (
            .O(N__18381),
            .I(\Lab_UT.dictrl.N_120 ));
    InMux I__4083 (
            .O(N__18378),
            .I(N__18375));
    LocalMux I__4082 (
            .O(N__18375),
            .I(N__18371));
    InMux I__4081 (
            .O(N__18374),
            .I(N__18368));
    Odrv4 I__4080 (
            .O(N__18371),
            .I(\Lab_UT.dictrl.N_99 ));
    LocalMux I__4079 (
            .O(N__18368),
            .I(\Lab_UT.dictrl.N_99 ));
    InMux I__4078 (
            .O(N__18363),
            .I(N__18360));
    LocalMux I__4077 (
            .O(N__18360),
            .I(N__18356));
    InMux I__4076 (
            .O(N__18359),
            .I(N__18353));
    Odrv4 I__4075 (
            .O(N__18356),
            .I(\Lab_UT.dictrl.N_96 ));
    LocalMux I__4074 (
            .O(N__18353),
            .I(\Lab_UT.dictrl.N_96 ));
    CascadeMux I__4073 (
            .O(N__18348),
            .I(\Lab_UT.dictrl.N_99_cascade_ ));
    InMux I__4072 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__4071 (
            .O(N__18342),
            .I(N__18339));
    Odrv4 I__4070 (
            .O(N__18339),
            .I(\Lab_UT.dictrl.N_101 ));
    CascadeMux I__4069 (
            .O(N__18336),
            .I(\Lab_UT.dictrl.N_100_cascade_ ));
    InMux I__4068 (
            .O(N__18333),
            .I(N__18330));
    LocalMux I__4067 (
            .O(N__18330),
            .I(N__18327));
    Odrv4 I__4066 (
            .O(N__18327),
            .I(\Lab_UT.dictrl.next_state_0_1 ));
    CascadeMux I__4065 (
            .O(N__18324),
            .I(\Lab_UT.dictrl.N_104_cascade_ ));
    CascadeMux I__4064 (
            .O(N__18321),
            .I(\Lab_UT.dictrl.N_101_cascade_ ));
    InMux I__4063 (
            .O(N__18318),
            .I(N__18314));
    InMux I__4062 (
            .O(N__18317),
            .I(N__18311));
    LocalMux I__4061 (
            .O(N__18314),
            .I(N__18306));
    LocalMux I__4060 (
            .O(N__18311),
            .I(N__18306));
    Odrv4 I__4059 (
            .O(N__18306),
            .I(\Lab_UT.dictrl.N_5_0 ));
    CascadeMux I__4058 (
            .O(N__18303),
            .I(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_ ));
    InMux I__4057 (
            .O(N__18300),
            .I(N__18297));
    LocalMux I__4056 (
            .O(N__18297),
            .I(N__18294));
    Span4Mux_h I__4055 (
            .O(N__18294),
            .I(N__18291));
    Odrv4 I__4054 (
            .O(N__18291),
            .I(\Lab_UT.dictrl.state_fast_3 ));
    InMux I__4053 (
            .O(N__18288),
            .I(N__18283));
    InMux I__4052 (
            .O(N__18287),
            .I(N__18276));
    InMux I__4051 (
            .O(N__18286),
            .I(N__18276));
    LocalMux I__4050 (
            .O(N__18283),
            .I(N__18273));
    InMux I__4049 (
            .O(N__18282),
            .I(N__18268));
    InMux I__4048 (
            .O(N__18281),
            .I(N__18268));
    LocalMux I__4047 (
            .O(N__18276),
            .I(N__18265));
    Span4Mux_h I__4046 (
            .O(N__18273),
            .I(N__18262));
    LocalMux I__4045 (
            .O(N__18268),
            .I(N__18257));
    Span4Mux_h I__4044 (
            .O(N__18265),
            .I(N__18257));
    Odrv4 I__4043 (
            .O(N__18262),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    Odrv4 I__4042 (
            .O(N__18257),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    CEMux I__4041 (
            .O(N__18252),
            .I(N__18237));
    CEMux I__4040 (
            .O(N__18251),
            .I(N__18237));
    CEMux I__4039 (
            .O(N__18250),
            .I(N__18237));
    CEMux I__4038 (
            .O(N__18249),
            .I(N__18237));
    CEMux I__4037 (
            .O(N__18248),
            .I(N__18237));
    GlobalMux I__4036 (
            .O(N__18237),
            .I(N__18234));
    gio2CtrlBuf I__4035 (
            .O(N__18234),
            .I(bu_rx_data_rdy_0_g));
    InMux I__4034 (
            .O(N__18231),
            .I(N__18228));
    LocalMux I__4033 (
            .O(N__18228),
            .I(N__18220));
    InMux I__4032 (
            .O(N__18227),
            .I(N__18217));
    InMux I__4031 (
            .O(N__18226),
            .I(N__18211));
    InMux I__4030 (
            .O(N__18225),
            .I(N__18208));
    CascadeMux I__4029 (
            .O(N__18224),
            .I(N__18205));
    CascadeMux I__4028 (
            .O(N__18223),
            .I(N__18202));
    Span4Mux_s1_v I__4027 (
            .O(N__18220),
            .I(N__18195));
    LocalMux I__4026 (
            .O(N__18217),
            .I(N__18195));
    InMux I__4025 (
            .O(N__18216),
            .I(N__18192));
    InMux I__4024 (
            .O(N__18215),
            .I(N__18188));
    InMux I__4023 (
            .O(N__18214),
            .I(N__18185));
    LocalMux I__4022 (
            .O(N__18211),
            .I(N__18180));
    LocalMux I__4021 (
            .O(N__18208),
            .I(N__18180));
    InMux I__4020 (
            .O(N__18205),
            .I(N__18177));
    InMux I__4019 (
            .O(N__18202),
            .I(N__18174));
    InMux I__4018 (
            .O(N__18201),
            .I(N__18169));
    InMux I__4017 (
            .O(N__18200),
            .I(N__18169));
    Span4Mux_v I__4016 (
            .O(N__18195),
            .I(N__18164));
    LocalMux I__4015 (
            .O(N__18192),
            .I(N__18164));
    InMux I__4014 (
            .O(N__18191),
            .I(N__18161));
    LocalMux I__4013 (
            .O(N__18188),
            .I(N__18158));
    LocalMux I__4012 (
            .O(N__18185),
            .I(N__18155));
    Span4Mux_v I__4011 (
            .O(N__18180),
            .I(N__18147));
    LocalMux I__4010 (
            .O(N__18177),
            .I(N__18147));
    LocalMux I__4009 (
            .O(N__18174),
            .I(N__18147));
    LocalMux I__4008 (
            .O(N__18169),
            .I(N__18144));
    Span4Mux_v I__4007 (
            .O(N__18164),
            .I(N__18141));
    LocalMux I__4006 (
            .O(N__18161),
            .I(N__18138));
    Span12Mux_s11_v I__4005 (
            .O(N__18158),
            .I(N__18132));
    Span12Mux_s6_v I__4004 (
            .O(N__18155),
            .I(N__18129));
    InMux I__4003 (
            .O(N__18154),
            .I(N__18126));
    Span4Mux_v I__4002 (
            .O(N__18147),
            .I(N__18123));
    Span4Mux_v I__4001 (
            .O(N__18144),
            .I(N__18116));
    Span4Mux_h I__4000 (
            .O(N__18141),
            .I(N__18116));
    Span4Mux_h I__3999 (
            .O(N__18138),
            .I(N__18116));
    InMux I__3998 (
            .O(N__18137),
            .I(N__18113));
    InMux I__3997 (
            .O(N__18136),
            .I(N__18108));
    InMux I__3996 (
            .O(N__18135),
            .I(N__18108));
    Odrv12 I__3995 (
            .O(N__18132),
            .I(bu_rx_data_0));
    Odrv12 I__3994 (
            .O(N__18129),
            .I(bu_rx_data_0));
    LocalMux I__3993 (
            .O(N__18126),
            .I(bu_rx_data_0));
    Odrv4 I__3992 (
            .O(N__18123),
            .I(bu_rx_data_0));
    Odrv4 I__3991 (
            .O(N__18116),
            .I(bu_rx_data_0));
    LocalMux I__3990 (
            .O(N__18113),
            .I(bu_rx_data_0));
    LocalMux I__3989 (
            .O(N__18108),
            .I(bu_rx_data_0));
    CascadeMux I__3988 (
            .O(N__18093),
            .I(N__18090));
    InMux I__3987 (
            .O(N__18090),
            .I(N__18087));
    LocalMux I__3986 (
            .O(N__18087),
            .I(N__18084));
    Odrv12 I__3985 (
            .O(N__18084),
            .I(\Lab_UT.dictrl.g0_9Z0Z_1 ));
    InMux I__3984 (
            .O(N__18081),
            .I(N__18078));
    LocalMux I__3983 (
            .O(N__18078),
            .I(N__18073));
    InMux I__3982 (
            .O(N__18077),
            .I(N__18068));
    InMux I__3981 (
            .O(N__18076),
            .I(N__18068));
    Span4Mux_h I__3980 (
            .O(N__18073),
            .I(N__18064));
    LocalMux I__3979 (
            .O(N__18068),
            .I(N__18061));
    InMux I__3978 (
            .O(N__18067),
            .I(N__18058));
    Odrv4 I__3977 (
            .O(N__18064),
            .I(\Lab_UT.dictrl.m25Z0Z_4 ));
    Odrv4 I__3976 (
            .O(N__18061),
            .I(\Lab_UT.dictrl.m25Z0Z_4 ));
    LocalMux I__3975 (
            .O(N__18058),
            .I(\Lab_UT.dictrl.m25Z0Z_4 ));
    CascadeMux I__3974 (
            .O(N__18051),
            .I(\Lab_UT.dictrl.N_116_mux_1_cascade_ ));
    InMux I__3973 (
            .O(N__18048),
            .I(N__18045));
    LocalMux I__3972 (
            .O(N__18045),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__3971 (
            .O(N__18042),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__3970 (
            .O(N__18039),
            .I(N__18036));
    LocalMux I__3969 (
            .O(N__18036),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__3968 (
            .O(N__18033),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__3967 (
            .O(N__18030),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__3966 (
            .O(N__18027),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__3965 (
            .O(N__18024),
            .I(N__18021));
    InMux I__3964 (
            .O(N__18021),
            .I(N__18017));
    InMux I__3963 (
            .O(N__18020),
            .I(N__18014));
    LocalMux I__3962 (
            .O(N__18017),
            .I(N__18011));
    LocalMux I__3961 (
            .O(N__18014),
            .I(N__18006));
    Span4Mux_h I__3960 (
            .O(N__18011),
            .I(N__18006));
    Odrv4 I__3959 (
            .O(N__18006),
            .I(\Lab_UT.dictrl.state_i_4_0 ));
    CascadeMux I__3958 (
            .O(N__18003),
            .I(\Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_ ));
    InMux I__3957 (
            .O(N__18000),
            .I(N__17997));
    LocalMux I__3956 (
            .O(N__17997),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    CascadeMux I__3955 (
            .O(N__17994),
            .I(N__17990));
    InMux I__3954 (
            .O(N__17993),
            .I(N__17985));
    InMux I__3953 (
            .O(N__17990),
            .I(N__17978));
    InMux I__3952 (
            .O(N__17989),
            .I(N__17978));
    InMux I__3951 (
            .O(N__17988),
            .I(N__17978));
    LocalMux I__3950 (
            .O(N__17985),
            .I(\Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2 ));
    LocalMux I__3949 (
            .O(N__17978),
            .I(\Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2 ));
    InMux I__3948 (
            .O(N__17973),
            .I(N__17970));
    LocalMux I__3947 (
            .O(N__17970),
            .I(N__17967));
    Span4Mux_v I__3946 (
            .O(N__17967),
            .I(N__17964));
    Span4Mux_v I__3945 (
            .O(N__17964),
            .I(N__17961));
    Odrv4 I__3944 (
            .O(N__17961),
            .I(\Lab_UT.dictrl.dicLdStens_1 ));
    CascadeMux I__3943 (
            .O(N__17958),
            .I(N__17954));
    InMux I__3942 (
            .O(N__17957),
            .I(N__17949));
    InMux I__3941 (
            .O(N__17954),
            .I(N__17949));
    LocalMux I__3940 (
            .O(N__17949),
            .I(N__17944));
    InMux I__3939 (
            .O(N__17948),
            .I(N__17941));
    InMux I__3938 (
            .O(N__17947),
            .I(N__17938));
    Odrv4 I__3937 (
            .O(N__17944),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    LocalMux I__3936 (
            .O(N__17941),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    LocalMux I__3935 (
            .O(N__17938),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    CascadeMux I__3934 (
            .O(N__17931),
            .I(\Lab_UT.didp.countrce2.q_5_1_cascade_ ));
    InMux I__3933 (
            .O(N__17928),
            .I(N__17922));
    InMux I__3932 (
            .O(N__17927),
            .I(N__17915));
    InMux I__3931 (
            .O(N__17926),
            .I(N__17915));
    InMux I__3930 (
            .O(N__17925),
            .I(N__17912));
    LocalMux I__3929 (
            .O(N__17922),
            .I(N__17909));
    InMux I__3928 (
            .O(N__17921),
            .I(N__17904));
    InMux I__3927 (
            .O(N__17920),
            .I(N__17904));
    LocalMux I__3926 (
            .O(N__17915),
            .I(\Lab_UT.didp.di_Stens_1 ));
    LocalMux I__3925 (
            .O(N__17912),
            .I(\Lab_UT.didp.di_Stens_1 ));
    Odrv12 I__3924 (
            .O(N__17909),
            .I(\Lab_UT.didp.di_Stens_1 ));
    LocalMux I__3923 (
            .O(N__17904),
            .I(\Lab_UT.didp.di_Stens_1 ));
    InMux I__3922 (
            .O(N__17895),
            .I(N__17891));
    CascadeMux I__3921 (
            .O(N__17894),
            .I(N__17887));
    LocalMux I__3920 (
            .O(N__17891),
            .I(N__17883));
    InMux I__3919 (
            .O(N__17890),
            .I(N__17876));
    InMux I__3918 (
            .O(N__17887),
            .I(N__17876));
    InMux I__3917 (
            .O(N__17886),
            .I(N__17876));
    Odrv4 I__3916 (
            .O(N__17883),
            .I(\Lab_UT.LdStens ));
    LocalMux I__3915 (
            .O(N__17876),
            .I(\Lab_UT.LdStens ));
    InMux I__3914 (
            .O(N__17871),
            .I(N__17868));
    LocalMux I__3913 (
            .O(N__17868),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__3912 (
            .O(N__17865),
            .I(N__17862));
    LocalMux I__3911 (
            .O(N__17862),
            .I(\Lab_UT.LdStens_i_4 ));
    InMux I__3910 (
            .O(N__17859),
            .I(N__17853));
    InMux I__3909 (
            .O(N__17858),
            .I(N__17853));
    LocalMux I__3908 (
            .O(N__17853),
            .I(N__17848));
    InMux I__3907 (
            .O(N__17852),
            .I(N__17845));
    InMux I__3906 (
            .O(N__17851),
            .I(N__17842));
    Odrv4 I__3905 (
            .O(N__17848),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    LocalMux I__3904 (
            .O(N__17845),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    LocalMux I__3903 (
            .O(N__17842),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    CascadeMux I__3902 (
            .O(N__17835),
            .I(N__17830));
    InMux I__3901 (
            .O(N__17834),
            .I(N__17825));
    InMux I__3900 (
            .O(N__17833),
            .I(N__17825));
    InMux I__3899 (
            .O(N__17830),
            .I(N__17822));
    LocalMux I__3898 (
            .O(N__17825),
            .I(N__17819));
    LocalMux I__3897 (
            .O(N__17822),
            .I(N__17816));
    Span4Mux_s2_v I__3896 (
            .O(N__17819),
            .I(N__17812));
    Span4Mux_s2_v I__3895 (
            .O(N__17816),
            .I(N__17809));
    InMux I__3894 (
            .O(N__17815),
            .I(N__17806));
    Odrv4 I__3893 (
            .O(N__17812),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__3892 (
            .O(N__17809),
            .I(\Lab_UT.LdSones ));
    LocalMux I__3891 (
            .O(N__17806),
            .I(\Lab_UT.LdSones ));
    InMux I__3890 (
            .O(N__17799),
            .I(N__17796));
    LocalMux I__3889 (
            .O(N__17796),
            .I(N__17787));
    InMux I__3888 (
            .O(N__17795),
            .I(N__17782));
    InMux I__3887 (
            .O(N__17794),
            .I(N__17782));
    InMux I__3886 (
            .O(N__17793),
            .I(N__17779));
    InMux I__3885 (
            .O(N__17792),
            .I(N__17772));
    InMux I__3884 (
            .O(N__17791),
            .I(N__17772));
    InMux I__3883 (
            .O(N__17790),
            .I(N__17772));
    Span4Mux_h I__3882 (
            .O(N__17787),
            .I(N__17767));
    LocalMux I__3881 (
            .O(N__17782),
            .I(N__17767));
    LocalMux I__3880 (
            .O(N__17779),
            .I(\Lab_UT.didp.di_Sones_0 ));
    LocalMux I__3879 (
            .O(N__17772),
            .I(\Lab_UT.didp.di_Sones_0 ));
    Odrv4 I__3878 (
            .O(N__17767),
            .I(\Lab_UT.didp.di_Sones_0 ));
    InMux I__3877 (
            .O(N__17760),
            .I(N__17757));
    LocalMux I__3876 (
            .O(N__17757),
            .I(N__17754));
    Span4Mux_s2_v I__3875 (
            .O(N__17754),
            .I(N__17751));
    Odrv4 I__3874 (
            .O(N__17751),
            .I(\Lab_UT.didp.countrce1.q_5_0 ));
    CascadeMux I__3873 (
            .O(N__17748),
            .I(N__17742));
    CascadeMux I__3872 (
            .O(N__17747),
            .I(N__17739));
    InMux I__3871 (
            .O(N__17746),
            .I(N__17732));
    InMux I__3870 (
            .O(N__17745),
            .I(N__17732));
    InMux I__3869 (
            .O(N__17742),
            .I(N__17732));
    InMux I__3868 (
            .O(N__17739),
            .I(N__17729));
    LocalMux I__3867 (
            .O(N__17732),
            .I(N__17726));
    LocalMux I__3866 (
            .O(N__17729),
            .I(N__17723));
    Span4Mux_s3_v I__3865 (
            .O(N__17726),
            .I(N__17717));
    Span4Mux_s3_h I__3864 (
            .O(N__17723),
            .I(N__17717));
    InMux I__3863 (
            .O(N__17722),
            .I(N__17714));
    Odrv4 I__3862 (
            .O(N__17717),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    LocalMux I__3861 (
            .O(N__17714),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2 ));
    InMux I__3860 (
            .O(N__17709),
            .I(N__17706));
    LocalMux I__3859 (
            .O(N__17706),
            .I(N__17703));
    Span4Mux_s3_v I__3858 (
            .O(N__17703),
            .I(N__17700));
    Odrv4 I__3857 (
            .O(N__17700),
            .I(\Lab_UT.LdSones_i_4 ));
    CascadeMux I__3856 (
            .O(N__17697),
            .I(\Lab_UT.didp.countrce2.un13_qPone_cascade_ ));
    CascadeMux I__3855 (
            .O(N__17694),
            .I(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ));
    CascadeMux I__3854 (
            .O(N__17691),
            .I(\Lab_UT.didp.countrce2.q_5_3_cascade_ ));
    CascadeMux I__3853 (
            .O(N__17688),
            .I(N__17684));
    CascadeMux I__3852 (
            .O(N__17687),
            .I(N__17681));
    InMux I__3851 (
            .O(N__17684),
            .I(N__17678));
    InMux I__3850 (
            .O(N__17681),
            .I(N__17672));
    LocalMux I__3849 (
            .O(N__17678),
            .I(N__17669));
    InMux I__3848 (
            .O(N__17677),
            .I(N__17666));
    InMux I__3847 (
            .O(N__17676),
            .I(N__17663));
    InMux I__3846 (
            .O(N__17675),
            .I(N__17660));
    LocalMux I__3845 (
            .O(N__17672),
            .I(N__17657));
    Span4Mux_h I__3844 (
            .O(N__17669),
            .I(N__17654));
    LocalMux I__3843 (
            .O(N__17666),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3842 (
            .O(N__17663),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3841 (
            .O(N__17660),
            .I(\Lab_UT.didp.di_Stens_3 ));
    Odrv12 I__3840 (
            .O(N__17657),
            .I(\Lab_UT.didp.di_Stens_3 ));
    Odrv4 I__3839 (
            .O(N__17654),
            .I(\Lab_UT.didp.di_Stens_3 ));
    InMux I__3838 (
            .O(N__17643),
            .I(N__17640));
    LocalMux I__3837 (
            .O(N__17640),
            .I(\Lab_UT.didp.countrce2.q_5_0 ));
    InMux I__3836 (
            .O(N__17637),
            .I(N__17630));
    InMux I__3835 (
            .O(N__17636),
            .I(N__17627));
    InMux I__3834 (
            .O(N__17635),
            .I(N__17624));
    InMux I__3833 (
            .O(N__17634),
            .I(N__17621));
    InMux I__3832 (
            .O(N__17633),
            .I(N__17617));
    LocalMux I__3831 (
            .O(N__17630),
            .I(N__17610));
    LocalMux I__3830 (
            .O(N__17627),
            .I(N__17610));
    LocalMux I__3829 (
            .O(N__17624),
            .I(N__17607));
    LocalMux I__3828 (
            .O(N__17621),
            .I(N__17604));
    InMux I__3827 (
            .O(N__17620),
            .I(N__17601));
    LocalMux I__3826 (
            .O(N__17617),
            .I(N__17597));
    InMux I__3825 (
            .O(N__17616),
            .I(N__17591));
    InMux I__3824 (
            .O(N__17615),
            .I(N__17591));
    Span4Mux_s2_v I__3823 (
            .O(N__17610),
            .I(N__17588));
    Span4Mux_h I__3822 (
            .O(N__17607),
            .I(N__17581));
    Span4Mux_s2_v I__3821 (
            .O(N__17604),
            .I(N__17581));
    LocalMux I__3820 (
            .O(N__17601),
            .I(N__17581));
    InMux I__3819 (
            .O(N__17600),
            .I(N__17578));
    Span4Mux_h I__3818 (
            .O(N__17597),
            .I(N__17575));
    InMux I__3817 (
            .O(N__17596),
            .I(N__17572));
    LocalMux I__3816 (
            .O(N__17591),
            .I(N__17567));
    Span4Mux_v I__3815 (
            .O(N__17588),
            .I(N__17567));
    Span4Mux_v I__3814 (
            .O(N__17581),
            .I(N__17558));
    LocalMux I__3813 (
            .O(N__17578),
            .I(N__17558));
    Span4Mux_v I__3812 (
            .O(N__17575),
            .I(N__17555));
    LocalMux I__3811 (
            .O(N__17572),
            .I(N__17552));
    Span4Mux_h I__3810 (
            .O(N__17567),
            .I(N__17549));
    InMux I__3809 (
            .O(N__17566),
            .I(N__17540));
    InMux I__3808 (
            .O(N__17565),
            .I(N__17540));
    InMux I__3807 (
            .O(N__17564),
            .I(N__17540));
    InMux I__3806 (
            .O(N__17563),
            .I(N__17540));
    Span4Mux_v I__3805 (
            .O(N__17558),
            .I(N__17537));
    Odrv4 I__3804 (
            .O(N__17555),
            .I(bu_rx_data_2));
    Odrv4 I__3803 (
            .O(N__17552),
            .I(bu_rx_data_2));
    Odrv4 I__3802 (
            .O(N__17549),
            .I(bu_rx_data_2));
    LocalMux I__3801 (
            .O(N__17540),
            .I(bu_rx_data_2));
    Odrv4 I__3800 (
            .O(N__17537),
            .I(bu_rx_data_2));
    InMux I__3799 (
            .O(N__17526),
            .I(N__17523));
    LocalMux I__3798 (
            .O(N__17523),
            .I(\Lab_UT.didp.countrce2.un13_qPone ));
    CascadeMux I__3797 (
            .O(N__17520),
            .I(\Lab_UT.didp.countrce2.q_5_2_cascade_ ));
    CascadeMux I__3796 (
            .O(N__17517),
            .I(N__17511));
    CascadeMux I__3795 (
            .O(N__17516),
            .I(N__17507));
    InMux I__3794 (
            .O(N__17515),
            .I(N__17504));
    InMux I__3793 (
            .O(N__17514),
            .I(N__17500));
    InMux I__3792 (
            .O(N__17511),
            .I(N__17497));
    InMux I__3791 (
            .O(N__17510),
            .I(N__17494));
    InMux I__3790 (
            .O(N__17507),
            .I(N__17491));
    LocalMux I__3789 (
            .O(N__17504),
            .I(N__17488));
    InMux I__3788 (
            .O(N__17503),
            .I(N__17485));
    LocalMux I__3787 (
            .O(N__17500),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__3786 (
            .O(N__17497),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__3785 (
            .O(N__17494),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__3784 (
            .O(N__17491),
            .I(\Lab_UT.didp.di_Stens_2 ));
    Odrv12 I__3783 (
            .O(N__17488),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__3782 (
            .O(N__17485),
            .I(\Lab_UT.didp.di_Stens_2 ));
    InMux I__3781 (
            .O(N__17472),
            .I(N__17467));
    InMux I__3780 (
            .O(N__17471),
            .I(N__17464));
    InMux I__3779 (
            .O(N__17470),
            .I(N__17457));
    LocalMux I__3778 (
            .O(N__17467),
            .I(N__17452));
    LocalMux I__3777 (
            .O(N__17464),
            .I(N__17452));
    InMux I__3776 (
            .O(N__17463),
            .I(N__17447));
    InMux I__3775 (
            .O(N__17462),
            .I(N__17447));
    InMux I__3774 (
            .O(N__17461),
            .I(N__17442));
    InMux I__3773 (
            .O(N__17460),
            .I(N__17442));
    LocalMux I__3772 (
            .O(N__17457),
            .I(N__17437));
    Span4Mux_h I__3771 (
            .O(N__17452),
            .I(N__17437));
    LocalMux I__3770 (
            .O(N__17447),
            .I(\Lab_UT.didp.di_Stens_0 ));
    LocalMux I__3769 (
            .O(N__17442),
            .I(\Lab_UT.didp.di_Stens_0 ));
    Odrv4 I__3768 (
            .O(N__17437),
            .I(\Lab_UT.didp.di_Stens_0 ));
    InMux I__3767 (
            .O(N__17430),
            .I(N__17424));
    InMux I__3766 (
            .O(N__17429),
            .I(N__17421));
    CascadeMux I__3765 (
            .O(N__17428),
            .I(N__17417));
    CascadeMux I__3764 (
            .O(N__17427),
            .I(N__17414));
    LocalMux I__3763 (
            .O(N__17424),
            .I(N__17409));
    LocalMux I__3762 (
            .O(N__17421),
            .I(N__17409));
    InMux I__3761 (
            .O(N__17420),
            .I(N__17402));
    InMux I__3760 (
            .O(N__17417),
            .I(N__17402));
    InMux I__3759 (
            .O(N__17414),
            .I(N__17402));
    Span4Mux_v I__3758 (
            .O(N__17409),
            .I(N__17397));
    LocalMux I__3757 (
            .O(N__17402),
            .I(N__17397));
    Span4Mux_h I__3756 (
            .O(N__17397),
            .I(N__17394));
    Odrv4 I__3755 (
            .O(N__17394),
            .I(buart__rx_shifter_0_fast_3));
    InMux I__3754 (
            .O(N__17391),
            .I(N__17388));
    LocalMux I__3753 (
            .O(N__17388),
            .I(N__17384));
    InMux I__3752 (
            .O(N__17387),
            .I(N__17381));
    Span4Mux_v I__3751 (
            .O(N__17384),
            .I(N__17372));
    LocalMux I__3750 (
            .O(N__17381),
            .I(N__17369));
    InMux I__3749 (
            .O(N__17380),
            .I(N__17362));
    InMux I__3748 (
            .O(N__17379),
            .I(N__17362));
    InMux I__3747 (
            .O(N__17378),
            .I(N__17362));
    InMux I__3746 (
            .O(N__17377),
            .I(N__17355));
    InMux I__3745 (
            .O(N__17376),
            .I(N__17355));
    InMux I__3744 (
            .O(N__17375),
            .I(N__17355));
    Odrv4 I__3743 (
            .O(N__17372),
            .I(bu_rx_data_5_rep1));
    Odrv4 I__3742 (
            .O(N__17369),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3741 (
            .O(N__17362),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3740 (
            .O(N__17355),
            .I(bu_rx_data_5_rep1));
    InMux I__3739 (
            .O(N__17346),
            .I(N__17343));
    LocalMux I__3738 (
            .O(N__17343),
            .I(N__17339));
    InMux I__3737 (
            .O(N__17342),
            .I(N__17332));
    Span4Mux_v I__3736 (
            .O(N__17339),
            .I(N__17329));
    InMux I__3735 (
            .O(N__17338),
            .I(N__17320));
    InMux I__3734 (
            .O(N__17337),
            .I(N__17320));
    InMux I__3733 (
            .O(N__17336),
            .I(N__17320));
    InMux I__3732 (
            .O(N__17335),
            .I(N__17320));
    LocalMux I__3731 (
            .O(N__17332),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__3730 (
            .O(N__17329),
            .I(bu_rx_data_4_rep1));
    LocalMux I__3729 (
            .O(N__17320),
            .I(bu_rx_data_4_rep1));
    InMux I__3728 (
            .O(N__17313),
            .I(N__17308));
    CascadeMux I__3727 (
            .O(N__17312),
            .I(N__17303));
    InMux I__3726 (
            .O(N__17311),
            .I(N__17300));
    LocalMux I__3725 (
            .O(N__17308),
            .I(N__17297));
    InMux I__3724 (
            .O(N__17307),
            .I(N__17292));
    InMux I__3723 (
            .O(N__17306),
            .I(N__17292));
    InMux I__3722 (
            .O(N__17303),
            .I(N__17289));
    LocalMux I__3721 (
            .O(N__17300),
            .I(N__17286));
    Odrv4 I__3720 (
            .O(N__17297),
            .I(bu_rx_data_fast_5));
    LocalMux I__3719 (
            .O(N__17292),
            .I(bu_rx_data_fast_5));
    LocalMux I__3718 (
            .O(N__17289),
            .I(bu_rx_data_fast_5));
    Odrv4 I__3717 (
            .O(N__17286),
            .I(bu_rx_data_fast_5));
    CascadeMux I__3716 (
            .O(N__17277),
            .I(N__17272));
    CascadeMux I__3715 (
            .O(N__17276),
            .I(N__17266));
    InMux I__3714 (
            .O(N__17275),
            .I(N__17263));
    InMux I__3713 (
            .O(N__17272),
            .I(N__17256));
    InMux I__3712 (
            .O(N__17271),
            .I(N__17256));
    InMux I__3711 (
            .O(N__17270),
            .I(N__17256));
    InMux I__3710 (
            .O(N__17269),
            .I(N__17251));
    InMux I__3709 (
            .O(N__17266),
            .I(N__17251));
    LocalMux I__3708 (
            .O(N__17263),
            .I(bu_rx_data_i_4_7_rep1));
    LocalMux I__3707 (
            .O(N__17256),
            .I(bu_rx_data_i_4_7_rep1));
    LocalMux I__3706 (
            .O(N__17251),
            .I(bu_rx_data_i_4_7_rep1));
    CascadeMux I__3705 (
            .O(N__17244),
            .I(N__17241));
    InMux I__3704 (
            .O(N__17241),
            .I(N__17238));
    LocalMux I__3703 (
            .O(N__17238),
            .I(\Lab_UT.dictrl.g0_28_1Z0Z_0 ));
    InMux I__3702 (
            .O(N__17235),
            .I(N__17229));
    InMux I__3701 (
            .O(N__17234),
            .I(N__17226));
    InMux I__3700 (
            .O(N__17233),
            .I(N__17223));
    InMux I__3699 (
            .O(N__17232),
            .I(N__17220));
    LocalMux I__3698 (
            .O(N__17229),
            .I(N__17217));
    LocalMux I__3697 (
            .O(N__17226),
            .I(N__17210));
    LocalMux I__3696 (
            .O(N__17223),
            .I(N__17210));
    LocalMux I__3695 (
            .O(N__17220),
            .I(N__17210));
    Span4Mux_h I__3694 (
            .O(N__17217),
            .I(N__17207));
    Odrv4 I__3693 (
            .O(N__17210),
            .I(bu_rx_data_fast_6));
    Odrv4 I__3692 (
            .O(N__17207),
            .I(bu_rx_data_fast_6));
    InMux I__3691 (
            .O(N__17202),
            .I(N__17199));
    LocalMux I__3690 (
            .O(N__17199),
            .I(\Lab_UT.dictrl.m31_xZ0Z0 ));
    InMux I__3689 (
            .O(N__17196),
            .I(N__17185));
    InMux I__3688 (
            .O(N__17195),
            .I(N__17185));
    InMux I__3687 (
            .O(N__17194),
            .I(N__17185));
    InMux I__3686 (
            .O(N__17193),
            .I(N__17180));
    InMux I__3685 (
            .O(N__17192),
            .I(N__17180));
    LocalMux I__3684 (
            .O(N__17185),
            .I(N__17177));
    LocalMux I__3683 (
            .O(N__17180),
            .I(N__17171));
    Span4Mux_h I__3682 (
            .O(N__17177),
            .I(N__17171));
    InMux I__3681 (
            .O(N__17176),
            .I(N__17168));
    Odrv4 I__3680 (
            .O(N__17171),
            .I(bu_rx_data_6_rep1));
    LocalMux I__3679 (
            .O(N__17168),
            .I(bu_rx_data_6_rep1));
    InMux I__3678 (
            .O(N__17163),
            .I(N__17160));
    LocalMux I__3677 (
            .O(N__17160),
            .I(N__17157));
    Odrv4 I__3676 (
            .O(N__17157),
            .I(\Lab_UT.dictrl.g0_43_xZ0 ));
    CascadeMux I__3675 (
            .O(N__17154),
            .I(\Lab_UT.dictrl.N_84_cascade_ ));
    InMux I__3674 (
            .O(N__17151),
            .I(N__17148));
    LocalMux I__3673 (
            .O(N__17148),
            .I(N__17144));
    InMux I__3672 (
            .O(N__17147),
            .I(N__17141));
    Span4Mux_h I__3671 (
            .O(N__17144),
            .I(N__17138));
    LocalMux I__3670 (
            .O(N__17141),
            .I(N__17135));
    Odrv4 I__3669 (
            .O(N__17138),
            .I(\Lab_UT.dictrl.alarmstate8_2 ));
    Odrv4 I__3668 (
            .O(N__17135),
            .I(\Lab_UT.dictrl.alarmstate8_2 ));
    CascadeMux I__3667 (
            .O(N__17130),
            .I(N__17127));
    InMux I__3666 (
            .O(N__17127),
            .I(N__17124));
    LocalMux I__3665 (
            .O(N__17124),
            .I(\Lab_UT.dictrl.g1_0_0_0_0 ));
    InMux I__3664 (
            .O(N__17121),
            .I(N__17118));
    LocalMux I__3663 (
            .O(N__17118),
            .I(N__17115));
    Odrv4 I__3662 (
            .O(N__17115),
            .I(\Lab_UT.dictrl.g0_4_a4Z0Z_5 ));
    InMux I__3661 (
            .O(N__17112),
            .I(N__17108));
    CascadeMux I__3660 (
            .O(N__17111),
            .I(N__17105));
    LocalMux I__3659 (
            .O(N__17108),
            .I(N__17101));
    InMux I__3658 (
            .O(N__17105),
            .I(N__17096));
    InMux I__3657 (
            .O(N__17104),
            .I(N__17096));
    Sp12to4 I__3656 (
            .O(N__17101),
            .I(N__17091));
    LocalMux I__3655 (
            .O(N__17096),
            .I(N__17091));
    Odrv12 I__3654 (
            .O(N__17091),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    CascadeMux I__3653 (
            .O(N__17088),
            .I(N__17083));
    CascadeMux I__3652 (
            .O(N__17087),
            .I(N__17079));
    InMux I__3651 (
            .O(N__17086),
            .I(N__17075));
    InMux I__3650 (
            .O(N__17083),
            .I(N__17068));
    InMux I__3649 (
            .O(N__17082),
            .I(N__17068));
    InMux I__3648 (
            .O(N__17079),
            .I(N__17068));
    CascadeMux I__3647 (
            .O(N__17078),
            .I(N__17065));
    LocalMux I__3646 (
            .O(N__17075),
            .I(N__17060));
    LocalMux I__3645 (
            .O(N__17068),
            .I(N__17060));
    InMux I__3644 (
            .O(N__17065),
            .I(N__17057));
    Span4Mux_h I__3643 (
            .O(N__17060),
            .I(N__17054));
    LocalMux I__3642 (
            .O(N__17057),
            .I(bu_rx_data_i_4_0));
    Odrv4 I__3641 (
            .O(N__17054),
            .I(bu_rx_data_i_4_0));
    InMux I__3640 (
            .O(N__17049),
            .I(N__17046));
    LocalMux I__3639 (
            .O(N__17046),
            .I(\Lab_UT.dictrl.g1_5 ));
    InMux I__3638 (
            .O(N__17043),
            .I(N__17040));
    LocalMux I__3637 (
            .O(N__17040),
            .I(\Lab_UT.dictrl.g0_5_4 ));
    CascadeMux I__3636 (
            .O(N__17037),
            .I(N__17031));
    CascadeMux I__3635 (
            .O(N__17036),
            .I(N__17027));
    CascadeMux I__3634 (
            .O(N__17035),
            .I(N__17022));
    CascadeMux I__3633 (
            .O(N__17034),
            .I(N__17018));
    InMux I__3632 (
            .O(N__17031),
            .I(N__17007));
    InMux I__3631 (
            .O(N__17030),
            .I(N__17007));
    InMux I__3630 (
            .O(N__17027),
            .I(N__17007));
    InMux I__3629 (
            .O(N__17026),
            .I(N__17007));
    InMux I__3628 (
            .O(N__17025),
            .I(N__17007));
    InMux I__3627 (
            .O(N__17022),
            .I(N__16999));
    InMux I__3626 (
            .O(N__17021),
            .I(N__16999));
    InMux I__3625 (
            .O(N__17018),
            .I(N__16999));
    LocalMux I__3624 (
            .O(N__17007),
            .I(N__16995));
    InMux I__3623 (
            .O(N__17006),
            .I(N__16990));
    LocalMux I__3622 (
            .O(N__16999),
            .I(N__16987));
    InMux I__3621 (
            .O(N__16998),
            .I(N__16984));
    Span4Mux_v I__3620 (
            .O(N__16995),
            .I(N__16981));
    InMux I__3619 (
            .O(N__16994),
            .I(N__16978));
    InMux I__3618 (
            .O(N__16993),
            .I(N__16975));
    LocalMux I__3617 (
            .O(N__16990),
            .I(N__16972));
    Span4Mux_v I__3616 (
            .O(N__16987),
            .I(N__16967));
    LocalMux I__3615 (
            .O(N__16984),
            .I(N__16967));
    Odrv4 I__3614 (
            .O(N__16981),
            .I(\Lab_UT.dicLdMones_1 ));
    LocalMux I__3613 (
            .O(N__16978),
            .I(\Lab_UT.dicLdMones_1 ));
    LocalMux I__3612 (
            .O(N__16975),
            .I(\Lab_UT.dicLdMones_1 ));
    Odrv4 I__3611 (
            .O(N__16972),
            .I(\Lab_UT.dicLdMones_1 ));
    Odrv4 I__3610 (
            .O(N__16967),
            .I(\Lab_UT.dicLdMones_1 ));
    CascadeMux I__3609 (
            .O(N__16956),
            .I(\Lab_UT.dictrl.N_1300_0_cascade_ ));
    InMux I__3608 (
            .O(N__16953),
            .I(N__16950));
    LocalMux I__3607 (
            .O(N__16950),
            .I(\Lab_UT.dictrl.g1_2_0 ));
    CascadeMux I__3606 (
            .O(N__16947),
            .I(\Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_ ));
    InMux I__3605 (
            .O(N__16944),
            .I(N__16934));
    InMux I__3604 (
            .O(N__16943),
            .I(N__16934));
    InMux I__3603 (
            .O(N__16942),
            .I(N__16934));
    InMux I__3602 (
            .O(N__16941),
            .I(N__16931));
    LocalMux I__3601 (
            .O(N__16934),
            .I(N__16928));
    LocalMux I__3600 (
            .O(N__16931),
            .I(buart__rx_shifter_0_fast_2));
    Odrv4 I__3599 (
            .O(N__16928),
            .I(buart__rx_shifter_0_fast_2));
    InMux I__3598 (
            .O(N__16923),
            .I(N__16920));
    LocalMux I__3597 (
            .O(N__16920),
            .I(\Lab_UT.dictrl.g0_5_5 ));
    InMux I__3596 (
            .O(N__16917),
            .I(N__16914));
    LocalMux I__3595 (
            .O(N__16914),
            .I(\Lab_UT.dictrl.N_7 ));
    InMux I__3594 (
            .O(N__16911),
            .I(N__16908));
    LocalMux I__3593 (
            .O(N__16908),
            .I(\Lab_UT.dictrl.g0_4_a4_4 ));
    InMux I__3592 (
            .O(N__16905),
            .I(N__16902));
    LocalMux I__3591 (
            .O(N__16902),
            .I(\Lab_UT.dictrl.N_5_2 ));
    InMux I__3590 (
            .O(N__16899),
            .I(N__16896));
    LocalMux I__3589 (
            .O(N__16896),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6 ));
    CascadeMux I__3588 (
            .O(N__16893),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_ ));
    CascadeMux I__3587 (
            .O(N__16890),
            .I(\Lab_UT.dictrl.N_96_1_cascade_ ));
    InMux I__3586 (
            .O(N__16887),
            .I(N__16884));
    LocalMux I__3585 (
            .O(N__16884),
            .I(\Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3 ));
    InMux I__3584 (
            .O(N__16881),
            .I(N__16877));
    InMux I__3583 (
            .O(N__16880),
            .I(N__16874));
    LocalMux I__3582 (
            .O(N__16877),
            .I(N__16871));
    LocalMux I__3581 (
            .O(N__16874),
            .I(\Lab_UT.dictrl.m36_0 ));
    Odrv4 I__3580 (
            .O(N__16871),
            .I(\Lab_UT.dictrl.m36_0 ));
    InMux I__3579 (
            .O(N__16866),
            .I(N__16860));
    InMux I__3578 (
            .O(N__16865),
            .I(N__16860));
    LocalMux I__3577 (
            .O(N__16860),
            .I(N__16857));
    Odrv4 I__3576 (
            .O(N__16857),
            .I(\Lab_UT.dictrl.g1_5_0 ));
    InMux I__3575 (
            .O(N__16854),
            .I(N__16851));
    LocalMux I__3574 (
            .O(N__16851),
            .I(\Lab_UT.dictrl.m45_1 ));
    InMux I__3573 (
            .O(N__16848),
            .I(N__16843));
    InMux I__3572 (
            .O(N__16847),
            .I(N__16838));
    InMux I__3571 (
            .O(N__16846),
            .I(N__16838));
    LocalMux I__3570 (
            .O(N__16843),
            .I(N__16832));
    LocalMux I__3569 (
            .O(N__16838),
            .I(N__16832));
    InMux I__3568 (
            .O(N__16837),
            .I(N__16829));
    Span4Mux_h I__3567 (
            .O(N__16832),
            .I(N__16824));
    LocalMux I__3566 (
            .O(N__16829),
            .I(N__16821));
    InMux I__3565 (
            .O(N__16828),
            .I(N__16818));
    InMux I__3564 (
            .O(N__16827),
            .I(N__16815));
    Odrv4 I__3563 (
            .O(N__16824),
            .I(\Lab_UT.dictrl.m25Z0Z_0 ));
    Odrv4 I__3562 (
            .O(N__16821),
            .I(\Lab_UT.dictrl.m25Z0Z_0 ));
    LocalMux I__3561 (
            .O(N__16818),
            .I(\Lab_UT.dictrl.m25Z0Z_0 ));
    LocalMux I__3560 (
            .O(N__16815),
            .I(\Lab_UT.dictrl.m25Z0Z_0 ));
    InMux I__3559 (
            .O(N__16806),
            .I(N__16803));
    LocalMux I__3558 (
            .O(N__16803),
            .I(N__16800));
    Odrv4 I__3557 (
            .O(N__16800),
            .I(\Lab_UT.dictrl.N_6_0 ));
    InMux I__3556 (
            .O(N__16797),
            .I(N__16794));
    LocalMux I__3555 (
            .O(N__16794),
            .I(N__16791));
    Odrv4 I__3554 (
            .O(N__16791),
            .I(\Lab_UT.dictrl.N_5 ));
    CascadeMux I__3553 (
            .O(N__16788),
            .I(N__16785));
    InMux I__3552 (
            .O(N__16785),
            .I(N__16782));
    LocalMux I__3551 (
            .O(N__16782),
            .I(N__16779));
    Odrv12 I__3550 (
            .O(N__16779),
            .I(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ));
    InMux I__3549 (
            .O(N__16776),
            .I(N__16773));
    LocalMux I__3548 (
            .O(N__16773),
            .I(\Lab_UT.dictrl.state_i_4_2 ));
    InMux I__3547 (
            .O(N__16770),
            .I(N__16750));
    InMux I__3546 (
            .O(N__16769),
            .I(N__16750));
    InMux I__3545 (
            .O(N__16768),
            .I(N__16750));
    InMux I__3544 (
            .O(N__16767),
            .I(N__16750));
    InMux I__3543 (
            .O(N__16766),
            .I(N__16750));
    InMux I__3542 (
            .O(N__16765),
            .I(N__16745));
    InMux I__3541 (
            .O(N__16764),
            .I(N__16745));
    InMux I__3540 (
            .O(N__16763),
            .I(N__16738));
    InMux I__3539 (
            .O(N__16762),
            .I(N__16738));
    InMux I__3538 (
            .O(N__16761),
            .I(N__16738));
    LocalMux I__3537 (
            .O(N__16750),
            .I(N__16733));
    LocalMux I__3536 (
            .O(N__16745),
            .I(N__16733));
    LocalMux I__3535 (
            .O(N__16738),
            .I(N__16730));
    Span4Mux_h I__3534 (
            .O(N__16733),
            .I(N__16727));
    Odrv4 I__3533 (
            .O(N__16730),
            .I(\Lab_UT.dicLdAMones_2 ));
    Odrv4 I__3532 (
            .O(N__16727),
            .I(\Lab_UT.dicLdAMones_2 ));
    InMux I__3531 (
            .O(N__16722),
            .I(N__16719));
    LocalMux I__3530 (
            .O(N__16719),
            .I(N__16715));
    InMux I__3529 (
            .O(N__16718),
            .I(N__16712));
    Span4Mux_h I__3528 (
            .O(N__16715),
            .I(N__16709));
    LocalMux I__3527 (
            .O(N__16712),
            .I(\Lab_UT.dictrl.N_94_0 ));
    Odrv4 I__3526 (
            .O(N__16709),
            .I(\Lab_UT.dictrl.N_94_0 ));
    InMux I__3525 (
            .O(N__16704),
            .I(N__16701));
    LocalMux I__3524 (
            .O(N__16701),
            .I(\Lab_UT.dictrl.N_2000_0 ));
    InMux I__3523 (
            .O(N__16698),
            .I(N__16695));
    LocalMux I__3522 (
            .O(N__16695),
            .I(N__16692));
    Odrv4 I__3521 (
            .O(N__16692),
            .I(\Lab_UT.dictrl.g1 ));
    InMux I__3520 (
            .O(N__16689),
            .I(N__16686));
    LocalMux I__3519 (
            .O(N__16686),
            .I(\Lab_UT.dictrl.g1_3_1 ));
    InMux I__3518 (
            .O(N__16683),
            .I(N__16679));
    InMux I__3517 (
            .O(N__16682),
            .I(N__16676));
    LocalMux I__3516 (
            .O(N__16679),
            .I(N__16673));
    LocalMux I__3515 (
            .O(N__16676),
            .I(N__16670));
    Span4Mux_v I__3514 (
            .O(N__16673),
            .I(N__16667));
    Span4Mux_v I__3513 (
            .O(N__16670),
            .I(N__16664));
    Odrv4 I__3512 (
            .O(N__16667),
            .I(\Lab_UT.dictrl.N_88_0 ));
    Odrv4 I__3511 (
            .O(N__16664),
            .I(\Lab_UT.dictrl.N_88_0 ));
    CascadeMux I__3510 (
            .O(N__16659),
            .I(\Lab_UT.dictrl.g1Z0Z_1_cascade_ ));
    CascadeMux I__3509 (
            .O(N__16656),
            .I(\Lab_UT.dictrl.i9_mux_0_1_0_cascade_ ));
    InMux I__3508 (
            .O(N__16653),
            .I(N__16650));
    LocalMux I__3507 (
            .O(N__16650),
            .I(\Lab_UT.dictrl.N_94_0_1_0 ));
    CascadeMux I__3506 (
            .O(N__16647),
            .I(\Lab_UT.dictrl.N_2000_0_1_0_cascade_ ));
    InMux I__3505 (
            .O(N__16644),
            .I(N__16641));
    LocalMux I__3504 (
            .O(N__16641),
            .I(N__16638));
    Span4Mux_h I__3503 (
            .O(N__16638),
            .I(N__16630));
    InMux I__3502 (
            .O(N__16637),
            .I(N__16627));
    InMux I__3501 (
            .O(N__16636),
            .I(N__16624));
    InMux I__3500 (
            .O(N__16635),
            .I(N__16611));
    InMux I__3499 (
            .O(N__16634),
            .I(N__16611));
    InMux I__3498 (
            .O(N__16633),
            .I(N__16611));
    Span4Mux_v I__3497 (
            .O(N__16630),
            .I(N__16608));
    LocalMux I__3496 (
            .O(N__16627),
            .I(N__16605));
    LocalMux I__3495 (
            .O(N__16624),
            .I(N__16602));
    InMux I__3494 (
            .O(N__16623),
            .I(N__16595));
    InMux I__3493 (
            .O(N__16622),
            .I(N__16595));
    InMux I__3492 (
            .O(N__16621),
            .I(N__16595));
    InMux I__3491 (
            .O(N__16620),
            .I(N__16590));
    InMux I__3490 (
            .O(N__16619),
            .I(N__16590));
    InMux I__3489 (
            .O(N__16618),
            .I(N__16587));
    LocalMux I__3488 (
            .O(N__16611),
            .I(N__16582));
    Span4Mux_h I__3487 (
            .O(N__16608),
            .I(N__16582));
    Odrv12 I__3486 (
            .O(N__16605),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__3485 (
            .O(N__16602),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__3484 (
            .O(N__16595),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__3483 (
            .O(N__16590),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__3482 (
            .O(N__16587),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__3481 (
            .O(N__16582),
            .I(\uu0.un4_l_count_0 ));
    IoInMux I__3480 (
            .O(N__16569),
            .I(N__16566));
    LocalMux I__3479 (
            .O(N__16566),
            .I(N__16563));
    IoSpan4Mux I__3478 (
            .O(N__16563),
            .I(N__16560));
    Span4Mux_s1_h I__3477 (
            .O(N__16560),
            .I(N__16557));
    Span4Mux_h I__3476 (
            .O(N__16557),
            .I(N__16554));
    Odrv4 I__3475 (
            .O(N__16554),
            .I(\uu0.un11_l_count_i ));
    InMux I__3474 (
            .O(N__16551),
            .I(N__16538));
    InMux I__3473 (
            .O(N__16550),
            .I(N__16538));
    InMux I__3472 (
            .O(N__16549),
            .I(N__16538));
    InMux I__3471 (
            .O(N__16548),
            .I(N__16538));
    InMux I__3470 (
            .O(N__16547),
            .I(N__16535));
    LocalMux I__3469 (
            .O(N__16538),
            .I(N__16532));
    LocalMux I__3468 (
            .O(N__16535),
            .I(N__16529));
    Span4Mux_h I__3467 (
            .O(N__16532),
            .I(N__16524));
    Span4Mux_h I__3466 (
            .O(N__16529),
            .I(N__16524));
    Odrv4 I__3465 (
            .O(N__16524),
            .I(\Lab_UT.dicLdASones_0 ));
    CascadeMux I__3464 (
            .O(N__16521),
            .I(N__16518));
    InMux I__3463 (
            .O(N__16518),
            .I(N__16515));
    LocalMux I__3462 (
            .O(N__16515),
            .I(\Lab_UT.dictrl.g3_1 ));
    CascadeMux I__3461 (
            .O(N__16512),
            .I(\Lab_UT.dictrl.i9_mux_0_cascade_ ));
    CascadeMux I__3460 (
            .O(N__16509),
            .I(\Lab_UT.dictrl.N_2000_0_cascade_ ));
    CascadeMux I__3459 (
            .O(N__16506),
            .I(\resetGen.un241_ci_cascade_ ));
    CascadeMux I__3458 (
            .O(N__16503),
            .I(N__16500));
    InMux I__3457 (
            .O(N__16500),
            .I(N__16494));
    InMux I__3456 (
            .O(N__16499),
            .I(N__16494));
    LocalMux I__3455 (
            .O(N__16494),
            .I(\resetGen.reset_countZ0Z_3 ));
    CascadeMux I__3454 (
            .O(N__16491),
            .I(\resetGen.reset_count_2_0_4_cascade_ ));
    InMux I__3453 (
            .O(N__16488),
            .I(N__16485));
    LocalMux I__3452 (
            .O(N__16485),
            .I(\resetGen.un241_ci ));
    CascadeMux I__3451 (
            .O(N__16482),
            .I(N__16475));
    InMux I__3450 (
            .O(N__16481),
            .I(N__16471));
    InMux I__3449 (
            .O(N__16480),
            .I(N__16460));
    InMux I__3448 (
            .O(N__16479),
            .I(N__16460));
    InMux I__3447 (
            .O(N__16478),
            .I(N__16460));
    InMux I__3446 (
            .O(N__16475),
            .I(N__16460));
    InMux I__3445 (
            .O(N__16474),
            .I(N__16460));
    LocalMux I__3444 (
            .O(N__16471),
            .I(N__16457));
    LocalMux I__3443 (
            .O(N__16460),
            .I(\resetGen.reset_countZ0Z_4 ));
    Odrv4 I__3442 (
            .O(N__16457),
            .I(\resetGen.reset_countZ0Z_4 ));
    CascadeMux I__3441 (
            .O(N__16452),
            .I(N__16446));
    CascadeMux I__3440 (
            .O(N__16451),
            .I(N__16441));
    CascadeMux I__3439 (
            .O(N__16450),
            .I(N__16437));
    InMux I__3438 (
            .O(N__16449),
            .I(N__16433));
    InMux I__3437 (
            .O(N__16446),
            .I(N__16418));
    InMux I__3436 (
            .O(N__16445),
            .I(N__16418));
    InMux I__3435 (
            .O(N__16444),
            .I(N__16418));
    InMux I__3434 (
            .O(N__16441),
            .I(N__16418));
    InMux I__3433 (
            .O(N__16440),
            .I(N__16418));
    InMux I__3432 (
            .O(N__16437),
            .I(N__16418));
    InMux I__3431 (
            .O(N__16436),
            .I(N__16418));
    LocalMux I__3430 (
            .O(N__16433),
            .I(N__16414));
    LocalMux I__3429 (
            .O(N__16418),
            .I(N__16411));
    CascadeMux I__3428 (
            .O(N__16417),
            .I(N__16408));
    Span4Mux_h I__3427 (
            .O(N__16414),
            .I(N__16404));
    Span4Mux_v I__3426 (
            .O(N__16411),
            .I(N__16401));
    InMux I__3425 (
            .O(N__16408),
            .I(N__16398));
    InMux I__3424 (
            .O(N__16407),
            .I(N__16395));
    Span4Mux_v I__3423 (
            .O(N__16404),
            .I(N__16392));
    Odrv4 I__3422 (
            .O(N__16401),
            .I(\Lab_UT.dicRun_1 ));
    LocalMux I__3421 (
            .O(N__16398),
            .I(\Lab_UT.dicRun_1 ));
    LocalMux I__3420 (
            .O(N__16395),
            .I(\Lab_UT.dicRun_1 ));
    Odrv4 I__3419 (
            .O(N__16392),
            .I(\Lab_UT.dicRun_1 ));
    InMux I__3418 (
            .O(N__16383),
            .I(N__16376));
    InMux I__3417 (
            .O(N__16382),
            .I(N__16376));
    InMux I__3416 (
            .O(N__16381),
            .I(N__16373));
    LocalMux I__3415 (
            .O(N__16376),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__3414 (
            .O(N__16373),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__3413 (
            .O(N__16368),
            .I(N__16364));
    InMux I__3412 (
            .O(N__16367),
            .I(N__16359));
    InMux I__3411 (
            .O(N__16364),
            .I(N__16356));
    InMux I__3410 (
            .O(N__16363),
            .I(N__16351));
    InMux I__3409 (
            .O(N__16362),
            .I(N__16351));
    LocalMux I__3408 (
            .O(N__16359),
            .I(N__16348));
    LocalMux I__3407 (
            .O(N__16356),
            .I(\resetGen.reset_countZ0Z_0 ));
    LocalMux I__3406 (
            .O(N__16351),
            .I(\resetGen.reset_countZ0Z_0 ));
    Odrv4 I__3405 (
            .O(N__16348),
            .I(\resetGen.reset_countZ0Z_0 ));
    InMux I__3404 (
            .O(N__16341),
            .I(N__16336));
    InMux I__3403 (
            .O(N__16340),
            .I(N__16331));
    InMux I__3402 (
            .O(N__16339),
            .I(N__16331));
    LocalMux I__3401 (
            .O(N__16336),
            .I(\resetGen.reset_countZ0Z_2 ));
    LocalMux I__3400 (
            .O(N__16331),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__3399 (
            .O(N__16326),
            .I(N__16323));
    LocalMux I__3398 (
            .O(N__16323),
            .I(\resetGen.un252_ci ));
    InMux I__3397 (
            .O(N__16320),
            .I(N__16317));
    LocalMux I__3396 (
            .O(N__16317),
            .I(N__16313));
    InMux I__3395 (
            .O(N__16316),
            .I(N__16310));
    Sp12to4 I__3394 (
            .O(N__16313),
            .I(N__16307));
    LocalMux I__3393 (
            .O(N__16310),
            .I(N__16304));
    Span12Mux_s9_v I__3392 (
            .O(N__16307),
            .I(N__16301));
    Odrv4 I__3391 (
            .O(N__16304),
            .I(\uu0.delay_lineZ0Z_0 ));
    Odrv12 I__3390 (
            .O(N__16301),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__3389 (
            .O(N__16296),
            .I(N__16293));
    LocalMux I__3388 (
            .O(N__16293),
            .I(N__16290));
    Span4Mux_h I__3387 (
            .O(N__16290),
            .I(N__16287));
    Span4Mux_h I__3386 (
            .O(N__16287),
            .I(N__16284));
    Odrv4 I__3385 (
            .O(N__16284),
            .I(\uu0.delay_lineZ0Z_1 ));
    CascadeMux I__3384 (
            .O(N__16281),
            .I(N__16277));
    InMux I__3383 (
            .O(N__16280),
            .I(N__16274));
    InMux I__3382 (
            .O(N__16277),
            .I(N__16271));
    LocalMux I__3381 (
            .O(N__16274),
            .I(N__16264));
    LocalMux I__3380 (
            .O(N__16271),
            .I(N__16264));
    InMux I__3379 (
            .O(N__16270),
            .I(N__16261));
    InMux I__3378 (
            .O(N__16269),
            .I(N__16258));
    Span4Mux_h I__3377 (
            .O(N__16264),
            .I(N__16255));
    LocalMux I__3376 (
            .O(N__16261),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    LocalMux I__3375 (
            .O(N__16258),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    Odrv4 I__3374 (
            .O(N__16255),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    InMux I__3373 (
            .O(N__16248),
            .I(N__16245));
    LocalMux I__3372 (
            .O(N__16245),
            .I(N__16242));
    Span4Mux_s2_v I__3371 (
            .O(N__16242),
            .I(N__16238));
    InMux I__3370 (
            .O(N__16241),
            .I(N__16235));
    Odrv4 I__3369 (
            .O(N__16238),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    LocalMux I__3368 (
            .O(N__16235),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__3367 (
            .O(N__16230),
            .I(N__16225));
    InMux I__3366 (
            .O(N__16229),
            .I(N__16220));
    InMux I__3365 (
            .O(N__16228),
            .I(N__16220));
    LocalMux I__3364 (
            .O(N__16225),
            .I(\Lab_UT.didp.countrce3.ce_12_2_3 ));
    LocalMux I__3363 (
            .O(N__16220),
            .I(\Lab_UT.didp.countrce3.ce_12_2_3 ));
    CascadeMux I__3362 (
            .O(N__16215),
            .I(N__16210));
    CascadeMux I__3361 (
            .O(N__16214),
            .I(N__16206));
    CascadeMux I__3360 (
            .O(N__16213),
            .I(N__16202));
    InMux I__3359 (
            .O(N__16210),
            .I(N__16197));
    InMux I__3358 (
            .O(N__16209),
            .I(N__16197));
    InMux I__3357 (
            .O(N__16206),
            .I(N__16190));
    InMux I__3356 (
            .O(N__16205),
            .I(N__16190));
    InMux I__3355 (
            .O(N__16202),
            .I(N__16190));
    LocalMux I__3354 (
            .O(N__16197),
            .I(N__16185));
    LocalMux I__3353 (
            .O(N__16190),
            .I(N__16185));
    Odrv12 I__3352 (
            .O(N__16185),
            .I(\Lab_UT.didp.un24_ce_2 ));
    InMux I__3351 (
            .O(N__16182),
            .I(N__16179));
    LocalMux I__3350 (
            .O(N__16179),
            .I(\Lab_UT.didp.reset_12_1_3 ));
    InMux I__3349 (
            .O(N__16176),
            .I(N__16172));
    InMux I__3348 (
            .O(N__16175),
            .I(N__16168));
    LocalMux I__3347 (
            .O(N__16172),
            .I(N__16165));
    InMux I__3346 (
            .O(N__16171),
            .I(N__16160));
    LocalMux I__3345 (
            .O(N__16168),
            .I(N__16154));
    Span4Mux_s3_v I__3344 (
            .O(N__16165),
            .I(N__16154));
    InMux I__3343 (
            .O(N__16164),
            .I(N__16149));
    InMux I__3342 (
            .O(N__16163),
            .I(N__16149));
    LocalMux I__3341 (
            .O(N__16160),
            .I(N__16146));
    InMux I__3340 (
            .O(N__16159),
            .I(N__16143));
    Odrv4 I__3339 (
            .O(N__16154),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__3338 (
            .O(N__16149),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    Odrv4 I__3337 (
            .O(N__16146),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__3336 (
            .O(N__16143),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    CascadeMux I__3335 (
            .O(N__16134),
            .I(\Lab_UT.didp.ce_12_3_cascade_ ));
    InMux I__3334 (
            .O(N__16131),
            .I(N__16125));
    CascadeMux I__3333 (
            .O(N__16130),
            .I(N__16122));
    CascadeMux I__3332 (
            .O(N__16129),
            .I(N__16119));
    CascadeMux I__3331 (
            .O(N__16128),
            .I(N__16115));
    LocalMux I__3330 (
            .O(N__16125),
            .I(N__16112));
    InMux I__3329 (
            .O(N__16122),
            .I(N__16109));
    InMux I__3328 (
            .O(N__16119),
            .I(N__16106));
    InMux I__3327 (
            .O(N__16118),
            .I(N__16103));
    InMux I__3326 (
            .O(N__16115),
            .I(N__16100));
    Span4Mux_h I__3325 (
            .O(N__16112),
            .I(N__16093));
    LocalMux I__3324 (
            .O(N__16109),
            .I(N__16093));
    LocalMux I__3323 (
            .O(N__16106),
            .I(N__16093));
    LocalMux I__3322 (
            .O(N__16103),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    LocalMux I__3321 (
            .O(N__16100),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    Odrv4 I__3320 (
            .O(N__16093),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    InMux I__3319 (
            .O(N__16086),
            .I(N__16083));
    LocalMux I__3318 (
            .O(N__16083),
            .I(N__16077));
    InMux I__3317 (
            .O(N__16082),
            .I(N__16070));
    InMux I__3316 (
            .O(N__16081),
            .I(N__16070));
    InMux I__3315 (
            .O(N__16080),
            .I(N__16070));
    Span4Mux_h I__3314 (
            .O(N__16077),
            .I(N__16065));
    LocalMux I__3313 (
            .O(N__16070),
            .I(N__16065));
    Odrv4 I__3312 (
            .O(N__16065),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    InMux I__3311 (
            .O(N__16062),
            .I(N__16041));
    InMux I__3310 (
            .O(N__16061),
            .I(N__16041));
    InMux I__3309 (
            .O(N__16060),
            .I(N__16041));
    InMux I__3308 (
            .O(N__16059),
            .I(N__16041));
    InMux I__3307 (
            .O(N__16058),
            .I(N__16041));
    InMux I__3306 (
            .O(N__16057),
            .I(N__16041));
    InMux I__3305 (
            .O(N__16056),
            .I(N__16041));
    LocalMux I__3304 (
            .O(N__16041),
            .I(N__16038));
    Odrv4 I__3303 (
            .O(N__16038),
            .I(\Lab_UT.didp.un18_ce ));
    InMux I__3302 (
            .O(N__16035),
            .I(N__16014));
    InMux I__3301 (
            .O(N__16034),
            .I(N__16014));
    InMux I__3300 (
            .O(N__16033),
            .I(N__16014));
    InMux I__3299 (
            .O(N__16032),
            .I(N__16014));
    InMux I__3298 (
            .O(N__16031),
            .I(N__16014));
    InMux I__3297 (
            .O(N__16030),
            .I(N__16014));
    InMux I__3296 (
            .O(N__16029),
            .I(N__16014));
    LocalMux I__3295 (
            .O(N__16014),
            .I(N__16009));
    CascadeMux I__3294 (
            .O(N__16013),
            .I(N__16004));
    InMux I__3293 (
            .O(N__16012),
            .I(N__16001));
    Span4Mux_h I__3292 (
            .O(N__16009),
            .I(N__15998));
    InMux I__3291 (
            .O(N__16008),
            .I(N__15995));
    CascadeMux I__3290 (
            .O(N__16007),
            .I(N__15990));
    InMux I__3289 (
            .O(N__16004),
            .I(N__15985));
    LocalMux I__3288 (
            .O(N__16001),
            .I(N__15982));
    Span4Mux_v I__3287 (
            .O(N__15998),
            .I(N__15977));
    LocalMux I__3286 (
            .O(N__15995),
            .I(N__15977));
    InMux I__3285 (
            .O(N__15994),
            .I(N__15972));
    InMux I__3284 (
            .O(N__15993),
            .I(N__15972));
    InMux I__3283 (
            .O(N__15990),
            .I(N__15969));
    InMux I__3282 (
            .O(N__15989),
            .I(N__15964));
    InMux I__3281 (
            .O(N__15988),
            .I(N__15964));
    LocalMux I__3280 (
            .O(N__15985),
            .I(N__15961));
    Span4Mux_v I__3279 (
            .O(N__15982),
            .I(N__15958));
    Span4Mux_v I__3278 (
            .O(N__15977),
            .I(N__15953));
    LocalMux I__3277 (
            .O(N__15972),
            .I(N__15953));
    LocalMux I__3276 (
            .O(N__15969),
            .I(N__15948));
    LocalMux I__3275 (
            .O(N__15964),
            .I(N__15948));
    Span4Mux_v I__3274 (
            .O(N__15961),
            .I(N__15945));
    Span4Mux_h I__3273 (
            .O(N__15958),
            .I(N__15942));
    Span4Mux_h I__3272 (
            .O(N__15953),
            .I(N__15939));
    Odrv4 I__3271 (
            .O(N__15948),
            .I(oneSecStrb));
    Odrv4 I__3270 (
            .O(N__15945),
            .I(oneSecStrb));
    Odrv4 I__3269 (
            .O(N__15942),
            .I(oneSecStrb));
    Odrv4 I__3268 (
            .O(N__15939),
            .I(oneSecStrb));
    InMux I__3267 (
            .O(N__15930),
            .I(N__15924));
    InMux I__3266 (
            .O(N__15929),
            .I(N__15924));
    LocalMux I__3265 (
            .O(N__15924),
            .I(N__15919));
    InMux I__3264 (
            .O(N__15923),
            .I(N__15914));
    InMux I__3263 (
            .O(N__15922),
            .I(N__15914));
    Span4Mux_h I__3262 (
            .O(N__15919),
            .I(N__15909));
    LocalMux I__3261 (
            .O(N__15914),
            .I(N__15909));
    Span4Mux_s0_v I__3260 (
            .O(N__15909),
            .I(N__15906));
    Odrv4 I__3259 (
            .O(N__15906),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    InMux I__3258 (
            .O(N__15903),
            .I(N__15897));
    InMux I__3257 (
            .O(N__15902),
            .I(N__15892));
    InMux I__3256 (
            .O(N__15901),
            .I(N__15889));
    InMux I__3255 (
            .O(N__15900),
            .I(N__15886));
    LocalMux I__3254 (
            .O(N__15897),
            .I(N__15883));
    InMux I__3253 (
            .O(N__15896),
            .I(N__15878));
    InMux I__3252 (
            .O(N__15895),
            .I(N__15878));
    LocalMux I__3251 (
            .O(N__15892),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3250 (
            .O(N__15889),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3249 (
            .O(N__15886),
            .I(\Lab_UT.didp.di_Mones_1 ));
    Odrv4 I__3248 (
            .O(N__15883),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3247 (
            .O(N__15878),
            .I(\Lab_UT.didp.di_Mones_1 ));
    InMux I__3246 (
            .O(N__15867),
            .I(N__15861));
    InMux I__3245 (
            .O(N__15866),
            .I(N__15861));
    LocalMux I__3244 (
            .O(N__15861),
            .I(N__15854));
    InMux I__3243 (
            .O(N__15860),
            .I(N__15851));
    InMux I__3242 (
            .O(N__15859),
            .I(N__15844));
    InMux I__3241 (
            .O(N__15858),
            .I(N__15844));
    InMux I__3240 (
            .O(N__15857),
            .I(N__15844));
    Odrv4 I__3239 (
            .O(N__15854),
            .I(\Lab_UT.didp.di_Mones_0 ));
    LocalMux I__3238 (
            .O(N__15851),
            .I(\Lab_UT.didp.di_Mones_0 ));
    LocalMux I__3237 (
            .O(N__15844),
            .I(\Lab_UT.didp.di_Mones_0 ));
    CascadeMux I__3236 (
            .O(N__15837),
            .I(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ));
    CascadeMux I__3235 (
            .O(N__15834),
            .I(\Lab_UT.didp.countrce3.q_5_2_cascade_ ));
    InMux I__3234 (
            .O(N__15831),
            .I(N__15828));
    LocalMux I__3233 (
            .O(N__15828),
            .I(\Lab_UT.didp.countrce3.un13_qPone ));
    CascadeMux I__3232 (
            .O(N__15825),
            .I(N__15817));
    InMux I__3231 (
            .O(N__15824),
            .I(N__15814));
    CascadeMux I__3230 (
            .O(N__15823),
            .I(N__15811));
    InMux I__3229 (
            .O(N__15822),
            .I(N__15802));
    InMux I__3228 (
            .O(N__15821),
            .I(N__15802));
    InMux I__3227 (
            .O(N__15820),
            .I(N__15802));
    InMux I__3226 (
            .O(N__15817),
            .I(N__15802));
    LocalMux I__3225 (
            .O(N__15814),
            .I(N__15799));
    InMux I__3224 (
            .O(N__15811),
            .I(N__15796));
    LocalMux I__3223 (
            .O(N__15802),
            .I(\Lab_UT.didp.di_Mones_2 ));
    Odrv4 I__3222 (
            .O(N__15799),
            .I(\Lab_UT.didp.di_Mones_2 ));
    LocalMux I__3221 (
            .O(N__15796),
            .I(\Lab_UT.didp.di_Mones_2 ));
    InMux I__3220 (
            .O(N__15789),
            .I(N__15783));
    InMux I__3219 (
            .O(N__15788),
            .I(N__15780));
    InMux I__3218 (
            .O(N__15787),
            .I(N__15777));
    CascadeMux I__3217 (
            .O(N__15786),
            .I(N__15773));
    LocalMux I__3216 (
            .O(N__15783),
            .I(N__15765));
    LocalMux I__3215 (
            .O(N__15780),
            .I(N__15765));
    LocalMux I__3214 (
            .O(N__15777),
            .I(N__15765));
    InMux I__3213 (
            .O(N__15776),
            .I(N__15758));
    InMux I__3212 (
            .O(N__15773),
            .I(N__15758));
    InMux I__3211 (
            .O(N__15772),
            .I(N__15758));
    Span4Mux_h I__3210 (
            .O(N__15765),
            .I(N__15755));
    LocalMux I__3209 (
            .O(N__15758),
            .I(N__15752));
    Span4Mux_v I__3208 (
            .O(N__15755),
            .I(N__15749));
    Span4Mux_v I__3207 (
            .O(N__15752),
            .I(N__15746));
    Odrv4 I__3206 (
            .O(N__15749),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3205 (
            .O(N__15746),
            .I(\Lab_UT.LdMones ));
    CascadeMux I__3204 (
            .O(N__15741),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    CascadeMux I__3203 (
            .O(N__15738),
            .I(\Lab_UT.didp.countrce3.q_5_3_cascade_ ));
    InMux I__3202 (
            .O(N__15735),
            .I(N__15729));
    InMux I__3201 (
            .O(N__15734),
            .I(N__15729));
    LocalMux I__3200 (
            .O(N__15729),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    InMux I__3199 (
            .O(N__15726),
            .I(N__15719));
    InMux I__3198 (
            .O(N__15725),
            .I(N__15716));
    InMux I__3197 (
            .O(N__15724),
            .I(N__15709));
    InMux I__3196 (
            .O(N__15723),
            .I(N__15709));
    InMux I__3195 (
            .O(N__15722),
            .I(N__15709));
    LocalMux I__3194 (
            .O(N__15719),
            .I(N__15706));
    LocalMux I__3193 (
            .O(N__15716),
            .I(N__15703));
    LocalMux I__3192 (
            .O(N__15709),
            .I(\Lab_UT.didp.di_Mones_3 ));
    Odrv4 I__3191 (
            .O(N__15706),
            .I(\Lab_UT.didp.di_Mones_3 ));
    Odrv4 I__3190 (
            .O(N__15703),
            .I(\Lab_UT.didp.di_Mones_3 ));
    InMux I__3189 (
            .O(N__15696),
            .I(N__15690));
    InMux I__3188 (
            .O(N__15695),
            .I(N__15690));
    LocalMux I__3187 (
            .O(N__15690),
            .I(N__15687));
    Span4Mux_v I__3186 (
            .O(N__15687),
            .I(N__15684));
    Odrv4 I__3185 (
            .O(N__15684),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    InMux I__3184 (
            .O(N__15681),
            .I(N__15674));
    InMux I__3183 (
            .O(N__15680),
            .I(N__15671));
    InMux I__3182 (
            .O(N__15679),
            .I(N__15668));
    InMux I__3181 (
            .O(N__15678),
            .I(N__15663));
    InMux I__3180 (
            .O(N__15677),
            .I(N__15663));
    LocalMux I__3179 (
            .O(N__15674),
            .I(N__15658));
    LocalMux I__3178 (
            .O(N__15671),
            .I(N__15658));
    LocalMux I__3177 (
            .O(N__15668),
            .I(\Lab_UT.dictrl.N_20_0 ));
    LocalMux I__3176 (
            .O(N__15663),
            .I(\Lab_UT.dictrl.N_20_0 ));
    Odrv4 I__3175 (
            .O(N__15658),
            .I(\Lab_UT.dictrl.N_20_0 ));
    InMux I__3174 (
            .O(N__15651),
            .I(N__15648));
    LocalMux I__3173 (
            .O(N__15648),
            .I(N__15645));
    Odrv12 I__3172 (
            .O(N__15645),
            .I(\Lab_UT.dictrl.g0_5_2 ));
    CascadeMux I__3171 (
            .O(N__15642),
            .I(N__15637));
    CascadeMux I__3170 (
            .O(N__15641),
            .I(N__15632));
    InMux I__3169 (
            .O(N__15640),
            .I(N__15629));
    InMux I__3168 (
            .O(N__15637),
            .I(N__15626));
    InMux I__3167 (
            .O(N__15636),
            .I(N__15621));
    InMux I__3166 (
            .O(N__15635),
            .I(N__15621));
    InMux I__3165 (
            .O(N__15632),
            .I(N__15618));
    LocalMux I__3164 (
            .O(N__15629),
            .I(N__15615));
    LocalMux I__3163 (
            .O(N__15626),
            .I(bu_rx_data_i_4_fast_7));
    LocalMux I__3162 (
            .O(N__15621),
            .I(bu_rx_data_i_4_fast_7));
    LocalMux I__3161 (
            .O(N__15618),
            .I(bu_rx_data_i_4_fast_7));
    Odrv4 I__3160 (
            .O(N__15615),
            .I(bu_rx_data_i_4_fast_7));
    CEMux I__3159 (
            .O(N__15606),
            .I(N__15579));
    CEMux I__3158 (
            .O(N__15605),
            .I(N__15579));
    CEMux I__3157 (
            .O(N__15604),
            .I(N__15579));
    CEMux I__3156 (
            .O(N__15603),
            .I(N__15579));
    CEMux I__3155 (
            .O(N__15602),
            .I(N__15579));
    CEMux I__3154 (
            .O(N__15601),
            .I(N__15579));
    CEMux I__3153 (
            .O(N__15600),
            .I(N__15579));
    CEMux I__3152 (
            .O(N__15599),
            .I(N__15579));
    CEMux I__3151 (
            .O(N__15598),
            .I(N__15579));
    GlobalMux I__3150 (
            .O(N__15579),
            .I(N__15576));
    gio2CtrlBuf I__3149 (
            .O(N__15576),
            .I(buart__rx_sample_g));
    InMux I__3148 (
            .O(N__15573),
            .I(N__15569));
    CascadeMux I__3147 (
            .O(N__15572),
            .I(N__15566));
    LocalMux I__3146 (
            .O(N__15569),
            .I(N__15563));
    InMux I__3145 (
            .O(N__15566),
            .I(N__15560));
    Span4Mux_h I__3144 (
            .O(N__15563),
            .I(N__15555));
    LocalMux I__3143 (
            .O(N__15560),
            .I(N__15552));
    InMux I__3142 (
            .O(N__15559),
            .I(N__15549));
    InMux I__3141 (
            .O(N__15558),
            .I(N__15546));
    Span4Mux_v I__3140 (
            .O(N__15555),
            .I(N__15543));
    Span4Mux_s2_v I__3139 (
            .O(N__15552),
            .I(N__15540));
    LocalMux I__3138 (
            .O(N__15549),
            .I(N__15537));
    LocalMux I__3137 (
            .O(N__15546),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__3136 (
            .O(N__15543),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__3135 (
            .O(N__15540),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__3134 (
            .O(N__15537),
            .I(\Lab_UT.di_AStens_1 ));
    CascadeMux I__3133 (
            .O(N__15528),
            .I(N__15525));
    InMux I__3132 (
            .O(N__15525),
            .I(N__15521));
    CascadeMux I__3131 (
            .O(N__15524),
            .I(N__15518));
    LocalMux I__3130 (
            .O(N__15521),
            .I(N__15513));
    InMux I__3129 (
            .O(N__15518),
            .I(N__15510));
    CascadeMux I__3128 (
            .O(N__15517),
            .I(N__15507));
    CascadeMux I__3127 (
            .O(N__15516),
            .I(N__15504));
    Span4Mux_h I__3126 (
            .O(N__15513),
            .I(N__15501));
    LocalMux I__3125 (
            .O(N__15510),
            .I(N__15498));
    InMux I__3124 (
            .O(N__15507),
            .I(N__15495));
    InMux I__3123 (
            .O(N__15504),
            .I(N__15492));
    Span4Mux_v I__3122 (
            .O(N__15501),
            .I(N__15487));
    Span4Mux_h I__3121 (
            .O(N__15498),
            .I(N__15487));
    LocalMux I__3120 (
            .O(N__15495),
            .I(N__15484));
    LocalMux I__3119 (
            .O(N__15492),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__3118 (
            .O(N__15487),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__3117 (
            .O(N__15484),
            .I(\Lab_UT.di_AStens_2 ));
    InMux I__3116 (
            .O(N__15477),
            .I(N__15474));
    LocalMux I__3115 (
            .O(N__15474),
            .I(N__15471));
    Span4Mux_v I__3114 (
            .O(N__15471),
            .I(N__15468));
    Odrv4 I__3113 (
            .O(N__15468),
            .I(\Lab_UT.didp.did_alarmMatch_2 ));
    InMux I__3112 (
            .O(N__15465),
            .I(N__15458));
    InMux I__3111 (
            .O(N__15464),
            .I(N__15454));
    InMux I__3110 (
            .O(N__15463),
            .I(N__15447));
    InMux I__3109 (
            .O(N__15462),
            .I(N__15447));
    InMux I__3108 (
            .O(N__15461),
            .I(N__15447));
    LocalMux I__3107 (
            .O(N__15458),
            .I(N__15444));
    InMux I__3106 (
            .O(N__15457),
            .I(N__15441));
    LocalMux I__3105 (
            .O(N__15454),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__3104 (
            .O(N__15447),
            .I(\Lab_UT.didp.di_Sones_1 ));
    Odrv4 I__3103 (
            .O(N__15444),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__3102 (
            .O(N__15441),
            .I(\Lab_UT.didp.di_Sones_1 ));
    InMux I__3101 (
            .O(N__15432),
            .I(N__15425));
    InMux I__3100 (
            .O(N__15431),
            .I(N__15422));
    InMux I__3099 (
            .O(N__15430),
            .I(N__15419));
    InMux I__3098 (
            .O(N__15429),
            .I(N__15416));
    InMux I__3097 (
            .O(N__15428),
            .I(N__15413));
    LocalMux I__3096 (
            .O(N__15425),
            .I(N__15410));
    LocalMux I__3095 (
            .O(N__15422),
            .I(N__15405));
    LocalMux I__3094 (
            .O(N__15419),
            .I(N__15405));
    LocalMux I__3093 (
            .O(N__15416),
            .I(\Lab_UT.didp.di_Sones_3 ));
    LocalMux I__3092 (
            .O(N__15413),
            .I(\Lab_UT.didp.di_Sones_3 ));
    Odrv4 I__3091 (
            .O(N__15410),
            .I(\Lab_UT.didp.di_Sones_3 ));
    Odrv4 I__3090 (
            .O(N__15405),
            .I(\Lab_UT.didp.di_Sones_3 ));
    CascadeMux I__3089 (
            .O(N__15396),
            .I(N__15391));
    InMux I__3088 (
            .O(N__15395),
            .I(N__15385));
    InMux I__3087 (
            .O(N__15394),
            .I(N__15385));
    InMux I__3086 (
            .O(N__15391),
            .I(N__15382));
    InMux I__3085 (
            .O(N__15390),
            .I(N__15379));
    LocalMux I__3084 (
            .O(N__15385),
            .I(N__15372));
    LocalMux I__3083 (
            .O(N__15382),
            .I(N__15372));
    LocalMux I__3082 (
            .O(N__15379),
            .I(N__15369));
    InMux I__3081 (
            .O(N__15378),
            .I(N__15364));
    InMux I__3080 (
            .O(N__15377),
            .I(N__15364));
    Odrv4 I__3079 (
            .O(N__15372),
            .I(\Lab_UT.didp.di_Sones_2 ));
    Odrv4 I__3078 (
            .O(N__15369),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__3077 (
            .O(N__15364),
            .I(\Lab_UT.didp.di_Sones_2 ));
    InMux I__3076 (
            .O(N__15357),
            .I(N__15354));
    LocalMux I__3075 (
            .O(N__15354),
            .I(\Lab_UT.dictrl.g1_1_1_0 ));
    InMux I__3074 (
            .O(N__15351),
            .I(N__15345));
    InMux I__3073 (
            .O(N__15350),
            .I(N__15345));
    LocalMux I__3072 (
            .O(N__15345),
            .I(N__15340));
    InMux I__3071 (
            .O(N__15344),
            .I(N__15337));
    InMux I__3070 (
            .O(N__15343),
            .I(N__15334));
    Odrv4 I__3069 (
            .O(N__15340),
            .I(bu_rx_data_fast_4));
    LocalMux I__3068 (
            .O(N__15337),
            .I(bu_rx_data_fast_4));
    LocalMux I__3067 (
            .O(N__15334),
            .I(bu_rx_data_fast_4));
    InMux I__3066 (
            .O(N__15327),
            .I(N__15324));
    LocalMux I__3065 (
            .O(N__15324),
            .I(\Lab_UT.dictrl.N_98_mux_0 ));
    CascadeMux I__3064 (
            .O(N__15321),
            .I(\Lab_UT.dictrl.g0_3_1_0_cascade_ ));
    InMux I__3063 (
            .O(N__15318),
            .I(N__15315));
    LocalMux I__3062 (
            .O(N__15315),
            .I(\Lab_UT.dictrl.g0_4Z0Z_1 ));
    CascadeMux I__3061 (
            .O(N__15312),
            .I(N__15307));
    InMux I__3060 (
            .O(N__15311),
            .I(N__15302));
    InMux I__3059 (
            .O(N__15310),
            .I(N__15302));
    InMux I__3058 (
            .O(N__15307),
            .I(N__15299));
    LocalMux I__3057 (
            .O(N__15302),
            .I(buart__rx_shifter_ret_1_fast));
    LocalMux I__3056 (
            .O(N__15299),
            .I(buart__rx_shifter_ret_1_fast));
    CascadeMux I__3055 (
            .O(N__15294),
            .I(\Lab_UT.dictrl.m25_xZ0Z1_cascade_ ));
    CascadeMux I__3054 (
            .O(N__15291),
            .I(\Lab_UT.dictrl.N_116_mux_cascade_ ));
    CascadeMux I__3053 (
            .O(N__15288),
            .I(\Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ));
    InMux I__3052 (
            .O(N__15285),
            .I(N__15282));
    LocalMux I__3051 (
            .O(N__15282),
            .I(N__15279));
    Odrv4 I__3050 (
            .O(N__15279),
            .I(\Lab_UT.dictrl.g0_0_0_a3_4 ));
    CascadeMux I__3049 (
            .O(N__15276),
            .I(\Lab_UT.dictrl.N_98_mux_4_cascade_ ));
    CascadeMux I__3048 (
            .O(N__15273),
            .I(\Lab_UT.dictrl.N_1304_0_0_cascade_ ));
    InMux I__3047 (
            .O(N__15270),
            .I(N__15267));
    LocalMux I__3046 (
            .O(N__15267),
            .I(N__15264));
    Span4Mux_v I__3045 (
            .O(N__15264),
            .I(N__15261));
    Odrv4 I__3044 (
            .O(N__15261),
            .I(\Lab_UT.dictrl.N_88_0_0 ));
    CascadeMux I__3043 (
            .O(N__15258),
            .I(\Lab_UT.dictrl.g1_1_1_cascade_ ));
    InMux I__3042 (
            .O(N__15255),
            .I(N__15252));
    LocalMux I__3041 (
            .O(N__15252),
            .I(\Lab_UT.dictrl.g1_0 ));
    CascadeMux I__3040 (
            .O(N__15249),
            .I(\Lab_UT.dictrl.N_116_mux_0_cascade_ ));
    InMux I__3039 (
            .O(N__15246),
            .I(N__15243));
    LocalMux I__3038 (
            .O(N__15243),
            .I(\Lab_UT.dictrl.N_116_mux_0_0_0 ));
    CascadeMux I__3037 (
            .O(N__15240),
            .I(\Lab_UT.dictrl.N_1304_0_1_0_cascade_ ));
    InMux I__3036 (
            .O(N__15237),
            .I(N__15234));
    LocalMux I__3035 (
            .O(N__15234),
            .I(\Lab_UT.dictrl.N_1304_0 ));
    CascadeMux I__3034 (
            .O(N__15231),
            .I(\Lab_UT.didp.countrce4.q_5_0_cascade_ ));
    InMux I__3033 (
            .O(N__15228),
            .I(N__15222));
    InMux I__3032 (
            .O(N__15227),
            .I(N__15219));
    CascadeMux I__3031 (
            .O(N__15226),
            .I(N__15216));
    InMux I__3030 (
            .O(N__15225),
            .I(N__15211));
    LocalMux I__3029 (
            .O(N__15222),
            .I(N__15206));
    LocalMux I__3028 (
            .O(N__15219),
            .I(N__15206));
    InMux I__3027 (
            .O(N__15216),
            .I(N__15199));
    InMux I__3026 (
            .O(N__15215),
            .I(N__15199));
    InMux I__3025 (
            .O(N__15214),
            .I(N__15199));
    LocalMux I__3024 (
            .O(N__15211),
            .I(N__15196));
    Span4Mux_s1_v I__3023 (
            .O(N__15206),
            .I(N__15193));
    LocalMux I__3022 (
            .O(N__15199),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    Odrv4 I__3021 (
            .O(N__15196),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    Odrv4 I__3020 (
            .O(N__15193),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    CascadeMux I__3019 (
            .O(N__15186),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__3018 (
            .O(N__15183),
            .I(N__15180));
    LocalMux I__3017 (
            .O(N__15180),
            .I(\Lab_UT.didp.countrce4.un20_qPone ));
    CascadeMux I__3016 (
            .O(N__15177),
            .I(\Lab_UT.didp.countrce4.q_5_3_cascade_ ));
    InMux I__3015 (
            .O(N__15174),
            .I(N__15166));
    InMux I__3014 (
            .O(N__15173),
            .I(N__15163));
    InMux I__3013 (
            .O(N__15172),
            .I(N__15154));
    InMux I__3012 (
            .O(N__15171),
            .I(N__15154));
    InMux I__3011 (
            .O(N__15170),
            .I(N__15154));
    InMux I__3010 (
            .O(N__15169),
            .I(N__15154));
    LocalMux I__3009 (
            .O(N__15166),
            .I(N__15147));
    LocalMux I__3008 (
            .O(N__15163),
            .I(N__15147));
    LocalMux I__3007 (
            .O(N__15154),
            .I(N__15147));
    Span4Mux_h I__3006 (
            .O(N__15147),
            .I(N__15144));
    Odrv4 I__3005 (
            .O(N__15144),
            .I(\Lab_UT.LdMtens ));
    InMux I__3004 (
            .O(N__15141),
            .I(N__15136));
    InMux I__3003 (
            .O(N__15140),
            .I(N__15131));
    InMux I__3002 (
            .O(N__15139),
            .I(N__15131));
    LocalMux I__3001 (
            .O(N__15136),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    LocalMux I__3000 (
            .O(N__15131),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    InMux I__2999 (
            .O(N__15126),
            .I(N__15123));
    LocalMux I__2998 (
            .O(N__15123),
            .I(N__15120));
    IoSpan4Mux I__2997 (
            .O(N__15120),
            .I(N__15117));
    Odrv4 I__2996 (
            .O(N__15117),
            .I(\Lab_UT.didp.did_alarmMatch_3 ));
    CascadeMux I__2995 (
            .O(N__15114),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_ ));
    InMux I__2994 (
            .O(N__15111),
            .I(N__15108));
    LocalMux I__2993 (
            .O(N__15108),
            .I(N__15105));
    Span4Mux_h I__2992 (
            .O(N__15105),
            .I(N__15102));
    Odrv4 I__2991 (
            .O(N__15102),
            .I(\Lab_UT.didp.did_alarmMatch_1 ));
    InMux I__2990 (
            .O(N__15099),
            .I(N__15096));
    LocalMux I__2989 (
            .O(N__15096),
            .I(N__15093));
    Odrv4 I__2988 (
            .O(N__15093),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_12 ));
    InMux I__2987 (
            .O(N__15090),
            .I(N__15086));
    CascadeMux I__2986 (
            .O(N__15089),
            .I(N__15083));
    LocalMux I__2985 (
            .O(N__15086),
            .I(N__15080));
    InMux I__2984 (
            .O(N__15083),
            .I(N__15075));
    Span12Mux_s6_h I__2983 (
            .O(N__15080),
            .I(N__15072));
    InMux I__2982 (
            .O(N__15079),
            .I(N__15067));
    InMux I__2981 (
            .O(N__15078),
            .I(N__15067));
    LocalMux I__2980 (
            .O(N__15075),
            .I(\Lab_UT.di_AMtens_3 ));
    Odrv12 I__2979 (
            .O(N__15072),
            .I(\Lab_UT.di_AMtens_3 ));
    LocalMux I__2978 (
            .O(N__15067),
            .I(\Lab_UT.di_AMtens_3 ));
    CascadeMux I__2977 (
            .O(N__15060),
            .I(N__15056));
    CascadeMux I__2976 (
            .O(N__15059),
            .I(N__15052));
    InMux I__2975 (
            .O(N__15056),
            .I(N__15039));
    InMux I__2974 (
            .O(N__15055),
            .I(N__15039));
    InMux I__2973 (
            .O(N__15052),
            .I(N__15039));
    InMux I__2972 (
            .O(N__15051),
            .I(N__15039));
    CascadeMux I__2971 (
            .O(N__15050),
            .I(N__15036));
    CascadeMux I__2970 (
            .O(N__15049),
            .I(N__15032));
    CascadeMux I__2969 (
            .O(N__15048),
            .I(N__15027));
    LocalMux I__2968 (
            .O(N__15039),
            .I(N__15018));
    InMux I__2967 (
            .O(N__15036),
            .I(N__15015));
    InMux I__2966 (
            .O(N__15035),
            .I(N__15010));
    InMux I__2965 (
            .O(N__15032),
            .I(N__15010));
    InMux I__2964 (
            .O(N__15031),
            .I(N__15003));
    InMux I__2963 (
            .O(N__15030),
            .I(N__15003));
    InMux I__2962 (
            .O(N__15027),
            .I(N__15003));
    InMux I__2961 (
            .O(N__15026),
            .I(N__14990));
    InMux I__2960 (
            .O(N__15025),
            .I(N__14990));
    InMux I__2959 (
            .O(N__15024),
            .I(N__14990));
    InMux I__2958 (
            .O(N__15023),
            .I(N__14990));
    InMux I__2957 (
            .O(N__15022),
            .I(N__14990));
    InMux I__2956 (
            .O(N__15021),
            .I(N__14990));
    Span4Mux_s2_v I__2955 (
            .O(N__15018),
            .I(N__14987));
    LocalMux I__2954 (
            .O(N__15015),
            .I(\Lab_UT.loadalarm_1 ));
    LocalMux I__2953 (
            .O(N__15010),
            .I(\Lab_UT.loadalarm_1 ));
    LocalMux I__2952 (
            .O(N__15003),
            .I(\Lab_UT.loadalarm_1 ));
    LocalMux I__2951 (
            .O(N__14990),
            .I(\Lab_UT.loadalarm_1 ));
    Odrv4 I__2950 (
            .O(N__14987),
            .I(\Lab_UT.loadalarm_1 ));
    InMux I__2949 (
            .O(N__14976),
            .I(N__14970));
    InMux I__2948 (
            .O(N__14975),
            .I(N__14963));
    InMux I__2947 (
            .O(N__14974),
            .I(N__14963));
    InMux I__2946 (
            .O(N__14973),
            .I(N__14963));
    LocalMux I__2945 (
            .O(N__14970),
            .I(N__14955));
    LocalMux I__2944 (
            .O(N__14963),
            .I(N__14955));
    CascadeMux I__2943 (
            .O(N__14962),
            .I(N__14945));
    InMux I__2942 (
            .O(N__14961),
            .I(N__14941));
    InMux I__2941 (
            .O(N__14960),
            .I(N__14938));
    Span4Mux_s2_v I__2940 (
            .O(N__14955),
            .I(N__14935));
    InMux I__2939 (
            .O(N__14954),
            .I(N__14930));
    InMux I__2938 (
            .O(N__14953),
            .I(N__14930));
    InMux I__2937 (
            .O(N__14952),
            .I(N__14917));
    InMux I__2936 (
            .O(N__14951),
            .I(N__14917));
    InMux I__2935 (
            .O(N__14950),
            .I(N__14917));
    InMux I__2934 (
            .O(N__14949),
            .I(N__14917));
    InMux I__2933 (
            .O(N__14948),
            .I(N__14917));
    InMux I__2932 (
            .O(N__14945),
            .I(N__14917));
    InMux I__2931 (
            .O(N__14944),
            .I(N__14914));
    LocalMux I__2930 (
            .O(N__14941),
            .I(\Lab_UT.loadalarm_0_0 ));
    LocalMux I__2929 (
            .O(N__14938),
            .I(\Lab_UT.loadalarm_0_0 ));
    Odrv4 I__2928 (
            .O(N__14935),
            .I(\Lab_UT.loadalarm_0_0 ));
    LocalMux I__2927 (
            .O(N__14930),
            .I(\Lab_UT.loadalarm_0_0 ));
    LocalMux I__2926 (
            .O(N__14917),
            .I(\Lab_UT.loadalarm_0_0 ));
    LocalMux I__2925 (
            .O(N__14914),
            .I(\Lab_UT.loadalarm_0_0 ));
    CascadeMux I__2924 (
            .O(N__14901),
            .I(N__14896));
    CascadeMux I__2923 (
            .O(N__14900),
            .I(N__14893));
    CascadeMux I__2922 (
            .O(N__14899),
            .I(N__14890));
    InMux I__2921 (
            .O(N__14896),
            .I(N__14876));
    InMux I__2920 (
            .O(N__14893),
            .I(N__14876));
    InMux I__2919 (
            .O(N__14890),
            .I(N__14876));
    InMux I__2918 (
            .O(N__14889),
            .I(N__14876));
    InMux I__2917 (
            .O(N__14888),
            .I(N__14876));
    CascadeMux I__2916 (
            .O(N__14887),
            .I(N__14872));
    LocalMux I__2915 (
            .O(N__14876),
            .I(N__14869));
    InMux I__2914 (
            .O(N__14875),
            .I(N__14864));
    InMux I__2913 (
            .O(N__14872),
            .I(N__14864));
    Span4Mux_v I__2912 (
            .O(N__14869),
            .I(N__14861));
    LocalMux I__2911 (
            .O(N__14864),
            .I(N__14858));
    Odrv4 I__2910 (
            .O(N__14861),
            .I(\Lab_UT.min1_3 ));
    Odrv12 I__2909 (
            .O(N__14858),
            .I(\Lab_UT.min1_3 ));
    InMux I__2908 (
            .O(N__14853),
            .I(N__14850));
    LocalMux I__2907 (
            .O(N__14850),
            .I(N__14847));
    Span4Mux_s0_v I__2906 (
            .O(N__14847),
            .I(N__14844));
    Odrv4 I__2905 (
            .O(N__14844),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__2904 (
            .O(N__14841),
            .I(N__14838));
    LocalMux I__2903 (
            .O(N__14838),
            .I(N__14835));
    Span4Mux_v I__2902 (
            .O(N__14835),
            .I(N__14830));
    InMux I__2901 (
            .O(N__14834),
            .I(N__14826));
    InMux I__2900 (
            .O(N__14833),
            .I(N__14823));
    Span4Mux_h I__2899 (
            .O(N__14830),
            .I(N__14820));
    InMux I__2898 (
            .O(N__14829),
            .I(N__14817));
    LocalMux I__2897 (
            .O(N__14826),
            .I(N__14814));
    LocalMux I__2896 (
            .O(N__14823),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__2895 (
            .O(N__14820),
            .I(\Lab_UT.di_AMtens_0 ));
    LocalMux I__2894 (
            .O(N__14817),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__2893 (
            .O(N__14814),
            .I(\Lab_UT.di_AMtens_0 ));
    InMux I__2892 (
            .O(N__14805),
            .I(N__14802));
    LocalMux I__2891 (
            .O(N__14802),
            .I(N__14799));
    Span4Mux_v I__2890 (
            .O(N__14799),
            .I(N__14795));
    InMux I__2889 (
            .O(N__14798),
            .I(N__14790));
    Span4Mux_h I__2888 (
            .O(N__14795),
            .I(N__14787));
    InMux I__2887 (
            .O(N__14794),
            .I(N__14784));
    InMux I__2886 (
            .O(N__14793),
            .I(N__14781));
    LocalMux I__2885 (
            .O(N__14790),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv4 I__2884 (
            .O(N__14787),
            .I(\Lab_UT.di_AMtens_1 ));
    LocalMux I__2883 (
            .O(N__14784),
            .I(\Lab_UT.di_AMtens_1 ));
    LocalMux I__2882 (
            .O(N__14781),
            .I(\Lab_UT.di_AMtens_1 ));
    CascadeMux I__2881 (
            .O(N__14772),
            .I(N__14767));
    InMux I__2880 (
            .O(N__14771),
            .I(N__14760));
    InMux I__2879 (
            .O(N__14770),
            .I(N__14757));
    InMux I__2878 (
            .O(N__14767),
            .I(N__14754));
    InMux I__2877 (
            .O(N__14766),
            .I(N__14745));
    InMux I__2876 (
            .O(N__14765),
            .I(N__14745));
    InMux I__2875 (
            .O(N__14764),
            .I(N__14745));
    InMux I__2874 (
            .O(N__14763),
            .I(N__14745));
    LocalMux I__2873 (
            .O(N__14760),
            .I(N__14740));
    LocalMux I__2872 (
            .O(N__14757),
            .I(N__14740));
    LocalMux I__2871 (
            .O(N__14754),
            .I(\Lab_UT.dicRun_2 ));
    LocalMux I__2870 (
            .O(N__14745),
            .I(\Lab_UT.dicRun_2 ));
    Odrv4 I__2869 (
            .O(N__14740),
            .I(\Lab_UT.dicRun_2 ));
    CascadeMux I__2868 (
            .O(N__14733),
            .I(N__14729));
    InMux I__2867 (
            .O(N__14732),
            .I(N__14726));
    InMux I__2866 (
            .O(N__14729),
            .I(N__14723));
    LocalMux I__2865 (
            .O(N__14726),
            .I(N__14719));
    LocalMux I__2864 (
            .O(N__14723),
            .I(N__14716));
    InMux I__2863 (
            .O(N__14722),
            .I(N__14712));
    Span4Mux_v I__2862 (
            .O(N__14719),
            .I(N__14709));
    Span4Mux_h I__2861 (
            .O(N__14716),
            .I(N__14706));
    InMux I__2860 (
            .O(N__14715),
            .I(N__14703));
    LocalMux I__2859 (
            .O(N__14712),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__2858 (
            .O(N__14709),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__2857 (
            .O(N__14706),
            .I(\Lab_UT.di_AMtens_2 ));
    LocalMux I__2856 (
            .O(N__14703),
            .I(\Lab_UT.di_AMtens_2 ));
    CascadeMux I__2855 (
            .O(N__14694),
            .I(N__14691));
    InMux I__2854 (
            .O(N__14691),
            .I(N__14685));
    InMux I__2853 (
            .O(N__14690),
            .I(N__14685));
    LocalMux I__2852 (
            .O(N__14685),
            .I(\Lab_UT.didp.countrce4.un13_qPone ));
    InMux I__2851 (
            .O(N__14682),
            .I(N__14678));
    CascadeMux I__2850 (
            .O(N__14681),
            .I(N__14675));
    LocalMux I__2849 (
            .O(N__14678),
            .I(N__14672));
    InMux I__2848 (
            .O(N__14675),
            .I(N__14668));
    Span4Mux_v I__2847 (
            .O(N__14672),
            .I(N__14665));
    CascadeMux I__2846 (
            .O(N__14671),
            .I(N__14661));
    LocalMux I__2845 (
            .O(N__14668),
            .I(N__14656));
    Span4Mux_v I__2844 (
            .O(N__14665),
            .I(N__14656));
    InMux I__2843 (
            .O(N__14664),
            .I(N__14653));
    InMux I__2842 (
            .O(N__14661),
            .I(N__14650));
    Odrv4 I__2841 (
            .O(N__14656),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__2840 (
            .O(N__14653),
            .I(\Lab_UT.di_AStens_0 ));
    LocalMux I__2839 (
            .O(N__14650),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__2838 (
            .O(N__14643),
            .I(N__14640));
    LocalMux I__2837 (
            .O(N__14640),
            .I(N__14637));
    Span4Mux_v I__2836 (
            .O(N__14637),
            .I(N__14632));
    InMux I__2835 (
            .O(N__14636),
            .I(N__14627));
    InMux I__2834 (
            .O(N__14635),
            .I(N__14627));
    Span4Mux_v I__2833 (
            .O(N__14632),
            .I(N__14623));
    LocalMux I__2832 (
            .O(N__14627),
            .I(N__14620));
    InMux I__2831 (
            .O(N__14626),
            .I(N__14617));
    Span4Mux_v I__2830 (
            .O(N__14623),
            .I(N__14612));
    Span4Mux_s2_v I__2829 (
            .O(N__14620),
            .I(N__14612));
    LocalMux I__2828 (
            .O(N__14617),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv4 I__2827 (
            .O(N__14612),
            .I(\Lab_UT.di_AStens_3 ));
    InMux I__2826 (
            .O(N__14607),
            .I(N__14604));
    LocalMux I__2825 (
            .O(N__14604),
            .I(N__14600));
    CascadeMux I__2824 (
            .O(N__14603),
            .I(N__14597));
    Span4Mux_v I__2823 (
            .O(N__14600),
            .I(N__14594));
    InMux I__2822 (
            .O(N__14597),
            .I(N__14591));
    Span4Mux_v I__2821 (
            .O(N__14594),
            .I(N__14585));
    LocalMux I__2820 (
            .O(N__14591),
            .I(N__14585));
    InMux I__2819 (
            .O(N__14590),
            .I(N__14581));
    Span4Mux_s2_v I__2818 (
            .O(N__14585),
            .I(N__14578));
    InMux I__2817 (
            .O(N__14584),
            .I(N__14575));
    LocalMux I__2816 (
            .O(N__14581),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__2815 (
            .O(N__14578),
            .I(\Lab_UT.di_AMones_1 ));
    LocalMux I__2814 (
            .O(N__14575),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__2813 (
            .O(N__14568),
            .I(N__14557));
    InMux I__2812 (
            .O(N__14567),
            .I(N__14557));
    InMux I__2811 (
            .O(N__14566),
            .I(N__14546));
    InMux I__2810 (
            .O(N__14565),
            .I(N__14546));
    InMux I__2809 (
            .O(N__14564),
            .I(N__14546));
    InMux I__2808 (
            .O(N__14563),
            .I(N__14546));
    InMux I__2807 (
            .O(N__14562),
            .I(N__14546));
    LocalMux I__2806 (
            .O(N__14557),
            .I(N__14543));
    LocalMux I__2805 (
            .O(N__14546),
            .I(\Lab_UT.min1_0 ));
    Odrv12 I__2804 (
            .O(N__14543),
            .I(\Lab_UT.min1_0 ));
    InMux I__2803 (
            .O(N__14538),
            .I(N__14527));
    InMux I__2802 (
            .O(N__14537),
            .I(N__14527));
    InMux I__2801 (
            .O(N__14536),
            .I(N__14516));
    InMux I__2800 (
            .O(N__14535),
            .I(N__14516));
    InMux I__2799 (
            .O(N__14534),
            .I(N__14516));
    InMux I__2798 (
            .O(N__14533),
            .I(N__14516));
    InMux I__2797 (
            .O(N__14532),
            .I(N__14516));
    LocalMux I__2796 (
            .O(N__14527),
            .I(N__14513));
    LocalMux I__2795 (
            .O(N__14516),
            .I(\Lab_UT.min1_1 ));
    Odrv4 I__2794 (
            .O(N__14513),
            .I(\Lab_UT.min1_1 ));
    CascadeMux I__2793 (
            .O(N__14508),
            .I(N__14504));
    InMux I__2792 (
            .O(N__14507),
            .I(N__14500));
    InMux I__2791 (
            .O(N__14504),
            .I(N__14497));
    InMux I__2790 (
            .O(N__14503),
            .I(N__14494));
    LocalMux I__2789 (
            .O(N__14500),
            .I(N__14490));
    LocalMux I__2788 (
            .O(N__14497),
            .I(N__14487));
    LocalMux I__2787 (
            .O(N__14494),
            .I(N__14484));
    InMux I__2786 (
            .O(N__14493),
            .I(N__14481));
    Span12Mux_s5_h I__2785 (
            .O(N__14490),
            .I(N__14478));
    Span12Mux_s6_v I__2784 (
            .O(N__14487),
            .I(N__14475));
    Span4Mux_v I__2783 (
            .O(N__14484),
            .I(N__14472));
    LocalMux I__2782 (
            .O(N__14481),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv12 I__2781 (
            .O(N__14478),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv12 I__2780 (
            .O(N__14475),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__2779 (
            .O(N__14472),
            .I(\Lab_UT.di_AMones_3 ));
    CascadeMux I__2778 (
            .O(N__14463),
            .I(\Lab_UT.didp.countrce1.q_5_1_cascade_ ));
    CascadeMux I__2777 (
            .O(N__14460),
            .I(N__14456));
    CascadeMux I__2776 (
            .O(N__14459),
            .I(N__14453));
    InMux I__2775 (
            .O(N__14456),
            .I(N__14448));
    InMux I__2774 (
            .O(N__14453),
            .I(N__14448));
    LocalMux I__2773 (
            .O(N__14448),
            .I(\Lab_UT.didp.countrce1.un13_qPone ));
    InMux I__2772 (
            .O(N__14445),
            .I(N__14438));
    InMux I__2771 (
            .O(N__14444),
            .I(N__14438));
    InMux I__2770 (
            .O(N__14443),
            .I(N__14435));
    LocalMux I__2769 (
            .O(N__14438),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    LocalMux I__2768 (
            .O(N__14435),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    CascadeMux I__2767 (
            .O(N__14430),
            .I(\Lab_UT.didp.un1_dicLdSones_0_cascade_ ));
    InMux I__2766 (
            .O(N__14427),
            .I(N__14424));
    LocalMux I__2765 (
            .O(N__14424),
            .I(N__14419));
    InMux I__2764 (
            .O(N__14423),
            .I(N__14416));
    CascadeMux I__2763 (
            .O(N__14422),
            .I(N__14410));
    Span4Mux_s2_v I__2762 (
            .O(N__14419),
            .I(N__14407));
    LocalMux I__2761 (
            .O(N__14416),
            .I(N__14404));
    InMux I__2760 (
            .O(N__14415),
            .I(N__14395));
    InMux I__2759 (
            .O(N__14414),
            .I(N__14395));
    InMux I__2758 (
            .O(N__14413),
            .I(N__14395));
    InMux I__2757 (
            .O(N__14410),
            .I(N__14395));
    Odrv4 I__2756 (
            .O(N__14407),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    Odrv12 I__2755 (
            .O(N__14404),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    LocalMux I__2754 (
            .O(N__14395),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    CascadeMux I__2753 (
            .O(N__14388),
            .I(N__14384));
    CascadeMux I__2752 (
            .O(N__14387),
            .I(N__14380));
    InMux I__2751 (
            .O(N__14384),
            .I(N__14376));
    InMux I__2750 (
            .O(N__14383),
            .I(N__14373));
    InMux I__2749 (
            .O(N__14380),
            .I(N__14370));
    InMux I__2748 (
            .O(N__14379),
            .I(N__14367));
    LocalMux I__2747 (
            .O(N__14376),
            .I(N__14364));
    LocalMux I__2746 (
            .O(N__14373),
            .I(N__14361));
    LocalMux I__2745 (
            .O(N__14370),
            .I(N__14356));
    LocalMux I__2744 (
            .O(N__14367),
            .I(N__14356));
    Span4Mux_s3_v I__2743 (
            .O(N__14364),
            .I(N__14353));
    Span4Mux_s3_v I__2742 (
            .O(N__14361),
            .I(N__14350));
    Odrv4 I__2741 (
            .O(N__14356),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__2740 (
            .O(N__14353),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__2739 (
            .O(N__14350),
            .I(\Lab_UT.di_AMones_2 ));
    InMux I__2738 (
            .O(N__14343),
            .I(N__14340));
    LocalMux I__2737 (
            .O(N__14340),
            .I(N__14337));
    Span4Mux_v I__2736 (
            .O(N__14337),
            .I(N__14334));
    Odrv4 I__2735 (
            .O(N__14334),
            .I(\Lab_UT.didp.did_alarmMatch_5 ));
    CascadeMux I__2734 (
            .O(N__14331),
            .I(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ));
    InMux I__2733 (
            .O(N__14328),
            .I(N__14325));
    LocalMux I__2732 (
            .O(N__14325),
            .I(N__14322));
    Odrv4 I__2731 (
            .O(N__14322),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    InMux I__2730 (
            .O(N__14319),
            .I(N__14316));
    LocalMux I__2729 (
            .O(N__14316),
            .I(bu_rx_data_i_4_fast_3));
    CascadeMux I__2728 (
            .O(N__14313),
            .I(N__14309));
    CascadeMux I__2727 (
            .O(N__14312),
            .I(N__14306));
    InMux I__2726 (
            .O(N__14309),
            .I(N__14303));
    InMux I__2725 (
            .O(N__14306),
            .I(N__14300));
    LocalMux I__2724 (
            .O(N__14303),
            .I(buart__rx_shifter_ret_5_fast));
    LocalMux I__2723 (
            .O(N__14300),
            .I(buart__rx_shifter_ret_5_fast));
    CascadeMux I__2722 (
            .O(N__14295),
            .I(\Lab_UT.dictrl.g1_1Z0Z_4_cascade_ ));
    CascadeMux I__2721 (
            .O(N__14292),
            .I(N__14289));
    InMux I__2720 (
            .O(N__14289),
            .I(N__14286));
    LocalMux I__2719 (
            .O(N__14286),
            .I(\Lab_UT.dictrl.N_98_mux_1 ));
    InMux I__2718 (
            .O(N__14283),
            .I(N__14280));
    LocalMux I__2717 (
            .O(N__14280),
            .I(\Lab_UT.dictrl.N_98_mux_0_0 ));
    CascadeMux I__2716 (
            .O(N__14277),
            .I(\Lab_UT.dictrl.g0_3_1_cascade_ ));
    CascadeMux I__2715 (
            .O(N__14274),
            .I(N__14268));
    InMux I__2714 (
            .O(N__14273),
            .I(N__14259));
    InMux I__2713 (
            .O(N__14272),
            .I(N__14259));
    InMux I__2712 (
            .O(N__14271),
            .I(N__14259));
    InMux I__2711 (
            .O(N__14268),
            .I(N__14259));
    LocalMux I__2710 (
            .O(N__14259),
            .I(bu_rx_data_7));
    InMux I__2709 (
            .O(N__14256),
            .I(N__14253));
    LocalMux I__2708 (
            .O(N__14253),
            .I(N__14250));
    Odrv12 I__2707 (
            .O(N__14250),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_6 ));
    CascadeMux I__2706 (
            .O(N__14247),
            .I(N__14244));
    InMux I__2705 (
            .O(N__14244),
            .I(N__14241));
    LocalMux I__2704 (
            .O(N__14241),
            .I(N__14238));
    Odrv4 I__2703 (
            .O(N__14238),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_7 ));
    CascadeMux I__2702 (
            .O(N__14235),
            .I(\Lab_UT.dictrl.N_127_0_0_cascade_ ));
    InMux I__2701 (
            .O(N__14232),
            .I(N__14226));
    InMux I__2700 (
            .O(N__14231),
            .I(N__14226));
    LocalMux I__2699 (
            .O(N__14226),
            .I(\Lab_UT.dictrl.justentered_0 ));
    CascadeMux I__2698 (
            .O(N__14223),
            .I(N__14215));
    InMux I__2697 (
            .O(N__14222),
            .I(N__14211));
    InMux I__2696 (
            .O(N__14221),
            .I(N__14208));
    InMux I__2695 (
            .O(N__14220),
            .I(N__14197));
    InMux I__2694 (
            .O(N__14219),
            .I(N__14197));
    InMux I__2693 (
            .O(N__14218),
            .I(N__14197));
    InMux I__2692 (
            .O(N__14215),
            .I(N__14197));
    InMux I__2691 (
            .O(N__14214),
            .I(N__14197));
    LocalMux I__2690 (
            .O(N__14211),
            .I(\Lab_UT.shifter_ret_3_RNIK5FS8_0 ));
    LocalMux I__2689 (
            .O(N__14208),
            .I(\Lab_UT.shifter_ret_3_RNIK5FS8_0 ));
    LocalMux I__2688 (
            .O(N__14197),
            .I(\Lab_UT.shifter_ret_3_RNIK5FS8_0 ));
    InMux I__2687 (
            .O(N__14190),
            .I(N__14181));
    InMux I__2686 (
            .O(N__14189),
            .I(N__14178));
    InMux I__2685 (
            .O(N__14188),
            .I(N__14167));
    InMux I__2684 (
            .O(N__14187),
            .I(N__14167));
    InMux I__2683 (
            .O(N__14186),
            .I(N__14167));
    InMux I__2682 (
            .O(N__14185),
            .I(N__14167));
    InMux I__2681 (
            .O(N__14184),
            .I(N__14167));
    LocalMux I__2680 (
            .O(N__14181),
            .I(\Lab_UT.shifter_ret_3_RNIQBH29_0 ));
    LocalMux I__2679 (
            .O(N__14178),
            .I(\Lab_UT.shifter_ret_3_RNIQBH29_0 ));
    LocalMux I__2678 (
            .O(N__14167),
            .I(\Lab_UT.shifter_ret_3_RNIQBH29_0 ));
    InMux I__2677 (
            .O(N__14160),
            .I(N__14154));
    InMux I__2676 (
            .O(N__14159),
            .I(N__14154));
    LocalMux I__2675 (
            .O(N__14154),
            .I(\Lab_UT.armed ));
    CascadeMux I__2674 (
            .O(N__14151),
            .I(\Lab_UT.armed_cascade_ ));
    InMux I__2673 (
            .O(N__14148),
            .I(N__14141));
    InMux I__2672 (
            .O(N__14147),
            .I(N__14141));
    InMux I__2671 (
            .O(N__14146),
            .I(N__14138));
    LocalMux I__2670 (
            .O(N__14141),
            .I(N__14135));
    LocalMux I__2669 (
            .O(N__14138),
            .I(N__14132));
    Odrv4 I__2668 (
            .O(N__14135),
            .I(\Lab_UT.alarmMatch ));
    Odrv12 I__2667 (
            .O(N__14132),
            .I(\Lab_UT.alarmMatch ));
    InMux I__2666 (
            .O(N__14127),
            .I(N__14124));
    LocalMux I__2665 (
            .O(N__14124),
            .I(G_203));
    InMux I__2664 (
            .O(N__14121),
            .I(N__14118));
    LocalMux I__2663 (
            .O(N__14118),
            .I(\Lab_UT.dictrl.alarmstate8_2_reti ));
    CascadeMux I__2662 (
            .O(N__14115),
            .I(\Lab_UT.dictrl.alarmstate8_10_3_cascade_ ));
    InMux I__2661 (
            .O(N__14112),
            .I(N__14109));
    LocalMux I__2660 (
            .O(N__14109),
            .I(N__14105));
    InMux I__2659 (
            .O(N__14108),
            .I(N__14102));
    Odrv4 I__2658 (
            .O(N__14105),
            .I(\Lab_UT.dictrl.alarmstate8 ));
    LocalMux I__2657 (
            .O(N__14102),
            .I(\Lab_UT.dictrl.alarmstate8 ));
    CascadeMux I__2656 (
            .O(N__14097),
            .I(\Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_ ));
    CascadeMux I__2655 (
            .O(N__14094),
            .I(\Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_ ));
    InMux I__2654 (
            .O(N__14091),
            .I(N__14088));
    LocalMux I__2653 (
            .O(N__14088),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i ));
    InMux I__2652 (
            .O(N__14085),
            .I(N__14079));
    InMux I__2651 (
            .O(N__14084),
            .I(N__14079));
    LocalMux I__2650 (
            .O(N__14079),
            .I(\Lab_UT.dictrl.alarmstate_0_sqmuxa_1 ));
    CascadeMux I__2649 (
            .O(N__14076),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_ ));
    InMux I__2648 (
            .O(N__14073),
            .I(N__14070));
    LocalMux I__2647 (
            .O(N__14070),
            .I(\Lab_UT.dictrl.alarmstate_1_0_i_0 ));
    CascadeMux I__2646 (
            .O(N__14067),
            .I(\Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_ ));
    InMux I__2645 (
            .O(N__14064),
            .I(N__14061));
    LocalMux I__2644 (
            .O(N__14061),
            .I(\Lab_UT.dictrl.g0_0_0_a3_0_0 ));
    CascadeMux I__2643 (
            .O(N__14058),
            .I(N__14055));
    InMux I__2642 (
            .O(N__14055),
            .I(N__14052));
    LocalMux I__2641 (
            .O(N__14052),
            .I(\Lab_UT.dictrl.N_127_0_0 ));
    InMux I__2640 (
            .O(N__14049),
            .I(N__14044));
    InMux I__2639 (
            .O(N__14048),
            .I(N__14039));
    InMux I__2638 (
            .O(N__14047),
            .I(N__14039));
    LocalMux I__2637 (
            .O(N__14044),
            .I(\Lab_UT.trig ));
    LocalMux I__2636 (
            .O(N__14039),
            .I(\Lab_UT.trig ));
    InMux I__2635 (
            .O(N__14034),
            .I(N__14030));
    InMux I__2634 (
            .O(N__14033),
            .I(N__14027));
    LocalMux I__2633 (
            .O(N__14030),
            .I(N__14024));
    LocalMux I__2632 (
            .O(N__14027),
            .I(N__14019));
    Span4Mux_s2_v I__2631 (
            .O(N__14024),
            .I(N__14016));
    InMux I__2630 (
            .O(N__14023),
            .I(N__14013));
    InMux I__2629 (
            .O(N__14022),
            .I(N__14010));
    Span4Mux_v I__2628 (
            .O(N__14019),
            .I(N__14005));
    Span4Mux_v I__2627 (
            .O(N__14016),
            .I(N__14005));
    LocalMux I__2626 (
            .O(N__14013),
            .I(N__14002));
    LocalMux I__2625 (
            .O(N__14010),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__2624 (
            .O(N__14005),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv12 I__2623 (
            .O(N__14002),
            .I(\Lab_UT.di_ASones_1 ));
    CascadeMux I__2622 (
            .O(N__13995),
            .I(N__13992));
    InMux I__2621 (
            .O(N__13992),
            .I(N__13988));
    InMux I__2620 (
            .O(N__13991),
            .I(N__13983));
    LocalMux I__2619 (
            .O(N__13988),
            .I(N__13980));
    CascadeMux I__2618 (
            .O(N__13987),
            .I(N__13977));
    CascadeMux I__2617 (
            .O(N__13986),
            .I(N__13974));
    LocalMux I__2616 (
            .O(N__13983),
            .I(N__13971));
    Span4Mux_s2_v I__2615 (
            .O(N__13980),
            .I(N__13968));
    InMux I__2614 (
            .O(N__13977),
            .I(N__13965));
    InMux I__2613 (
            .O(N__13974),
            .I(N__13962));
    Span4Mux_v I__2612 (
            .O(N__13971),
            .I(N__13957));
    Span4Mux_v I__2611 (
            .O(N__13968),
            .I(N__13957));
    LocalMux I__2610 (
            .O(N__13965),
            .I(N__13954));
    LocalMux I__2609 (
            .O(N__13962),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__2608 (
            .O(N__13957),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv12 I__2607 (
            .O(N__13954),
            .I(\Lab_UT.di_ASones_2 ));
    InMux I__2606 (
            .O(N__13947),
            .I(N__13942));
    InMux I__2605 (
            .O(N__13946),
            .I(N__13937));
    InMux I__2604 (
            .O(N__13945),
            .I(N__13937));
    LocalMux I__2603 (
            .O(N__13942),
            .I(N__13933));
    LocalMux I__2602 (
            .O(N__13937),
            .I(N__13930));
    InMux I__2601 (
            .O(N__13936),
            .I(N__13927));
    Span4Mux_v I__2600 (
            .O(N__13933),
            .I(N__13922));
    Span4Mux_s2_v I__2599 (
            .O(N__13930),
            .I(N__13922));
    LocalMux I__2598 (
            .O(N__13927),
            .I(N__13917));
    Span4Mux_v I__2597 (
            .O(N__13922),
            .I(N__13917));
    Odrv4 I__2596 (
            .O(N__13917),
            .I(\Lab_UT.di_ASones_3 ));
    CascadeMux I__2595 (
            .O(N__13914),
            .I(N__13908));
    InMux I__2594 (
            .O(N__13913),
            .I(N__13905));
    InMux I__2593 (
            .O(N__13912),
            .I(N__13902));
    InMux I__2592 (
            .O(N__13911),
            .I(N__13899));
    InMux I__2591 (
            .O(N__13908),
            .I(N__13896));
    LocalMux I__2590 (
            .O(N__13905),
            .I(N__13893));
    LocalMux I__2589 (
            .O(N__13902),
            .I(N__13888));
    LocalMux I__2588 (
            .O(N__13899),
            .I(N__13888));
    LocalMux I__2587 (
            .O(N__13896),
            .I(N__13885));
    Span4Mux_h I__2586 (
            .O(N__13893),
            .I(N__13882));
    Span4Mux_s2_v I__2585 (
            .O(N__13888),
            .I(N__13879));
    Odrv4 I__2584 (
            .O(N__13885),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__2583 (
            .O(N__13882),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__2582 (
            .O(N__13879),
            .I(\Lab_UT.di_AMones_0 ));
    CascadeMux I__2581 (
            .O(N__13872),
            .I(N__13867));
    CascadeMux I__2580 (
            .O(N__13871),
            .I(N__13864));
    CascadeMux I__2579 (
            .O(N__13870),
            .I(N__13858));
    InMux I__2578 (
            .O(N__13867),
            .I(N__13846));
    InMux I__2577 (
            .O(N__13864),
            .I(N__13846));
    InMux I__2576 (
            .O(N__13863),
            .I(N__13846));
    InMux I__2575 (
            .O(N__13862),
            .I(N__13846));
    InMux I__2574 (
            .O(N__13861),
            .I(N__13846));
    InMux I__2573 (
            .O(N__13858),
            .I(N__13841));
    InMux I__2572 (
            .O(N__13857),
            .I(N__13841));
    LocalMux I__2571 (
            .O(N__13846),
            .I(N__13838));
    LocalMux I__2570 (
            .O(N__13841),
            .I(\Lab_UT.min1_2 ));
    Odrv4 I__2569 (
            .O(N__13838),
            .I(\Lab_UT.min1_2 ));
    InMux I__2568 (
            .O(N__13833),
            .I(N__13830));
    LocalMux I__2567 (
            .O(N__13830),
            .I(\uu2.bitmapZ0Z_34 ));
    InMux I__2566 (
            .O(N__13827),
            .I(N__13824));
    LocalMux I__2565 (
            .O(N__13824),
            .I(N__13820));
    InMux I__2564 (
            .O(N__13823),
            .I(N__13806));
    Span4Mux_h I__2563 (
            .O(N__13820),
            .I(N__13801));
    InMux I__2562 (
            .O(N__13819),
            .I(N__13798));
    InMux I__2561 (
            .O(N__13818),
            .I(N__13791));
    InMux I__2560 (
            .O(N__13817),
            .I(N__13791));
    InMux I__2559 (
            .O(N__13816),
            .I(N__13791));
    InMux I__2558 (
            .O(N__13815),
            .I(N__13784));
    InMux I__2557 (
            .O(N__13814),
            .I(N__13784));
    InMux I__2556 (
            .O(N__13813),
            .I(N__13784));
    InMux I__2555 (
            .O(N__13812),
            .I(N__13775));
    InMux I__2554 (
            .O(N__13811),
            .I(N__13775));
    InMux I__2553 (
            .O(N__13810),
            .I(N__13775));
    InMux I__2552 (
            .O(N__13809),
            .I(N__13775));
    LocalMux I__2551 (
            .O(N__13806),
            .I(N__13772));
    InMux I__2550 (
            .O(N__13805),
            .I(N__13769));
    InMux I__2549 (
            .O(N__13804),
            .I(N__13766));
    Odrv4 I__2548 (
            .O(N__13801),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2547 (
            .O(N__13798),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2546 (
            .O(N__13791),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2545 (
            .O(N__13784),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2544 (
            .O(N__13775),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv12 I__2543 (
            .O(N__13772),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2542 (
            .O(N__13769),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2541 (
            .O(N__13766),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    CascadeMux I__2540 (
            .O(N__13749),
            .I(N__13746));
    InMux I__2539 (
            .O(N__13746),
            .I(N__13743));
    LocalMux I__2538 (
            .O(N__13743),
            .I(\uu2.bitmapZ0Z_290 ));
    InMux I__2537 (
            .O(N__13740),
            .I(N__13737));
    LocalMux I__2536 (
            .O(N__13737),
            .I(N__13734));
    Span4Mux_h I__2535 (
            .O(N__13734),
            .I(N__13731));
    Odrv4 I__2534 (
            .O(N__13731),
            .I(\uu2.bitmap_pmux_26_bm_1 ));
    InMux I__2533 (
            .O(N__13728),
            .I(N__13725));
    LocalMux I__2532 (
            .O(N__13725),
            .I(N__13722));
    Span4Mux_h I__2531 (
            .O(N__13722),
            .I(N__13717));
    InMux I__2530 (
            .O(N__13721),
            .I(N__13714));
    InMux I__2529 (
            .O(N__13720),
            .I(N__13711));
    Span4Mux_v I__2528 (
            .O(N__13717),
            .I(N__13693));
    LocalMux I__2527 (
            .O(N__13714),
            .I(N__13690));
    LocalMux I__2526 (
            .O(N__13711),
            .I(N__13687));
    InMux I__2525 (
            .O(N__13710),
            .I(N__13684));
    InMux I__2524 (
            .O(N__13709),
            .I(N__13677));
    InMux I__2523 (
            .O(N__13708),
            .I(N__13677));
    InMux I__2522 (
            .O(N__13707),
            .I(N__13677));
    InMux I__2521 (
            .O(N__13706),
            .I(N__13668));
    InMux I__2520 (
            .O(N__13705),
            .I(N__13668));
    InMux I__2519 (
            .O(N__13704),
            .I(N__13668));
    InMux I__2518 (
            .O(N__13703),
            .I(N__13668));
    InMux I__2517 (
            .O(N__13702),
            .I(N__13665));
    InMux I__2516 (
            .O(N__13701),
            .I(N__13662));
    InMux I__2515 (
            .O(N__13700),
            .I(N__13657));
    InMux I__2514 (
            .O(N__13699),
            .I(N__13657));
    InMux I__2513 (
            .O(N__13698),
            .I(N__13650));
    InMux I__2512 (
            .O(N__13697),
            .I(N__13650));
    InMux I__2511 (
            .O(N__13696),
            .I(N__13650));
    Odrv4 I__2510 (
            .O(N__13693),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv12 I__2509 (
            .O(N__13690),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__2508 (
            .O(N__13687),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2507 (
            .O(N__13684),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2506 (
            .O(N__13677),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2505 (
            .O(N__13668),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2504 (
            .O(N__13665),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2503 (
            .O(N__13662),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2502 (
            .O(N__13657),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__2501 (
            .O(N__13650),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__2500 (
            .O(N__13629),
            .I(N__13626));
    LocalMux I__2499 (
            .O(N__13626),
            .I(N__13623));
    Odrv4 I__2498 (
            .O(N__13623),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__2497 (
            .O(N__13620),
            .I(N__13617));
    LocalMux I__2496 (
            .O(N__13617),
            .I(\uu2.bitmapZ0Z_162 ));
    InMux I__2495 (
            .O(N__13614),
            .I(N__13611));
    LocalMux I__2494 (
            .O(N__13611),
            .I(N__13608));
    Odrv4 I__2493 (
            .O(N__13608),
            .I(\uu2.N_217 ));
    CascadeMux I__2492 (
            .O(N__13605),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ));
    InMux I__2491 (
            .O(N__13602),
            .I(N__13599));
    LocalMux I__2490 (
            .O(N__13599),
            .I(N__13596));
    Odrv12 I__2489 (
            .O(N__13596),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_11 ));
    CascadeMux I__2488 (
            .O(N__13593),
            .I(\Lab_UT.didp.countrce4.q_5_2_cascade_ ));
    CascadeMux I__2487 (
            .O(N__13590),
            .I(N__13584));
    InMux I__2486 (
            .O(N__13589),
            .I(N__13581));
    InMux I__2485 (
            .O(N__13588),
            .I(N__13578));
    InMux I__2484 (
            .O(N__13587),
            .I(N__13575));
    InMux I__2483 (
            .O(N__13584),
            .I(N__13572));
    LocalMux I__2482 (
            .O(N__13581),
            .I(N__13569));
    LocalMux I__2481 (
            .O(N__13578),
            .I(N__13564));
    LocalMux I__2480 (
            .O(N__13575),
            .I(N__13564));
    LocalMux I__2479 (
            .O(N__13572),
            .I(N__13559));
    Span4Mux_v I__2478 (
            .O(N__13569),
            .I(N__13559));
    Span4Mux_s2_v I__2477 (
            .O(N__13564),
            .I(N__13556));
    Odrv4 I__2476 (
            .O(N__13559),
            .I(\Lab_UT.di_ASones_0 ));
    Odrv4 I__2475 (
            .O(N__13556),
            .I(\Lab_UT.di_ASones_0 ));
    CascadeMux I__2474 (
            .O(N__13551),
            .I(\uu2.o_adder_vbuf_w_addr_displaying_6_cascade_ ));
    CEMux I__2473 (
            .O(N__13548),
            .I(N__13544));
    CEMux I__2472 (
            .O(N__13547),
            .I(N__13541));
    LocalMux I__2471 (
            .O(N__13544),
            .I(N__13538));
    LocalMux I__2470 (
            .O(N__13541),
            .I(N__13535));
    Span4Mux_v I__2469 (
            .O(N__13538),
            .I(N__13532));
    Span4Mux_v I__2468 (
            .O(N__13535),
            .I(N__13529));
    Span4Mux_h I__2467 (
            .O(N__13532),
            .I(N__13526));
    Odrv4 I__2466 (
            .O(N__13529),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    Odrv4 I__2465 (
            .O(N__13526),
            .I(\uu2.un21_w_addr_displaying_i_0 ));
    CascadeMux I__2464 (
            .O(N__13521),
            .I(N__13518));
    InMux I__2463 (
            .O(N__13518),
            .I(N__13515));
    LocalMux I__2462 (
            .O(N__13515),
            .I(N__13512));
    Span4Mux_v I__2461 (
            .O(N__13512),
            .I(N__13509));
    Odrv4 I__2460 (
            .O(N__13509),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    InMux I__2459 (
            .O(N__13506),
            .I(N__13503));
    LocalMux I__2458 (
            .O(N__13503),
            .I(N__13499));
    CascadeMux I__2457 (
            .O(N__13502),
            .I(N__13495));
    Span4Mux_v I__2456 (
            .O(N__13499),
            .I(N__13490));
    InMux I__2455 (
            .O(N__13498),
            .I(N__13487));
    InMux I__2454 (
            .O(N__13495),
            .I(N__13482));
    InMux I__2453 (
            .O(N__13494),
            .I(N__13482));
    CascadeMux I__2452 (
            .O(N__13493),
            .I(N__13479));
    Span4Mux_v I__2451 (
            .O(N__13490),
            .I(N__13468));
    LocalMux I__2450 (
            .O(N__13487),
            .I(N__13468));
    LocalMux I__2449 (
            .O(N__13482),
            .I(N__13468));
    InMux I__2448 (
            .O(N__13479),
            .I(N__13461));
    InMux I__2447 (
            .O(N__13478),
            .I(N__13461));
    InMux I__2446 (
            .O(N__13477),
            .I(N__13461));
    InMux I__2445 (
            .O(N__13476),
            .I(N__13458));
    InMux I__2444 (
            .O(N__13475),
            .I(N__13455));
    Span4Mux_h I__2443 (
            .O(N__13468),
            .I(N__13452));
    LocalMux I__2442 (
            .O(N__13461),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2441 (
            .O(N__13458),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2440 (
            .O(N__13455),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2439 (
            .O(N__13452),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__2438 (
            .O(N__13443),
            .I(N__13438));
    InMux I__2437 (
            .O(N__13442),
            .I(N__13435));
    InMux I__2436 (
            .O(N__13441),
            .I(N__13432));
    InMux I__2435 (
            .O(N__13438),
            .I(N__13428));
    LocalMux I__2434 (
            .O(N__13435),
            .I(N__13425));
    LocalMux I__2433 (
            .O(N__13432),
            .I(N__13421));
    CascadeMux I__2432 (
            .O(N__13431),
            .I(N__13417));
    LocalMux I__2431 (
            .O(N__13428),
            .I(N__13412));
    Span4Mux_h I__2430 (
            .O(N__13425),
            .I(N__13412));
    InMux I__2429 (
            .O(N__13424),
            .I(N__13409));
    Span4Mux_h I__2428 (
            .O(N__13421),
            .I(N__13406));
    InMux I__2427 (
            .O(N__13420),
            .I(N__13401));
    InMux I__2426 (
            .O(N__13417),
            .I(N__13401));
    Span4Mux_v I__2425 (
            .O(N__13412),
            .I(N__13398));
    LocalMux I__2424 (
            .O(N__13409),
            .I(\uu2.un15_w_data_displaying_6 ));
    Odrv4 I__2423 (
            .O(N__13406),
            .I(\uu2.un15_w_data_displaying_6 ));
    LocalMux I__2422 (
            .O(N__13401),
            .I(\uu2.un15_w_data_displaying_6 ));
    Odrv4 I__2421 (
            .O(N__13398),
            .I(\uu2.un15_w_data_displaying_6 ));
    InMux I__2420 (
            .O(N__13389),
            .I(N__13386));
    LocalMux I__2419 (
            .O(N__13386),
            .I(N__13381));
    InMux I__2418 (
            .O(N__13385),
            .I(N__13374));
    InMux I__2417 (
            .O(N__13384),
            .I(N__13371));
    Span4Mux_h I__2416 (
            .O(N__13381),
            .I(N__13368));
    InMux I__2415 (
            .O(N__13380),
            .I(N__13359));
    InMux I__2414 (
            .O(N__13379),
            .I(N__13359));
    InMux I__2413 (
            .O(N__13378),
            .I(N__13359));
    InMux I__2412 (
            .O(N__13377),
            .I(N__13359));
    LocalMux I__2411 (
            .O(N__13374),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2410 (
            .O(N__13371),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__2409 (
            .O(N__13368),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2408 (
            .O(N__13359),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__2407 (
            .O(N__13350),
            .I(N__13347));
    LocalMux I__2406 (
            .O(N__13347),
            .I(N__13343));
    CascadeMux I__2405 (
            .O(N__13346),
            .I(N__13339));
    Span4Mux_v I__2404 (
            .O(N__13343),
            .I(N__13333));
    InMux I__2403 (
            .O(N__13342),
            .I(N__13330));
    InMux I__2402 (
            .O(N__13339),
            .I(N__13327));
    InMux I__2401 (
            .O(N__13338),
            .I(N__13324));
    InMux I__2400 (
            .O(N__13337),
            .I(N__13314));
    InMux I__2399 (
            .O(N__13336),
            .I(N__13314));
    Span4Mux_h I__2398 (
            .O(N__13333),
            .I(N__13308));
    LocalMux I__2397 (
            .O(N__13330),
            .I(N__13301));
    LocalMux I__2396 (
            .O(N__13327),
            .I(N__13301));
    LocalMux I__2395 (
            .O(N__13324),
            .I(N__13301));
    InMux I__2394 (
            .O(N__13323),
            .I(N__13298));
    InMux I__2393 (
            .O(N__13322),
            .I(N__13295));
    InMux I__2392 (
            .O(N__13321),
            .I(N__13292));
    InMux I__2391 (
            .O(N__13320),
            .I(N__13287));
    InMux I__2390 (
            .O(N__13319),
            .I(N__13287));
    LocalMux I__2389 (
            .O(N__13314),
            .I(N__13284));
    InMux I__2388 (
            .O(N__13313),
            .I(N__13277));
    InMux I__2387 (
            .O(N__13312),
            .I(N__13277));
    InMux I__2386 (
            .O(N__13311),
            .I(N__13277));
    Odrv4 I__2385 (
            .O(N__13308),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2384 (
            .O(N__13301),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2383 (
            .O(N__13298),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2382 (
            .O(N__13295),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2381 (
            .O(N__13292),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2380 (
            .O(N__13287),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2379 (
            .O(N__13284),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2378 (
            .O(N__13277),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__2377 (
            .O(N__13260),
            .I(N__13257));
    LocalMux I__2376 (
            .O(N__13257),
            .I(N__13254));
    Span4Mux_h I__2375 (
            .O(N__13254),
            .I(N__13247));
    CascadeMux I__2374 (
            .O(N__13253),
            .I(N__13243));
    CascadeMux I__2373 (
            .O(N__13252),
            .I(N__13240));
    CascadeMux I__2372 (
            .O(N__13251),
            .I(N__13237));
    InMux I__2371 (
            .O(N__13250),
            .I(N__13234));
    Span4Mux_v I__2370 (
            .O(N__13247),
            .I(N__13231));
    InMux I__2369 (
            .O(N__13246),
            .I(N__13226));
    InMux I__2368 (
            .O(N__13243),
            .I(N__13226));
    InMux I__2367 (
            .O(N__13240),
            .I(N__13221));
    InMux I__2366 (
            .O(N__13237),
            .I(N__13221));
    LocalMux I__2365 (
            .O(N__13234),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    Odrv4 I__2364 (
            .O(N__13231),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2363 (
            .O(N__13226),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2362 (
            .O(N__13221),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__2361 (
            .O(N__13212),
            .I(N__13209));
    LocalMux I__2360 (
            .O(N__13209),
            .I(N__13206));
    Span4Mux_h I__2359 (
            .O(N__13206),
            .I(N__13203));
    Odrv4 I__2358 (
            .O(N__13203),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    InMux I__2357 (
            .O(N__13200),
            .I(N__13197));
    LocalMux I__2356 (
            .O(N__13197),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__2355 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__2354 (
            .O(N__13191),
            .I(\uu2.bitmap_pmux_25_am_1 ));
    CascadeMux I__2353 (
            .O(N__13188),
            .I(N__13185));
    InMux I__2352 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__2351 (
            .O(N__13182),
            .I(N__13179));
    Odrv4 I__2350 (
            .O(N__13179),
            .I(\uu2.bitmapZ0Z_194 ));
    CascadeMux I__2349 (
            .O(N__13176),
            .I(N__13173));
    InMux I__2348 (
            .O(N__13173),
            .I(N__13165));
    InMux I__2347 (
            .O(N__13172),
            .I(N__13162));
    InMux I__2346 (
            .O(N__13171),
            .I(N__13156));
    InMux I__2345 (
            .O(N__13170),
            .I(N__13152));
    InMux I__2344 (
            .O(N__13169),
            .I(N__13145));
    InMux I__2343 (
            .O(N__13168),
            .I(N__13145));
    LocalMux I__2342 (
            .O(N__13165),
            .I(N__13140));
    LocalMux I__2341 (
            .O(N__13162),
            .I(N__13140));
    InMux I__2340 (
            .O(N__13161),
            .I(N__13133));
    InMux I__2339 (
            .O(N__13160),
            .I(N__13133));
    InMux I__2338 (
            .O(N__13159),
            .I(N__13133));
    LocalMux I__2337 (
            .O(N__13156),
            .I(N__13130));
    InMux I__2336 (
            .O(N__13155),
            .I(N__13127));
    LocalMux I__2335 (
            .O(N__13152),
            .I(N__13124));
    CascadeMux I__2334 (
            .O(N__13151),
            .I(N__13121));
    InMux I__2333 (
            .O(N__13150),
            .I(N__13110));
    LocalMux I__2332 (
            .O(N__13145),
            .I(N__13101));
    Span4Mux_v I__2331 (
            .O(N__13140),
            .I(N__13101));
    LocalMux I__2330 (
            .O(N__13133),
            .I(N__13101));
    Span4Mux_h I__2329 (
            .O(N__13130),
            .I(N__13101));
    LocalMux I__2328 (
            .O(N__13127),
            .I(N__13096));
    Span4Mux_s0_v I__2327 (
            .O(N__13124),
            .I(N__13096));
    InMux I__2326 (
            .O(N__13121),
            .I(N__13093));
    InMux I__2325 (
            .O(N__13120),
            .I(N__13088));
    InMux I__2324 (
            .O(N__13119),
            .I(N__13088));
    InMux I__2323 (
            .O(N__13118),
            .I(N__13079));
    InMux I__2322 (
            .O(N__13117),
            .I(N__13079));
    InMux I__2321 (
            .O(N__13116),
            .I(N__13079));
    InMux I__2320 (
            .O(N__13115),
            .I(N__13079));
    InMux I__2319 (
            .O(N__13114),
            .I(N__13074));
    InMux I__2318 (
            .O(N__13113),
            .I(N__13074));
    LocalMux I__2317 (
            .O(N__13110),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2316 (
            .O(N__13101),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2315 (
            .O(N__13096),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2314 (
            .O(N__13093),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2313 (
            .O(N__13088),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2312 (
            .O(N__13079),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2311 (
            .O(N__13074),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__2310 (
            .O(N__13059),
            .I(N__13056));
    LocalMux I__2309 (
            .O(N__13056),
            .I(N__13053));
    Span4Mux_h I__2308 (
            .O(N__13053),
            .I(N__13050));
    Odrv4 I__2307 (
            .O(N__13050),
            .I(\uu2.bitmap_RNIV8902Z0Z_66 ));
    CascadeMux I__2306 (
            .O(N__13047),
            .I(\Lab_UT.didp.un2_did_alarmMatch_0_cascade_ ));
    InMux I__2305 (
            .O(N__13044),
            .I(N__13038));
    InMux I__2304 (
            .O(N__13043),
            .I(N__13038));
    LocalMux I__2303 (
            .O(N__13038),
            .I(N__13030));
    InMux I__2302 (
            .O(N__13037),
            .I(N__13019));
    InMux I__2301 (
            .O(N__13036),
            .I(N__13019));
    InMux I__2300 (
            .O(N__13035),
            .I(N__13019));
    InMux I__2299 (
            .O(N__13034),
            .I(N__13019));
    InMux I__2298 (
            .O(N__13033),
            .I(N__13019));
    Span4Mux_s2_v I__2297 (
            .O(N__13030),
            .I(N__13016));
    LocalMux I__2296 (
            .O(N__13019),
            .I(N__13013));
    Odrv4 I__2295 (
            .O(N__13016),
            .I(\Lab_UT.sec2_0 ));
    Odrv4 I__2294 (
            .O(N__13013),
            .I(\Lab_UT.sec2_0 ));
    CascadeMux I__2293 (
            .O(N__13008),
            .I(\Lab_UT.loadalarm_0_0_cascade_ ));
    InMux I__2292 (
            .O(N__13005),
            .I(N__12987));
    InMux I__2291 (
            .O(N__13004),
            .I(N__12987));
    InMux I__2290 (
            .O(N__13003),
            .I(N__12987));
    InMux I__2289 (
            .O(N__13002),
            .I(N__12987));
    InMux I__2288 (
            .O(N__13001),
            .I(N__12987));
    InMux I__2287 (
            .O(N__13000),
            .I(N__12987));
    LocalMux I__2286 (
            .O(N__12987),
            .I(N__12983));
    InMux I__2285 (
            .O(N__12986),
            .I(N__12980));
    Span4Mux_h I__2284 (
            .O(N__12983),
            .I(N__12977));
    LocalMux I__2283 (
            .O(N__12980),
            .I(N__12974));
    Odrv4 I__2282 (
            .O(N__12977),
            .I(\Lab_UT.sec1_0 ));
    Odrv4 I__2281 (
            .O(N__12974),
            .I(\Lab_UT.sec1_0 ));
    InMux I__2280 (
            .O(N__12969),
            .I(N__12966));
    LocalMux I__2279 (
            .O(N__12966),
            .I(\Lab_UT.didp.did_alarmMatch_7 ));
    CascadeMux I__2278 (
            .O(N__12963),
            .I(N__12957));
    InMux I__2277 (
            .O(N__12962),
            .I(N__12950));
    InMux I__2276 (
            .O(N__12961),
            .I(N__12950));
    InMux I__2275 (
            .O(N__12960),
            .I(N__12950));
    InMux I__2274 (
            .O(N__12957),
            .I(N__12947));
    LocalMux I__2273 (
            .O(N__12950),
            .I(N__12942));
    LocalMux I__2272 (
            .O(N__12947),
            .I(N__12942));
    Span4Mux_h I__2271 (
            .O(N__12942),
            .I(N__12936));
    InMux I__2270 (
            .O(N__12941),
            .I(N__12929));
    InMux I__2269 (
            .O(N__12940),
            .I(N__12929));
    InMux I__2268 (
            .O(N__12939),
            .I(N__12929));
    Odrv4 I__2267 (
            .O(N__12936),
            .I(\uu2.un15_w_data_displaying_5 ));
    LocalMux I__2266 (
            .O(N__12929),
            .I(\uu2.un15_w_data_displaying_5 ));
    CascadeMux I__2265 (
            .O(N__12924),
            .I(N__12921));
    InMux I__2264 (
            .O(N__12921),
            .I(N__12915));
    InMux I__2263 (
            .O(N__12920),
            .I(N__12915));
    LocalMux I__2262 (
            .O(N__12915),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__2261 (
            .O(N__12912),
            .I(N__12909));
    LocalMux I__2260 (
            .O(N__12909),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    CascadeMux I__2259 (
            .O(N__12906),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    CascadeMux I__2258 (
            .O(N__12903),
            .I(\Lab_UT.didp.countrce1.q_5_3_cascade_ ));
    CascadeMux I__2257 (
            .O(N__12900),
            .I(\Lab_UT.didp.countrce1.q_5_2_cascade_ ));
    InMux I__2256 (
            .O(N__12897),
            .I(N__12894));
    LocalMux I__2255 (
            .O(N__12894),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    InMux I__2254 (
            .O(N__12891),
            .I(N__12888));
    LocalMux I__2253 (
            .O(N__12888),
            .I(N__12884));
    InMux I__2252 (
            .O(N__12887),
            .I(N__12881));
    Span4Mux_s3_v I__2251 (
            .O(N__12884),
            .I(N__12875));
    LocalMux I__2250 (
            .O(N__12881),
            .I(N__12875));
    InMux I__2249 (
            .O(N__12880),
            .I(N__12872));
    Span4Mux_v I__2248 (
            .O(N__12875),
            .I(N__12869));
    LocalMux I__2247 (
            .O(N__12872),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    Odrv4 I__2246 (
            .O(N__12869),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__2245 (
            .O(N__12864),
            .I(N__12861));
    InMux I__2244 (
            .O(N__12861),
            .I(N__12857));
    CascadeMux I__2243 (
            .O(N__12860),
            .I(N__12854));
    LocalMux I__2242 (
            .O(N__12857),
            .I(N__12851));
    InMux I__2241 (
            .O(N__12854),
            .I(N__12848));
    Span4Mux_s3_v I__2240 (
            .O(N__12851),
            .I(N__12843));
    LocalMux I__2239 (
            .O(N__12848),
            .I(N__12843));
    Span4Mux_h I__2238 (
            .O(N__12843),
            .I(N__12838));
    InMux I__2237 (
            .O(N__12842),
            .I(N__12833));
    InMux I__2236 (
            .O(N__12841),
            .I(N__12833));
    Span4Mux_v I__2235 (
            .O(N__12838),
            .I(N__12830));
    LocalMux I__2234 (
            .O(N__12833),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    Odrv4 I__2233 (
            .O(N__12830),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    InMux I__2232 (
            .O(N__12825),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__2231 (
            .O(N__12822),
            .I(N__12818));
    InMux I__2230 (
            .O(N__12821),
            .I(N__12815));
    LocalMux I__2229 (
            .O(N__12818),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__2228 (
            .O(N__12815),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__2227 (
            .O(N__12810),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__2226 (
            .O(N__12807),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__2225 (
            .O(N__12804),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__2224 (
            .O(N__12801),
            .I(N__12791));
    InMux I__2223 (
            .O(N__12800),
            .I(N__12791));
    InMux I__2222 (
            .O(N__12799),
            .I(N__12791));
    InMux I__2221 (
            .O(N__12798),
            .I(N__12788));
    LocalMux I__2220 (
            .O(N__12791),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__2219 (
            .O(N__12788),
            .I(\buart.Z_tx.ser_clk ));
    InMux I__2218 (
            .O(N__12783),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__2217 (
            .O(N__12780),
            .I(N__12777));
    InMux I__2216 (
            .O(N__12777),
            .I(N__12771));
    InMux I__2215 (
            .O(N__12776),
            .I(N__12771));
    LocalMux I__2214 (
            .O(N__12771),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__2213 (
            .O(N__12768),
            .I(N__12765));
    InMux I__2212 (
            .O(N__12765),
            .I(N__12759));
    InMux I__2211 (
            .O(N__12764),
            .I(N__12759));
    LocalMux I__2210 (
            .O(N__12759),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__2209 (
            .O(N__12756),
            .I(N__12752));
    InMux I__2208 (
            .O(N__12755),
            .I(N__12749));
    InMux I__2207 (
            .O(N__12752),
            .I(N__12746));
    LocalMux I__2206 (
            .O(N__12749),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__2205 (
            .O(N__12746),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    CascadeMux I__2204 (
            .O(N__12741),
            .I(\Lab_UT.dispString.N_41_cascade_ ));
    CascadeMux I__2203 (
            .O(N__12738),
            .I(\Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_ ));
    InMux I__2202 (
            .O(N__12735),
            .I(N__12732));
    LocalMux I__2201 (
            .O(N__12732),
            .I(\Lab_UT.dispString.dOut_RNO_0Z0Z_0 ));
    InMux I__2200 (
            .O(N__12729),
            .I(N__12717));
    InMux I__2199 (
            .O(N__12728),
            .I(N__12717));
    InMux I__2198 (
            .O(N__12727),
            .I(N__12717));
    InMux I__2197 (
            .O(N__12726),
            .I(N__12717));
    LocalMux I__2196 (
            .O(N__12717),
            .I(L3_tx_data_0));
    InMux I__2195 (
            .O(N__12714),
            .I(N__12709));
    InMux I__2194 (
            .O(N__12713),
            .I(N__12704));
    InMux I__2193 (
            .O(N__12712),
            .I(N__12704));
    LocalMux I__2192 (
            .O(N__12709),
            .I(\Lab_UT.alarmchar_1 ));
    LocalMux I__2191 (
            .O(N__12704),
            .I(\Lab_UT.alarmchar_1 ));
    CascadeMux I__2190 (
            .O(N__12699),
            .I(N__12691));
    CascadeMux I__2189 (
            .O(N__12698),
            .I(N__12688));
    InMux I__2188 (
            .O(N__12697),
            .I(N__12682));
    InMux I__2187 (
            .O(N__12696),
            .I(N__12676));
    InMux I__2186 (
            .O(N__12695),
            .I(N__12676));
    InMux I__2185 (
            .O(N__12694),
            .I(N__12669));
    InMux I__2184 (
            .O(N__12691),
            .I(N__12669));
    InMux I__2183 (
            .O(N__12688),
            .I(N__12669));
    InMux I__2182 (
            .O(N__12687),
            .I(N__12659));
    InMux I__2181 (
            .O(N__12686),
            .I(N__12659));
    InMux I__2180 (
            .O(N__12685),
            .I(N__12659));
    LocalMux I__2179 (
            .O(N__12682),
            .I(N__12656));
    InMux I__2178 (
            .O(N__12681),
            .I(N__12653));
    LocalMux I__2177 (
            .O(N__12676),
            .I(N__12648));
    LocalMux I__2176 (
            .O(N__12669),
            .I(N__12648));
    InMux I__2175 (
            .O(N__12668),
            .I(N__12641));
    InMux I__2174 (
            .O(N__12667),
            .I(N__12641));
    InMux I__2173 (
            .O(N__12666),
            .I(N__12641));
    LocalMux I__2172 (
            .O(N__12659),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__2171 (
            .O(N__12656),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2170 (
            .O(N__12653),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__2169 (
            .O(N__12648),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2168 (
            .O(N__12641),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    CascadeMux I__2167 (
            .O(N__12630),
            .I(\Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_ ));
    InMux I__2166 (
            .O(N__12627),
            .I(N__12624));
    LocalMux I__2165 (
            .O(N__12624),
            .I(\Lab_UT.dispString.dOut_RNO_0Z0Z_2 ));
    InMux I__2164 (
            .O(N__12621),
            .I(N__12615));
    InMux I__2163 (
            .O(N__12620),
            .I(N__12608));
    InMux I__2162 (
            .O(N__12619),
            .I(N__12608));
    InMux I__2161 (
            .O(N__12618),
            .I(N__12608));
    LocalMux I__2160 (
            .O(N__12615),
            .I(L3_tx_data_2));
    LocalMux I__2159 (
            .O(N__12608),
            .I(L3_tx_data_2));
    InMux I__2158 (
            .O(N__12603),
            .I(N__12591));
    InMux I__2157 (
            .O(N__12602),
            .I(N__12591));
    InMux I__2156 (
            .O(N__12601),
            .I(N__12586));
    InMux I__2155 (
            .O(N__12600),
            .I(N__12586));
    InMux I__2154 (
            .O(N__12599),
            .I(N__12579));
    InMux I__2153 (
            .O(N__12598),
            .I(N__12579));
    InMux I__2152 (
            .O(N__12597),
            .I(N__12579));
    InMux I__2151 (
            .O(N__12596),
            .I(N__12576));
    LocalMux I__2150 (
            .O(N__12591),
            .I(N__12561));
    LocalMux I__2149 (
            .O(N__12586),
            .I(N__12561));
    LocalMux I__2148 (
            .O(N__12579),
            .I(N__12561));
    LocalMux I__2147 (
            .O(N__12576),
            .I(N__12558));
    InMux I__2146 (
            .O(N__12575),
            .I(N__12549));
    InMux I__2145 (
            .O(N__12574),
            .I(N__12549));
    InMux I__2144 (
            .O(N__12573),
            .I(N__12549));
    InMux I__2143 (
            .O(N__12572),
            .I(N__12549));
    InMux I__2142 (
            .O(N__12571),
            .I(N__12540));
    InMux I__2141 (
            .O(N__12570),
            .I(N__12540));
    InMux I__2140 (
            .O(N__12569),
            .I(N__12540));
    InMux I__2139 (
            .O(N__12568),
            .I(N__12540));
    Odrv4 I__2138 (
            .O(N__12561),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2137 (
            .O(N__12558),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2136 (
            .O(N__12549),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2135 (
            .O(N__12540),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    InMux I__2134 (
            .O(N__12531),
            .I(N__12528));
    LocalMux I__2133 (
            .O(N__12528),
            .I(\Lab_UT.dispString.N_32 ));
    CascadeMux I__2132 (
            .O(N__12525),
            .I(N__12514));
    CascadeMux I__2131 (
            .O(N__12524),
            .I(N__12508));
    CascadeMux I__2130 (
            .O(N__12523),
            .I(N__12499));
    CascadeMux I__2129 (
            .O(N__12522),
            .I(N__12496));
    CascadeMux I__2128 (
            .O(N__12521),
            .I(N__12493));
    InMux I__2127 (
            .O(N__12520),
            .I(N__12485));
    InMux I__2126 (
            .O(N__12519),
            .I(N__12485));
    InMux I__2125 (
            .O(N__12518),
            .I(N__12485));
    CascadeMux I__2124 (
            .O(N__12517),
            .I(N__12482));
    InMux I__2123 (
            .O(N__12514),
            .I(N__12471));
    InMux I__2122 (
            .O(N__12513),
            .I(N__12471));
    InMux I__2121 (
            .O(N__12512),
            .I(N__12471));
    InMux I__2120 (
            .O(N__12511),
            .I(N__12471));
    InMux I__2119 (
            .O(N__12508),
            .I(N__12471));
    CascadeMux I__2118 (
            .O(N__12507),
            .I(N__12468));
    CascadeMux I__2117 (
            .O(N__12506),
            .I(N__12465));
    CascadeMux I__2116 (
            .O(N__12505),
            .I(N__12462));
    CascadeMux I__2115 (
            .O(N__12504),
            .I(N__12459));
    InMux I__2114 (
            .O(N__12503),
            .I(N__12456));
    InMux I__2113 (
            .O(N__12502),
            .I(N__12449));
    InMux I__2112 (
            .O(N__12499),
            .I(N__12449));
    InMux I__2111 (
            .O(N__12496),
            .I(N__12449));
    InMux I__2110 (
            .O(N__12493),
            .I(N__12446));
    CascadeMux I__2109 (
            .O(N__12492),
            .I(N__12443));
    LocalMux I__2108 (
            .O(N__12485),
            .I(N__12438));
    InMux I__2107 (
            .O(N__12482),
            .I(N__12435));
    LocalMux I__2106 (
            .O(N__12471),
            .I(N__12432));
    InMux I__2105 (
            .O(N__12468),
            .I(N__12423));
    InMux I__2104 (
            .O(N__12465),
            .I(N__12423));
    InMux I__2103 (
            .O(N__12462),
            .I(N__12423));
    InMux I__2102 (
            .O(N__12459),
            .I(N__12423));
    LocalMux I__2101 (
            .O(N__12456),
            .I(N__12420));
    LocalMux I__2100 (
            .O(N__12449),
            .I(N__12417));
    LocalMux I__2099 (
            .O(N__12446),
            .I(N__12414));
    InMux I__2098 (
            .O(N__12443),
            .I(N__12407));
    InMux I__2097 (
            .O(N__12442),
            .I(N__12407));
    InMux I__2096 (
            .O(N__12441),
            .I(N__12407));
    Span4Mux_v I__2095 (
            .O(N__12438),
            .I(N__12400));
    LocalMux I__2094 (
            .O(N__12435),
            .I(N__12400));
    Span4Mux_h I__2093 (
            .O(N__12432),
            .I(N__12400));
    LocalMux I__2092 (
            .O(N__12423),
            .I(N__12395));
    Span4Mux_s3_h I__2091 (
            .O(N__12420),
            .I(N__12395));
    Odrv4 I__2090 (
            .O(N__12417),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv12 I__2089 (
            .O(N__12414),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    LocalMux I__2088 (
            .O(N__12407),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2087 (
            .O(N__12400),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2086 (
            .O(N__12395),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    InMux I__2085 (
            .O(N__12384),
            .I(N__12381));
    LocalMux I__2084 (
            .O(N__12381),
            .I(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ));
    InMux I__2083 (
            .O(N__12378),
            .I(N__12373));
    InMux I__2082 (
            .O(N__12377),
            .I(N__12368));
    InMux I__2081 (
            .O(N__12376),
            .I(N__12368));
    LocalMux I__2080 (
            .O(N__12373),
            .I(N__12365));
    LocalMux I__2079 (
            .O(N__12368),
            .I(\uu2.un28_w_addr_user_i_0 ));
    Odrv4 I__2078 (
            .O(N__12365),
            .I(\uu2.un28_w_addr_user_i_0 ));
    InMux I__2077 (
            .O(N__12360),
            .I(N__12357));
    LocalMux I__2076 (
            .O(N__12357),
            .I(N__12353));
    CascadeMux I__2075 (
            .O(N__12356),
            .I(N__12349));
    Span4Mux_v I__2074 (
            .O(N__12353),
            .I(N__12345));
    InMux I__2073 (
            .O(N__12352),
            .I(N__12342));
    InMux I__2072 (
            .O(N__12349),
            .I(N__12337));
    InMux I__2071 (
            .O(N__12348),
            .I(N__12337));
    Odrv4 I__2070 (
            .O(N__12345),
            .I(\uu2.N_115 ));
    LocalMux I__2069 (
            .O(N__12342),
            .I(\uu2.N_115 ));
    LocalMux I__2068 (
            .O(N__12337),
            .I(\uu2.N_115 ));
    InMux I__2067 (
            .O(N__12330),
            .I(N__12321));
    InMux I__2066 (
            .O(N__12329),
            .I(N__12321));
    InMux I__2065 (
            .O(N__12328),
            .I(N__12321));
    LocalMux I__2064 (
            .O(N__12321),
            .I(N__12312));
    InMux I__2063 (
            .O(N__12320),
            .I(N__12303));
    InMux I__2062 (
            .O(N__12319),
            .I(N__12303));
    InMux I__2061 (
            .O(N__12318),
            .I(N__12303));
    InMux I__2060 (
            .O(N__12317),
            .I(N__12303));
    InMux I__2059 (
            .O(N__12316),
            .I(N__12300));
    InMux I__2058 (
            .O(N__12315),
            .I(N__12297));
    Span4Mux_v I__2057 (
            .O(N__12312),
            .I(N__12292));
    LocalMux I__2056 (
            .O(N__12303),
            .I(N__12292));
    LocalMux I__2055 (
            .O(N__12300),
            .I(\uu2.N_144 ));
    LocalMux I__2054 (
            .O(N__12297),
            .I(\uu2.N_144 ));
    Odrv4 I__2053 (
            .O(N__12292),
            .I(\uu2.N_144 ));
    InMux I__2052 (
            .O(N__12285),
            .I(N__12277));
    InMux I__2051 (
            .O(N__12284),
            .I(N__12272));
    InMux I__2050 (
            .O(N__12283),
            .I(N__12272));
    InMux I__2049 (
            .O(N__12282),
            .I(N__12269));
    InMux I__2048 (
            .O(N__12281),
            .I(N__12266));
    CascadeMux I__2047 (
            .O(N__12280),
            .I(N__12263));
    LocalMux I__2046 (
            .O(N__12277),
            .I(N__12254));
    LocalMux I__2045 (
            .O(N__12272),
            .I(N__12254));
    LocalMux I__2044 (
            .O(N__12269),
            .I(N__12254));
    LocalMux I__2043 (
            .O(N__12266),
            .I(N__12254));
    InMux I__2042 (
            .O(N__12263),
            .I(N__12251));
    Span4Mux_v I__2041 (
            .O(N__12254),
            .I(N__12248));
    LocalMux I__2040 (
            .O(N__12251),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__2039 (
            .O(N__12248),
            .I(\uu2.w_addr_userZ0Z_4 ));
    InMux I__2038 (
            .O(N__12243),
            .I(N__12240));
    LocalMux I__2037 (
            .O(N__12240),
            .I(N__12235));
    InMux I__2036 (
            .O(N__12239),
            .I(N__12231));
    InMux I__2035 (
            .O(N__12238),
            .I(N__12228));
    Span4Mux_h I__2034 (
            .O(N__12235),
            .I(N__12225));
    InMux I__2033 (
            .O(N__12234),
            .I(N__12222));
    LocalMux I__2032 (
            .O(N__12231),
            .I(o_One_Sec_Pulse));
    LocalMux I__2031 (
            .O(N__12228),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2030 (
            .O(N__12225),
            .I(o_One_Sec_Pulse));
    LocalMux I__2029 (
            .O(N__12222),
            .I(o_One_Sec_Pulse));
    InMux I__2028 (
            .O(N__12213),
            .I(N__12210));
    LocalMux I__2027 (
            .O(N__12210),
            .I(\uu2.bitmapZ0Z_111 ));
    InMux I__2026 (
            .O(N__12207),
            .I(N__12203));
    InMux I__2025 (
            .O(N__12206),
            .I(N__12200));
    LocalMux I__2024 (
            .O(N__12203),
            .I(N__12193));
    LocalMux I__2023 (
            .O(N__12200),
            .I(N__12193));
    InMux I__2022 (
            .O(N__12199),
            .I(N__12190));
    InMux I__2021 (
            .O(N__12198),
            .I(N__12187));
    Span12Mux_s11_h I__2020 (
            .O(N__12193),
            .I(N__12184));
    LocalMux I__2019 (
            .O(N__12190),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__2018 (
            .O(N__12187),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv12 I__2017 (
            .O(N__12184),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__2016 (
            .O(N__12177),
            .I(N__12174));
    LocalMux I__2015 (
            .O(N__12174),
            .I(N__12171));
    Span4Mux_v I__2014 (
            .O(N__12171),
            .I(N__12167));
    InMux I__2013 (
            .O(N__12170),
            .I(N__12164));
    Span4Mux_h I__2012 (
            .O(N__12167),
            .I(N__12161));
    LocalMux I__2011 (
            .O(N__12164),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__2010 (
            .O(N__12161),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__2009 (
            .O(N__12156),
            .I(N__12153));
    LocalMux I__2008 (
            .O(N__12153),
            .I(N__12150));
    Span4Mux_v I__2007 (
            .O(N__12150),
            .I(N__12147));
    Span4Mux_h I__2006 (
            .O(N__12147),
            .I(N__12144));
    Odrv4 I__2005 (
            .O(N__12144),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__2004 (
            .O(N__12141),
            .I(N__12138));
    LocalMux I__2003 (
            .O(N__12138),
            .I(\Lab_UT.dispString.dOutP_1_iv_0_4 ));
    CascadeMux I__2002 (
            .O(N__12135),
            .I(\Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ));
    InMux I__2001 (
            .O(N__12132),
            .I(N__12129));
    LocalMux I__2000 (
            .O(N__12129),
            .I(N__12125));
    CascadeMux I__1999 (
            .O(N__12128),
            .I(N__12120));
    Span4Mux_h I__1998 (
            .O(N__12125),
            .I(N__12116));
    InMux I__1997 (
            .O(N__12124),
            .I(N__12107));
    InMux I__1996 (
            .O(N__12123),
            .I(N__12107));
    InMux I__1995 (
            .O(N__12120),
            .I(N__12107));
    InMux I__1994 (
            .O(N__12119),
            .I(N__12107));
    Odrv4 I__1993 (
            .O(N__12116),
            .I(L3_tx_data_1));
    LocalMux I__1992 (
            .O(N__12107),
            .I(L3_tx_data_1));
    InMux I__1991 (
            .O(N__12102),
            .I(N__12099));
    LocalMux I__1990 (
            .O(N__12099),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_5 ));
    InMux I__1989 (
            .O(N__12096),
            .I(N__12092));
    InMux I__1988 (
            .O(N__12095),
            .I(N__12089));
    LocalMux I__1987 (
            .O(N__12092),
            .I(N__12086));
    LocalMux I__1986 (
            .O(N__12089),
            .I(\uu2.bitmapZ0Z_314 ));
    Odrv12 I__1985 (
            .O(N__12086),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__1984 (
            .O(N__12081),
            .I(N__12078));
    LocalMux I__1983 (
            .O(N__12078),
            .I(N__12075));
    Odrv4 I__1982 (
            .O(N__12075),
            .I(\uu2.bitmapZ0Z_180 ));
    CascadeMux I__1981 (
            .O(N__12072),
            .I(\uu2.N_383_cascade_ ));
    InMux I__1980 (
            .O(N__12069),
            .I(N__12066));
    LocalMux I__1979 (
            .O(N__12066),
            .I(N__12063));
    Odrv4 I__1978 (
            .O(N__12063),
            .I(\uu2.N_215 ));
    InMux I__1977 (
            .O(N__12060),
            .I(N__12057));
    LocalMux I__1976 (
            .O(N__12057),
            .I(N__12054));
    Odrv4 I__1975 (
            .O(N__12054),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    CascadeMux I__1974 (
            .O(N__12051),
            .I(\uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_ ));
    InMux I__1973 (
            .O(N__12048),
            .I(N__12045));
    LocalMux I__1972 (
            .O(N__12045),
            .I(N__12042));
    Odrv12 I__1971 (
            .O(N__12042),
            .I(\uu2.bitmap_RNIS4UH1Z0Z_314 ));
    InMux I__1970 (
            .O(N__12039),
            .I(N__12036));
    LocalMux I__1969 (
            .O(N__12036),
            .I(\uu2.N_397 ));
    InMux I__1968 (
            .O(N__12033),
            .I(N__12030));
    LocalMux I__1967 (
            .O(N__12030),
            .I(\uu2.bitmap_pmux_sn_N_15 ));
    CascadeMux I__1966 (
            .O(N__12027),
            .I(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ));
    InMux I__1965 (
            .O(N__12024),
            .I(N__12021));
    LocalMux I__1964 (
            .O(N__12021),
            .I(\uu2.bitmap_RNIELSJ2Z0Z_111 ));
    InMux I__1963 (
            .O(N__12018),
            .I(N__12014));
    InMux I__1962 (
            .O(N__12017),
            .I(N__12007));
    LocalMux I__1961 (
            .O(N__12014),
            .I(N__12004));
    CascadeMux I__1960 (
            .O(N__12013),
            .I(N__12001));
    CascadeMux I__1959 (
            .O(N__12012),
            .I(N__11993));
    CascadeMux I__1958 (
            .O(N__12011),
            .I(N__11989));
    CascadeMux I__1957 (
            .O(N__12010),
            .I(N__11983));
    LocalMux I__1956 (
            .O(N__12007),
            .I(N__11980));
    Span4Mux_v I__1955 (
            .O(N__12004),
            .I(N__11977));
    InMux I__1954 (
            .O(N__12001),
            .I(N__11968));
    InMux I__1953 (
            .O(N__12000),
            .I(N__11968));
    InMux I__1952 (
            .O(N__11999),
            .I(N__11968));
    InMux I__1951 (
            .O(N__11998),
            .I(N__11968));
    InMux I__1950 (
            .O(N__11997),
            .I(N__11959));
    InMux I__1949 (
            .O(N__11996),
            .I(N__11959));
    InMux I__1948 (
            .O(N__11993),
            .I(N__11959));
    InMux I__1947 (
            .O(N__11992),
            .I(N__11959));
    InMux I__1946 (
            .O(N__11989),
            .I(N__11954));
    InMux I__1945 (
            .O(N__11988),
            .I(N__11954));
    InMux I__1944 (
            .O(N__11987),
            .I(N__11951));
    InMux I__1943 (
            .O(N__11986),
            .I(N__11946));
    InMux I__1942 (
            .O(N__11983),
            .I(N__11946));
    Odrv4 I__1941 (
            .O(N__11980),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1940 (
            .O(N__11977),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1939 (
            .O(N__11968),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1938 (
            .O(N__11959),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1937 (
            .O(N__11954),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1936 (
            .O(N__11951),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1935 (
            .O(N__11946),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__1934 (
            .O(N__11931),
            .I(N__11926));
    CascadeMux I__1933 (
            .O(N__11930),
            .I(N__11921));
    InMux I__1932 (
            .O(N__11929),
            .I(N__11917));
    InMux I__1931 (
            .O(N__11926),
            .I(N__11914));
    InMux I__1930 (
            .O(N__11925),
            .I(N__11905));
    InMux I__1929 (
            .O(N__11924),
            .I(N__11905));
    InMux I__1928 (
            .O(N__11921),
            .I(N__11905));
    InMux I__1927 (
            .O(N__11920),
            .I(N__11905));
    LocalMux I__1926 (
            .O(N__11917),
            .I(N__11902));
    LocalMux I__1925 (
            .O(N__11914),
            .I(\uu2.un21_w_addr_displaying_i ));
    LocalMux I__1924 (
            .O(N__11905),
            .I(\uu2.un21_w_addr_displaying_i ));
    Odrv4 I__1923 (
            .O(N__11902),
            .I(\uu2.un21_w_addr_displaying_i ));
    InMux I__1922 (
            .O(N__11895),
            .I(N__11890));
    CascadeMux I__1921 (
            .O(N__11894),
            .I(N__11883));
    InMux I__1920 (
            .O(N__11893),
            .I(N__11878));
    LocalMux I__1919 (
            .O(N__11890),
            .I(N__11875));
    InMux I__1918 (
            .O(N__11889),
            .I(N__11870));
    InMux I__1917 (
            .O(N__11888),
            .I(N__11870));
    InMux I__1916 (
            .O(N__11887),
            .I(N__11861));
    InMux I__1915 (
            .O(N__11886),
            .I(N__11861));
    InMux I__1914 (
            .O(N__11883),
            .I(N__11861));
    InMux I__1913 (
            .O(N__11882),
            .I(N__11861));
    InMux I__1912 (
            .O(N__11881),
            .I(N__11856));
    LocalMux I__1911 (
            .O(N__11878),
            .I(N__11853));
    Span4Mux_h I__1910 (
            .O(N__11875),
            .I(N__11850));
    LocalMux I__1909 (
            .O(N__11870),
            .I(N__11847));
    LocalMux I__1908 (
            .O(N__11861),
            .I(N__11844));
    InMux I__1907 (
            .O(N__11860),
            .I(N__11839));
    InMux I__1906 (
            .O(N__11859),
            .I(N__11839));
    LocalMux I__1905 (
            .O(N__11856),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__1904 (
            .O(N__11853),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__1903 (
            .O(N__11850),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__1902 (
            .O(N__11847),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__1901 (
            .O(N__11844),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__1900 (
            .O(N__11839),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    InMux I__1899 (
            .O(N__11826),
            .I(N__11821));
    InMux I__1898 (
            .O(N__11825),
            .I(N__11818));
    CascadeMux I__1897 (
            .O(N__11824),
            .I(N__11815));
    LocalMux I__1896 (
            .O(N__11821),
            .I(N__11808));
    LocalMux I__1895 (
            .O(N__11818),
            .I(N__11805));
    InMux I__1894 (
            .O(N__11815),
            .I(N__11802));
    InMux I__1893 (
            .O(N__11814),
            .I(N__11793));
    InMux I__1892 (
            .O(N__11813),
            .I(N__11793));
    InMux I__1891 (
            .O(N__11812),
            .I(N__11793));
    InMux I__1890 (
            .O(N__11811),
            .I(N__11793));
    Span4Mux_h I__1889 (
            .O(N__11808),
            .I(N__11788));
    Span4Mux_h I__1888 (
            .O(N__11805),
            .I(N__11788));
    LocalMux I__1887 (
            .O(N__11802),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1886 (
            .O(N__11793),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__1885 (
            .O(N__11788),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__1884 (
            .O(N__11781),
            .I(N__11776));
    CascadeMux I__1883 (
            .O(N__11780),
            .I(N__11772));
    CascadeMux I__1882 (
            .O(N__11779),
            .I(N__11769));
    InMux I__1881 (
            .O(N__11776),
            .I(N__11765));
    InMux I__1880 (
            .O(N__11775),
            .I(N__11758));
    InMux I__1879 (
            .O(N__11772),
            .I(N__11758));
    InMux I__1878 (
            .O(N__11769),
            .I(N__11758));
    CascadeMux I__1877 (
            .O(N__11768),
            .I(N__11755));
    LocalMux I__1876 (
            .O(N__11765),
            .I(N__11749));
    LocalMux I__1875 (
            .O(N__11758),
            .I(N__11749));
    InMux I__1874 (
            .O(N__11755),
            .I(N__11746));
    InMux I__1873 (
            .O(N__11754),
            .I(N__11743));
    Span4Mux_h I__1872 (
            .O(N__11749),
            .I(N__11740));
    LocalMux I__1871 (
            .O(N__11746),
            .I(\uu2.w_addr_userZ0Z_1 ));
    LocalMux I__1870 (
            .O(N__11743),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1869 (
            .O(N__11740),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__1868 (
            .O(N__11733),
            .I(N__11729));
    InMux I__1867 (
            .O(N__11732),
            .I(N__11726));
    InMux I__1866 (
            .O(N__11729),
            .I(N__11723));
    LocalMux I__1865 (
            .O(N__11726),
            .I(\uu2.un33_w_data_displaying ));
    LocalMux I__1864 (
            .O(N__11723),
            .I(\uu2.un33_w_data_displaying ));
    InMux I__1863 (
            .O(N__11718),
            .I(N__11714));
    CascadeMux I__1862 (
            .O(N__11717),
            .I(N__11701));
    LocalMux I__1861 (
            .O(N__11714),
            .I(N__11696));
    InMux I__1860 (
            .O(N__11713),
            .I(N__11693));
    InMux I__1859 (
            .O(N__11712),
            .I(N__11690));
    InMux I__1858 (
            .O(N__11711),
            .I(N__11685));
    InMux I__1857 (
            .O(N__11710),
            .I(N__11685));
    InMux I__1856 (
            .O(N__11709),
            .I(N__11680));
    InMux I__1855 (
            .O(N__11708),
            .I(N__11680));
    InMux I__1854 (
            .O(N__11707),
            .I(N__11675));
    InMux I__1853 (
            .O(N__11706),
            .I(N__11675));
    InMux I__1852 (
            .O(N__11705),
            .I(N__11670));
    InMux I__1851 (
            .O(N__11704),
            .I(N__11670));
    InMux I__1850 (
            .O(N__11701),
            .I(N__11667));
    InMux I__1849 (
            .O(N__11700),
            .I(N__11662));
    InMux I__1848 (
            .O(N__11699),
            .I(N__11662));
    Span4Mux_h I__1847 (
            .O(N__11696),
            .I(N__11653));
    LocalMux I__1846 (
            .O(N__11693),
            .I(N__11653));
    LocalMux I__1845 (
            .O(N__11690),
            .I(N__11653));
    LocalMux I__1844 (
            .O(N__11685),
            .I(N__11653));
    LocalMux I__1843 (
            .O(N__11680),
            .I(N__11650));
    LocalMux I__1842 (
            .O(N__11675),
            .I(N__11645));
    LocalMux I__1841 (
            .O(N__11670),
            .I(N__11645));
    LocalMux I__1840 (
            .O(N__11667),
            .I(N__11640));
    LocalMux I__1839 (
            .O(N__11662),
            .I(N__11640));
    Span4Mux_v I__1838 (
            .O(N__11653),
            .I(N__11635));
    Span4Mux_v I__1837 (
            .O(N__11650),
            .I(N__11635));
    Span4Mux_v I__1836 (
            .O(N__11645),
            .I(N__11632));
    Odrv12 I__1835 (
            .O(N__11640),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    Odrv4 I__1834 (
            .O(N__11635),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    Odrv4 I__1833 (
            .O(N__11632),
            .I(\uu2.w_addr_i_0_tzZ0Z_0 ));
    CascadeMux I__1832 (
            .O(N__11625),
            .I(\uu2.un21_w_addr_displaying_i_cascade_ ));
    InMux I__1831 (
            .O(N__11622),
            .I(N__11619));
    LocalMux I__1830 (
            .O(N__11619),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    InMux I__1829 (
            .O(N__11616),
            .I(N__11613));
    LocalMux I__1828 (
            .O(N__11613),
            .I(N__11610));
    Odrv12 I__1827 (
            .O(N__11610),
            .I(\uu2.bitmap_pmux_sn_N_65 ));
    CascadeMux I__1826 (
            .O(N__11607),
            .I(\uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ));
    CascadeMux I__1825 (
            .O(N__11604),
            .I(N__11600));
    InMux I__1824 (
            .O(N__11603),
            .I(N__11594));
    InMux I__1823 (
            .O(N__11600),
            .I(N__11594));
    InMux I__1822 (
            .O(N__11599),
            .I(N__11591));
    LocalMux I__1821 (
            .O(N__11594),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    LocalMux I__1820 (
            .O(N__11591),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    InMux I__1819 (
            .O(N__11586),
            .I(N__11583));
    LocalMux I__1818 (
            .O(N__11583),
            .I(\uu2.bitmap_pmux_sn_i7_mux_0 ));
    InMux I__1817 (
            .O(N__11580),
            .I(N__11577));
    LocalMux I__1816 (
            .O(N__11577),
            .I(N__11572));
    InMux I__1815 (
            .O(N__11576),
            .I(N__11567));
    InMux I__1814 (
            .O(N__11575),
            .I(N__11567));
    Odrv4 I__1813 (
            .O(N__11572),
            .I(\uu2.un15_w_data_displaying_2 ));
    LocalMux I__1812 (
            .O(N__11567),
            .I(\uu2.un15_w_data_displaying_2 ));
    InMux I__1811 (
            .O(N__11562),
            .I(N__11559));
    LocalMux I__1810 (
            .O(N__11559),
            .I(\uu2.bitmapZ0Z_69 ));
    CascadeMux I__1809 (
            .O(N__11556),
            .I(N__11553));
    InMux I__1808 (
            .O(N__11553),
            .I(N__11550));
    LocalMux I__1807 (
            .O(N__11550),
            .I(\uu2.bitmapZ0Z_197 ));
    CascadeMux I__1806 (
            .O(N__11547),
            .I(\uu2.un437_ci_0_cascade_ ));
    InMux I__1805 (
            .O(N__11544),
            .I(N__11539));
    CascadeMux I__1804 (
            .O(N__11543),
            .I(N__11536));
    CascadeMux I__1803 (
            .O(N__11542),
            .I(N__11533));
    LocalMux I__1802 (
            .O(N__11539),
            .I(N__11530));
    InMux I__1801 (
            .O(N__11536),
            .I(N__11525));
    InMux I__1800 (
            .O(N__11533),
            .I(N__11525));
    Span4Mux_v I__1799 (
            .O(N__11530),
            .I(N__11522));
    LocalMux I__1798 (
            .O(N__11525),
            .I(N__11519));
    Odrv4 I__1797 (
            .O(N__11522),
            .I(L3_tx_data_6));
    Odrv4 I__1796 (
            .O(N__11519),
            .I(L3_tx_data_6));
    InMux I__1795 (
            .O(N__11514),
            .I(N__11511));
    LocalMux I__1794 (
            .O(N__11511),
            .I(N__11508));
    Span4Mux_h I__1793 (
            .O(N__11508),
            .I(N__11505));
    Odrv4 I__1792 (
            .O(N__11505),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__1791 (
            .O(N__11502),
            .I(N__11499));
    LocalMux I__1790 (
            .O(N__11499),
            .I(\uu2.un31_w_data_displaying_2 ));
    CascadeMux I__1789 (
            .O(N__11496),
            .I(N__11493));
    InMux I__1788 (
            .O(N__11493),
            .I(N__11490));
    LocalMux I__1787 (
            .O(N__11490),
            .I(N__11487));
    Span4Mux_v I__1786 (
            .O(N__11487),
            .I(N__11484));
    Odrv4 I__1785 (
            .O(N__11484),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__1784 (
            .O(N__11481),
            .I(N__11478));
    LocalMux I__1783 (
            .O(N__11478),
            .I(\uu2.bitmapZ0Z_72 ));
    CascadeMux I__1782 (
            .O(N__11475),
            .I(N__11472));
    InMux I__1781 (
            .O(N__11472),
            .I(N__11469));
    LocalMux I__1780 (
            .O(N__11469),
            .I(\uu2.bitmapZ0Z_200 ));
    CascadeMux I__1779 (
            .O(N__11466),
            .I(\uu2.bitmap_pmux_24_i_m2_bm_1_cascade_ ));
    InMux I__1778 (
            .O(N__11463),
            .I(N__11460));
    LocalMux I__1777 (
            .O(N__11460),
            .I(\uu2.bitmap_RNI1UT12Z0Z_75 ));
    InMux I__1776 (
            .O(N__11457),
            .I(N__11454));
    LocalMux I__1775 (
            .O(N__11454),
            .I(\uu2.bitmapZ0Z_75 ));
    InMux I__1774 (
            .O(N__11451),
            .I(N__11448));
    LocalMux I__1773 (
            .O(N__11448),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__1772 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__1771 (
            .O(N__11442),
            .I(N__11439));
    Span4Mux_v I__1770 (
            .O(N__11439),
            .I(N__11430));
    InMux I__1769 (
            .O(N__11438),
            .I(N__11417));
    InMux I__1768 (
            .O(N__11437),
            .I(N__11417));
    InMux I__1767 (
            .O(N__11436),
            .I(N__11417));
    InMux I__1766 (
            .O(N__11435),
            .I(N__11417));
    InMux I__1765 (
            .O(N__11434),
            .I(N__11417));
    InMux I__1764 (
            .O(N__11433),
            .I(N__11417));
    Odrv4 I__1763 (
            .O(N__11430),
            .I(\Lab_UT.min2_2 ));
    LocalMux I__1762 (
            .O(N__11417),
            .I(\Lab_UT.min2_2 ));
    InMux I__1761 (
            .O(N__11412),
            .I(N__11409));
    LocalMux I__1760 (
            .O(N__11409),
            .I(N__11403));
    CascadeMux I__1759 (
            .O(N__11408),
            .I(N__11399));
    CascadeMux I__1758 (
            .O(N__11407),
            .I(N__11396));
    CascadeMux I__1757 (
            .O(N__11406),
            .I(N__11393));
    Sp12to4 I__1756 (
            .O(N__11403),
            .I(N__11388));
    InMux I__1755 (
            .O(N__11402),
            .I(N__11375));
    InMux I__1754 (
            .O(N__11399),
            .I(N__11375));
    InMux I__1753 (
            .O(N__11396),
            .I(N__11375));
    InMux I__1752 (
            .O(N__11393),
            .I(N__11375));
    InMux I__1751 (
            .O(N__11392),
            .I(N__11375));
    InMux I__1750 (
            .O(N__11391),
            .I(N__11375));
    Odrv12 I__1749 (
            .O(N__11388),
            .I(\Lab_UT.min2_1 ));
    LocalMux I__1748 (
            .O(N__11375),
            .I(\Lab_UT.min2_1 ));
    CascadeMux I__1747 (
            .O(N__11370),
            .I(N__11367));
    InMux I__1746 (
            .O(N__11367),
            .I(N__11364));
    LocalMux I__1745 (
            .O(N__11364),
            .I(N__11358));
    CascadeMux I__1744 (
            .O(N__11363),
            .I(N__11355));
    CascadeMux I__1743 (
            .O(N__11362),
            .I(N__11349));
    CascadeMux I__1742 (
            .O(N__11361),
            .I(N__11346));
    Span4Mux_v I__1741 (
            .O(N__11358),
            .I(N__11343));
    InMux I__1740 (
            .O(N__11355),
            .I(N__11330));
    InMux I__1739 (
            .O(N__11354),
            .I(N__11330));
    InMux I__1738 (
            .O(N__11353),
            .I(N__11330));
    InMux I__1737 (
            .O(N__11352),
            .I(N__11330));
    InMux I__1736 (
            .O(N__11349),
            .I(N__11330));
    InMux I__1735 (
            .O(N__11346),
            .I(N__11330));
    Odrv4 I__1734 (
            .O(N__11343),
            .I(\Lab_UT.min2_3 ));
    LocalMux I__1733 (
            .O(N__11330),
            .I(\Lab_UT.min2_3 ));
    InMux I__1732 (
            .O(N__11325),
            .I(N__11322));
    LocalMux I__1731 (
            .O(N__11322),
            .I(N__11319));
    Span4Mux_v I__1730 (
            .O(N__11319),
            .I(N__11310));
    InMux I__1729 (
            .O(N__11318),
            .I(N__11297));
    InMux I__1728 (
            .O(N__11317),
            .I(N__11297));
    InMux I__1727 (
            .O(N__11316),
            .I(N__11297));
    InMux I__1726 (
            .O(N__11315),
            .I(N__11297));
    InMux I__1725 (
            .O(N__11314),
            .I(N__11297));
    InMux I__1724 (
            .O(N__11313),
            .I(N__11297));
    Odrv4 I__1723 (
            .O(N__11310),
            .I(\Lab_UT.min2_0 ));
    LocalMux I__1722 (
            .O(N__11297),
            .I(\Lab_UT.min2_0 ));
    CascadeMux I__1721 (
            .O(N__11292),
            .I(N__11285));
    CascadeMux I__1720 (
            .O(N__11291),
            .I(N__11282));
    CascadeMux I__1719 (
            .O(N__11290),
            .I(N__11278));
    CascadeMux I__1718 (
            .O(N__11289),
            .I(N__11274));
    InMux I__1717 (
            .O(N__11288),
            .I(N__11269));
    InMux I__1716 (
            .O(N__11285),
            .I(N__11269));
    InMux I__1715 (
            .O(N__11282),
            .I(N__11258));
    InMux I__1714 (
            .O(N__11281),
            .I(N__11258));
    InMux I__1713 (
            .O(N__11278),
            .I(N__11258));
    InMux I__1712 (
            .O(N__11277),
            .I(N__11258));
    InMux I__1711 (
            .O(N__11274),
            .I(N__11258));
    LocalMux I__1710 (
            .O(N__11269),
            .I(\Lab_UT.sec2_3 ));
    LocalMux I__1709 (
            .O(N__11258),
            .I(\Lab_UT.sec2_3 ));
    CascadeMux I__1708 (
            .O(N__11253),
            .I(N__11248));
    CascadeMux I__1707 (
            .O(N__11252),
            .I(N__11244));
    InMux I__1706 (
            .O(N__11251),
            .I(N__11230));
    InMux I__1705 (
            .O(N__11248),
            .I(N__11230));
    InMux I__1704 (
            .O(N__11247),
            .I(N__11230));
    InMux I__1703 (
            .O(N__11244),
            .I(N__11230));
    InMux I__1702 (
            .O(N__11243),
            .I(N__11230));
    InMux I__1701 (
            .O(N__11242),
            .I(N__11225));
    InMux I__1700 (
            .O(N__11241),
            .I(N__11225));
    LocalMux I__1699 (
            .O(N__11230),
            .I(N__11222));
    LocalMux I__1698 (
            .O(N__11225),
            .I(\Lab_UT.sec2_2 ));
    Odrv4 I__1697 (
            .O(N__11222),
            .I(\Lab_UT.sec2_2 ));
    CascadeMux I__1696 (
            .O(N__11217),
            .I(N__11209));
    InMux I__1695 (
            .O(N__11216),
            .I(N__11197));
    InMux I__1694 (
            .O(N__11215),
            .I(N__11197));
    InMux I__1693 (
            .O(N__11214),
            .I(N__11197));
    InMux I__1692 (
            .O(N__11213),
            .I(N__11197));
    InMux I__1691 (
            .O(N__11212),
            .I(N__11197));
    InMux I__1690 (
            .O(N__11209),
            .I(N__11192));
    InMux I__1689 (
            .O(N__11208),
            .I(N__11192));
    LocalMux I__1688 (
            .O(N__11197),
            .I(N__11189));
    LocalMux I__1687 (
            .O(N__11192),
            .I(\Lab_UT.sec2_1 ));
    Odrv4 I__1686 (
            .O(N__11189),
            .I(\Lab_UT.sec2_1 ));
    InMux I__1685 (
            .O(N__11184),
            .I(N__11181));
    LocalMux I__1684 (
            .O(N__11181),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__1683 (
            .O(N__11178),
            .I(N__11175));
    LocalMux I__1682 (
            .O(N__11175),
            .I(\uu2.bitmapZ0Z_58 ));
    CascadeMux I__1681 (
            .O(N__11172),
            .I(\uu2.N_216_cascade_ ));
    InMux I__1680 (
            .O(N__11169),
            .I(N__11151));
    InMux I__1679 (
            .O(N__11168),
            .I(N__11151));
    InMux I__1678 (
            .O(N__11167),
            .I(N__11151));
    InMux I__1677 (
            .O(N__11166),
            .I(N__11151));
    InMux I__1676 (
            .O(N__11165),
            .I(N__11151));
    InMux I__1675 (
            .O(N__11164),
            .I(N__11151));
    LocalMux I__1674 (
            .O(N__11151),
            .I(N__11148));
    IoSpan4Mux I__1673 (
            .O(N__11148),
            .I(N__11144));
    InMux I__1672 (
            .O(N__11147),
            .I(N__11141));
    Odrv4 I__1671 (
            .O(N__11144),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__1670 (
            .O(N__11141),
            .I(\Lab_UT.sec1_1 ));
    CascadeMux I__1669 (
            .O(N__11136),
            .I(N__11130));
    CascadeMux I__1668 (
            .O(N__11135),
            .I(N__11127));
    CascadeMux I__1667 (
            .O(N__11134),
            .I(N__11124));
    CascadeMux I__1666 (
            .O(N__11133),
            .I(N__11121));
    InMux I__1665 (
            .O(N__11130),
            .I(N__11105));
    InMux I__1664 (
            .O(N__11127),
            .I(N__11105));
    InMux I__1663 (
            .O(N__11124),
            .I(N__11105));
    InMux I__1662 (
            .O(N__11121),
            .I(N__11105));
    InMux I__1661 (
            .O(N__11120),
            .I(N__11105));
    InMux I__1660 (
            .O(N__11119),
            .I(N__11105));
    CascadeMux I__1659 (
            .O(N__11118),
            .I(N__11102));
    LocalMux I__1658 (
            .O(N__11105),
            .I(N__11099));
    InMux I__1657 (
            .O(N__11102),
            .I(N__11096));
    Odrv4 I__1656 (
            .O(N__11099),
            .I(\Lab_UT.sec1_2 ));
    LocalMux I__1655 (
            .O(N__11096),
            .I(\Lab_UT.sec1_2 ));
    CascadeMux I__1654 (
            .O(N__11091),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    CascadeMux I__1653 (
            .O(N__11088),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    CascadeMux I__1652 (
            .O(N__11085),
            .I(\buart.Z_tx.un1_bitcount_c2_cascade_ ));
    InMux I__1651 (
            .O(N__11082),
            .I(N__11077));
    InMux I__1650 (
            .O(N__11081),
            .I(N__11072));
    InMux I__1649 (
            .O(N__11080),
            .I(N__11072));
    LocalMux I__1648 (
            .O(N__11077),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__1647 (
            .O(N__11072),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    InMux I__1646 (
            .O(N__11067),
            .I(N__11061));
    InMux I__1645 (
            .O(N__11066),
            .I(N__11058));
    InMux I__1644 (
            .O(N__11065),
            .I(N__11051));
    InMux I__1643 (
            .O(N__11064),
            .I(N__11051));
    LocalMux I__1642 (
            .O(N__11061),
            .I(N__11046));
    LocalMux I__1641 (
            .O(N__11058),
            .I(N__11046));
    InMux I__1640 (
            .O(N__11057),
            .I(N__11041));
    InMux I__1639 (
            .O(N__11056),
            .I(N__11041));
    LocalMux I__1638 (
            .O(N__11051),
            .I(N__11036));
    Span4Mux_v I__1637 (
            .O(N__11046),
            .I(N__11036));
    LocalMux I__1636 (
            .O(N__11041),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    Odrv4 I__1635 (
            .O(N__11036),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    CascadeMux I__1634 (
            .O(N__11031),
            .I(N__11028));
    InMux I__1633 (
            .O(N__11028),
            .I(N__11019));
    InMux I__1632 (
            .O(N__11027),
            .I(N__11019));
    InMux I__1631 (
            .O(N__11026),
            .I(N__11019));
    LocalMux I__1630 (
            .O(N__11019),
            .I(N__11016));
    Span4Mux_v I__1629 (
            .O(N__11016),
            .I(N__11004));
    InMux I__1628 (
            .O(N__11015),
            .I(N__10993));
    InMux I__1627 (
            .O(N__11014),
            .I(N__10993));
    InMux I__1626 (
            .O(N__11013),
            .I(N__10993));
    InMux I__1625 (
            .O(N__11012),
            .I(N__10993));
    InMux I__1624 (
            .O(N__11011),
            .I(N__10993));
    InMux I__1623 (
            .O(N__11010),
            .I(N__10990));
    InMux I__1622 (
            .O(N__11009),
            .I(N__10985));
    InMux I__1621 (
            .O(N__11008),
            .I(N__10985));
    CascadeMux I__1620 (
            .O(N__11007),
            .I(N__10978));
    Span4Mux_v I__1619 (
            .O(N__11004),
            .I(N__10975));
    LocalMux I__1618 (
            .O(N__10993),
            .I(N__10968));
    LocalMux I__1617 (
            .O(N__10990),
            .I(N__10968));
    LocalMux I__1616 (
            .O(N__10985),
            .I(N__10968));
    InMux I__1615 (
            .O(N__10984),
            .I(N__10959));
    InMux I__1614 (
            .O(N__10983),
            .I(N__10959));
    InMux I__1613 (
            .O(N__10982),
            .I(N__10959));
    InMux I__1612 (
            .O(N__10981),
            .I(N__10959));
    InMux I__1611 (
            .O(N__10978),
            .I(N__10956));
    Span4Mux_h I__1610 (
            .O(N__10975),
            .I(N__10953));
    Span4Mux_v I__1609 (
            .O(N__10968),
            .I(N__10948));
    LocalMux I__1608 (
            .O(N__10959),
            .I(N__10948));
    LocalMux I__1607 (
            .O(N__10956),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1606 (
            .O(N__10953),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__1605 (
            .O(N__10948),
            .I(vbuf_tx_data_rdy));
    CascadeMux I__1604 (
            .O(N__10941),
            .I(N__10937));
    InMux I__1603 (
            .O(N__10940),
            .I(N__10929));
    InMux I__1602 (
            .O(N__10937),
            .I(N__10929));
    InMux I__1601 (
            .O(N__10936),
            .I(N__10924));
    InMux I__1600 (
            .O(N__10935),
            .I(N__10924));
    InMux I__1599 (
            .O(N__10934),
            .I(N__10921));
    LocalMux I__1598 (
            .O(N__10929),
            .I(N__10916));
    LocalMux I__1597 (
            .O(N__10924),
            .I(N__10916));
    LocalMux I__1596 (
            .O(N__10921),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    Odrv4 I__1595 (
            .O(N__10916),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__1594 (
            .O(N__10911),
            .I(N__10899));
    InMux I__1593 (
            .O(N__10910),
            .I(N__10899));
    InMux I__1592 (
            .O(N__10909),
            .I(N__10899));
    InMux I__1591 (
            .O(N__10908),
            .I(N__10899));
    LocalMux I__1590 (
            .O(N__10899),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__1589 (
            .O(N__10896),
            .I(N__10893));
    LocalMux I__1588 (
            .O(N__10893),
            .I(\uu2.bitmapZ0Z_90 ));
    CascadeMux I__1587 (
            .O(N__10890),
            .I(N__10887));
    InMux I__1586 (
            .O(N__10887),
            .I(N__10884));
    LocalMux I__1585 (
            .O(N__10884),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__1584 (
            .O(N__10881),
            .I(N__10878));
    LocalMux I__1583 (
            .O(N__10878),
            .I(\uu2.bitmap_pmux_25_bm_1 ));
    InMux I__1582 (
            .O(N__10875),
            .I(N__10872));
    LocalMux I__1581 (
            .O(N__10872),
            .I(\Lab_UT.dispString.N_50 ));
    CascadeMux I__1580 (
            .O(N__10869),
            .I(\Lab_UT.dispString.N_28_cascade_ ));
    InMux I__1579 (
            .O(N__10866),
            .I(N__10863));
    LocalMux I__1578 (
            .O(N__10863),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_3 ));
    CascadeMux I__1577 (
            .O(N__10860),
            .I(\buart.Z_tx.un1_bitcount_c3_cascade_ ));
    InMux I__1576 (
            .O(N__10857),
            .I(N__10853));
    InMux I__1575 (
            .O(N__10856),
            .I(N__10850));
    LocalMux I__1574 (
            .O(N__10853),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__1573 (
            .O(N__10850),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__1572 (
            .O(N__10845),
            .I(N__10841));
    InMux I__1571 (
            .O(N__10844),
            .I(N__10838));
    InMux I__1570 (
            .O(N__10841),
            .I(N__10834));
    LocalMux I__1569 (
            .O(N__10838),
            .I(N__10831));
    InMux I__1568 (
            .O(N__10837),
            .I(N__10828));
    LocalMux I__1567 (
            .O(N__10834),
            .I(N__10825));
    Odrv4 I__1566 (
            .O(N__10831),
            .I(\uu2.N_361 ));
    LocalMux I__1565 (
            .O(N__10828),
            .I(\uu2.N_361 ));
    Odrv4 I__1564 (
            .O(N__10825),
            .I(\uu2.N_361 ));
    CascadeMux I__1563 (
            .O(N__10818),
            .I(\uu2.mem0.w_data_0_a2_0_4_cascade_ ));
    InMux I__1562 (
            .O(N__10815),
            .I(N__10812));
    LocalMux I__1561 (
            .O(N__10812),
            .I(N__10809));
    Span4Mux_s3_h I__1560 (
            .O(N__10809),
            .I(N__10806));
    Odrv4 I__1559 (
            .O(N__10806),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1558 (
            .O(N__10803),
            .I(N__10798));
    InMux I__1557 (
            .O(N__10802),
            .I(N__10795));
    InMux I__1556 (
            .O(N__10801),
            .I(N__10792));
    LocalMux I__1555 (
            .O(N__10798),
            .I(N__10789));
    LocalMux I__1554 (
            .O(N__10795),
            .I(N__10784));
    LocalMux I__1553 (
            .O(N__10792),
            .I(N__10784));
    Odrv4 I__1552 (
            .O(N__10789),
            .I(L3_tx_data_5));
    Odrv4 I__1551 (
            .O(N__10784),
            .I(L3_tx_data_5));
    InMux I__1550 (
            .O(N__10779),
            .I(N__10773));
    InMux I__1549 (
            .O(N__10778),
            .I(N__10773));
    LocalMux I__1548 (
            .O(N__10773),
            .I(N__10770));
    Odrv4 I__1547 (
            .O(N__10770),
            .I(L3_tx_data_4));
    InMux I__1546 (
            .O(N__10767),
            .I(N__10755));
    InMux I__1545 (
            .O(N__10766),
            .I(N__10755));
    InMux I__1544 (
            .O(N__10765),
            .I(N__10755));
    InMux I__1543 (
            .O(N__10764),
            .I(N__10755));
    LocalMux I__1542 (
            .O(N__10755),
            .I(\uu2.N_109 ));
    InMux I__1541 (
            .O(N__10752),
            .I(N__10746));
    InMux I__1540 (
            .O(N__10751),
            .I(N__10746));
    LocalMux I__1539 (
            .O(N__10746),
            .I(\uu2.N_111 ));
    CascadeMux I__1538 (
            .O(N__10743),
            .I(\uu2.N_109_cascade_ ));
    InMux I__1537 (
            .O(N__10740),
            .I(N__10730));
    InMux I__1536 (
            .O(N__10739),
            .I(N__10730));
    InMux I__1535 (
            .O(N__10738),
            .I(N__10727));
    InMux I__1534 (
            .O(N__10737),
            .I(N__10720));
    InMux I__1533 (
            .O(N__10736),
            .I(N__10720));
    InMux I__1532 (
            .O(N__10735),
            .I(N__10720));
    LocalMux I__1531 (
            .O(N__10730),
            .I(N__10717));
    LocalMux I__1530 (
            .O(N__10727),
            .I(L3_tx_data_rdy));
    LocalMux I__1529 (
            .O(N__10720),
            .I(L3_tx_data_rdy));
    Odrv4 I__1528 (
            .O(N__10717),
            .I(L3_tx_data_rdy));
    CascadeMux I__1527 (
            .O(N__10710),
            .I(N__10705));
    InMux I__1526 (
            .O(N__10709),
            .I(N__10701));
    InMux I__1525 (
            .O(N__10708),
            .I(N__10694));
    InMux I__1524 (
            .O(N__10705),
            .I(N__10694));
    InMux I__1523 (
            .O(N__10704),
            .I(N__10694));
    LocalMux I__1522 (
            .O(N__10701),
            .I(N__10691));
    LocalMux I__1521 (
            .O(N__10694),
            .I(N__10688));
    Span4Mux_v I__1520 (
            .O(N__10691),
            .I(N__10685));
    Odrv4 I__1519 (
            .O(N__10688),
            .I(\Lab_UT.dispString.N_61 ));
    Odrv4 I__1518 (
            .O(N__10685),
            .I(\Lab_UT.dispString.N_61 ));
    InMux I__1517 (
            .O(N__10680),
            .I(N__10677));
    LocalMux I__1516 (
            .O(N__10677),
            .I(N__10674));
    Span4Mux_h I__1515 (
            .O(N__10674),
            .I(N__10671));
    Odrv4 I__1514 (
            .O(N__10671),
            .I(\Lab_UT.dispString.un46_dOutP_i_m_3 ));
    CascadeMux I__1513 (
            .O(N__10668),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_3_cascade_ ));
    InMux I__1512 (
            .O(N__10665),
            .I(N__10662));
    LocalMux I__1511 (
            .O(N__10662),
            .I(\Lab_UT.dispString.dOutP_6 ));
    InMux I__1510 (
            .O(N__10659),
            .I(N__10656));
    LocalMux I__1509 (
            .O(N__10656),
            .I(N__10653));
    Span12Mux_s4_v I__1508 (
            .O(N__10653),
            .I(N__10648));
    InMux I__1507 (
            .O(N__10652),
            .I(N__10643));
    InMux I__1506 (
            .O(N__10651),
            .I(N__10643));
    Odrv12 I__1505 (
            .O(N__10648),
            .I(L3_tx_data_3));
    LocalMux I__1504 (
            .O(N__10643),
            .I(L3_tx_data_3));
    CascadeMux I__1503 (
            .O(N__10638),
            .I(\uu2.N_111_cascade_ ));
    SRMux I__1502 (
            .O(N__10635),
            .I(N__10631));
    CEMux I__1501 (
            .O(N__10634),
            .I(N__10628));
    LocalMux I__1500 (
            .O(N__10631),
            .I(N__10625));
    LocalMux I__1499 (
            .O(N__10628),
            .I(N__10622));
    Span4Mux_v I__1498 (
            .O(N__10625),
            .I(N__10617));
    Span4Mux_h I__1497 (
            .O(N__10622),
            .I(N__10617));
    Span4Mux_v I__1496 (
            .O(N__10617),
            .I(N__10614));
    Odrv4 I__1495 (
            .O(N__10614),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1494 (
            .O(N__10611),
            .I(\uu2.mem0.w_data_i_a2_1_0_cascade_ ));
    InMux I__1493 (
            .O(N__10608),
            .I(N__10605));
    LocalMux I__1492 (
            .O(N__10605),
            .I(N__10602));
    Span4Mux_s3_h I__1491 (
            .O(N__10602),
            .I(N__10599));
    Odrv4 I__1490 (
            .O(N__10599),
            .I(\uu2.mem0.N_82_i ));
    CascadeMux I__1489 (
            .O(N__10596),
            .I(N__10593));
    InMux I__1488 (
            .O(N__10593),
            .I(N__10590));
    LocalMux I__1487 (
            .O(N__10590),
            .I(\uu2.mem0.N_110 ));
    InMux I__1486 (
            .O(N__10587),
            .I(N__10579));
    InMux I__1485 (
            .O(N__10586),
            .I(N__10576));
    InMux I__1484 (
            .O(N__10585),
            .I(N__10567));
    InMux I__1483 (
            .O(N__10584),
            .I(N__10567));
    InMux I__1482 (
            .O(N__10583),
            .I(N__10567));
    InMux I__1481 (
            .O(N__10582),
            .I(N__10567));
    LocalMux I__1480 (
            .O(N__10579),
            .I(N__10564));
    LocalMux I__1479 (
            .O(N__10576),
            .I(N__10561));
    LocalMux I__1478 (
            .O(N__10567),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__1477 (
            .O(N__10564),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__1476 (
            .O(N__10561),
            .I(\uu2.w_addr_userZ0Z_6 ));
    InMux I__1475 (
            .O(N__10554),
            .I(N__10549));
    InMux I__1474 (
            .O(N__10553),
            .I(N__10546));
    InMux I__1473 (
            .O(N__10552),
            .I(N__10543));
    LocalMux I__1472 (
            .O(N__10549),
            .I(N__10540));
    LocalMux I__1471 (
            .O(N__10546),
            .I(N__10535));
    LocalMux I__1470 (
            .O(N__10543),
            .I(N__10535));
    Span4Mux_v I__1469 (
            .O(N__10540),
            .I(N__10532));
    Odrv4 I__1468 (
            .O(N__10535),
            .I(\uu2.N_225 ));
    Odrv4 I__1467 (
            .O(N__10532),
            .I(\uu2.N_225 ));
    CascadeMux I__1466 (
            .O(N__10527),
            .I(\uu2.N_144_cascade_ ));
    InMux I__1465 (
            .O(N__10524),
            .I(N__10521));
    LocalMux I__1464 (
            .O(N__10521),
            .I(\uu2.bitmapZ0Z_40 ));
    CascadeMux I__1463 (
            .O(N__10518),
            .I(\uu2.bitmap_RNI1PH82Z0Z_40_cascade_ ));
    CascadeMux I__1462 (
            .O(N__10515),
            .I(\uu2.N_401_cascade_ ));
    InMux I__1461 (
            .O(N__10512),
            .I(N__10509));
    LocalMux I__1460 (
            .O(N__10509),
            .I(\uu2.N_406 ));
    InMux I__1459 (
            .O(N__10506),
            .I(N__10503));
    LocalMux I__1458 (
            .O(N__10503),
            .I(N__10500));
    Odrv4 I__1457 (
            .O(N__10500),
            .I(\uu2.un31_w_data_displaying_1 ));
    CascadeMux I__1456 (
            .O(N__10497),
            .I(N__10494));
    InMux I__1455 (
            .O(N__10494),
            .I(N__10490));
    InMux I__1454 (
            .O(N__10493),
            .I(N__10487));
    LocalMux I__1453 (
            .O(N__10490),
            .I(N__10484));
    LocalMux I__1452 (
            .O(N__10487),
            .I(\uu2.un49_w_data_displaying_1 ));
    Odrv4 I__1451 (
            .O(N__10484),
            .I(\uu2.un49_w_data_displaying_1 ));
    CascadeMux I__1450 (
            .O(N__10479),
            .I(N__10476));
    InMux I__1449 (
            .O(N__10476),
            .I(N__10473));
    LocalMux I__1448 (
            .O(N__10473),
            .I(N__10470));
    Odrv4 I__1447 (
            .O(N__10470),
            .I(\uu2.mem0.N_81_i ));
    CascadeMux I__1446 (
            .O(N__10467),
            .I(N__10464));
    InMux I__1445 (
            .O(N__10464),
            .I(N__10461));
    LocalMux I__1444 (
            .O(N__10461),
            .I(N__10458));
    Span4Mux_v I__1443 (
            .O(N__10458),
            .I(N__10455));
    Odrv4 I__1442 (
            .O(N__10455),
            .I(\uu2.mem0.N_80_i ));
    InMux I__1441 (
            .O(N__10452),
            .I(N__10449));
    LocalMux I__1440 (
            .O(N__10449),
            .I(N__10446));
    Span4Mux_v I__1439 (
            .O(N__10446),
            .I(N__10443));
    Odrv4 I__1438 (
            .O(N__10443),
            .I(\uu2.mem0.N_72_i ));
    CascadeMux I__1437 (
            .O(N__10440),
            .I(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ));
    CascadeMux I__1436 (
            .O(N__10437),
            .I(\uu2.bitmap_pmux_sn_i5_mux_cascade_ ));
    InMux I__1435 (
            .O(N__10434),
            .I(N__10431));
    LocalMux I__1434 (
            .O(N__10431),
            .I(N__10428));
    Odrv12 I__1433 (
            .O(N__10428),
            .I(\uu2.N_404 ));
    CascadeMux I__1432 (
            .O(N__10425),
            .I(\uu2.bitmap_pmux_29_0_cascade_ ));
    InMux I__1431 (
            .O(N__10422),
            .I(N__10416));
    InMux I__1430 (
            .O(N__10421),
            .I(N__10416));
    LocalMux I__1429 (
            .O(N__10416),
            .I(\uu2.bitmap_pmux ));
    InMux I__1428 (
            .O(N__10413),
            .I(N__10410));
    LocalMux I__1427 (
            .O(N__10410),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__1426 (
            .O(N__10407),
            .I(N__10404));
    LocalMux I__1425 (
            .O(N__10404),
            .I(\uu2.bitmapZ0Z_52 ));
    CascadeMux I__1424 (
            .O(N__10401),
            .I(N__10393));
    CascadeMux I__1423 (
            .O(N__10400),
            .I(N__10390));
    InMux I__1422 (
            .O(N__10399),
            .I(N__10376));
    InMux I__1421 (
            .O(N__10398),
            .I(N__10376));
    InMux I__1420 (
            .O(N__10397),
            .I(N__10376));
    InMux I__1419 (
            .O(N__10396),
            .I(N__10376));
    InMux I__1418 (
            .O(N__10393),
            .I(N__10376));
    InMux I__1417 (
            .O(N__10390),
            .I(N__10376));
    InMux I__1416 (
            .O(N__10389),
            .I(N__10373));
    LocalMux I__1415 (
            .O(N__10376),
            .I(N__10370));
    LocalMux I__1414 (
            .O(N__10373),
            .I(N__10367));
    Odrv4 I__1413 (
            .O(N__10370),
            .I(\Lab_UT.sec1_3 ));
    Odrv12 I__1412 (
            .O(N__10367),
            .I(\Lab_UT.sec1_3 ));
    InMux I__1411 (
            .O(N__10362),
            .I(N__10359));
    LocalMux I__1410 (
            .O(N__10359),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__1409 (
            .O(N__10356),
            .I(N__10353));
    LocalMux I__1408 (
            .O(N__10353),
            .I(\uu2.bitmapZ0Z_84 ));
    InMux I__1407 (
            .O(N__10350),
            .I(N__10347));
    LocalMux I__1406 (
            .O(N__10347),
            .I(\uu2.bitmap_pmux_24_i_m2_am_1 ));
    CascadeMux I__1405 (
            .O(N__10344),
            .I(\uu2.un51_w_data_displaying_cascade_ ));
    InMux I__1404 (
            .O(N__10341),
            .I(N__10338));
    LocalMux I__1403 (
            .O(N__10338),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1402 (
            .O(N__10335),
            .I(N__10331));
    InMux I__1401 (
            .O(N__10334),
            .I(N__10328));
    LocalMux I__1400 (
            .O(N__10331),
            .I(N__10325));
    LocalMux I__1399 (
            .O(N__10328),
            .I(N__10322));
    Odrv4 I__1398 (
            .O(N__10325),
            .I(\uu2.w_addr_displaying_4_1 ));
    Odrv4 I__1397 (
            .O(N__10322),
            .I(\uu2.w_addr_displaying_4_1 ));
    InMux I__1396 (
            .O(N__10317),
            .I(N__10314));
    LocalMux I__1395 (
            .O(N__10314),
            .I(\uu2.un51_w_data_displaying ));
    InMux I__1394 (
            .O(N__10311),
            .I(N__10308));
    LocalMux I__1393 (
            .O(N__10308),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1392 (
            .O(N__10305),
            .I(N__10302));
    LocalMux I__1391 (
            .O(N__10302),
            .I(\uu2.mem0.w_data_1 ));
    CascadeMux I__1390 (
            .O(N__10299),
            .I(\uu2.bitmap_RNIAE522Z0Z_93_cascade_ ));
    CascadeMux I__1389 (
            .O(N__10296),
            .I(N__10293));
    InMux I__1388 (
            .O(N__10293),
            .I(N__10290));
    LocalMux I__1387 (
            .O(N__10290),
            .I(\uu2.bitmapZ0Z_215 ));
    CascadeMux I__1386 (
            .O(N__10287),
            .I(\uu2.bitmap_RNIKL222Z0Z_212_cascade_ ));
    InMux I__1385 (
            .O(N__10284),
            .I(N__10281));
    LocalMux I__1384 (
            .O(N__10281),
            .I(\uu2.bitmap_pmux_27_ns_1 ));
    InMux I__1383 (
            .O(N__10278),
            .I(N__10275));
    LocalMux I__1382 (
            .O(N__10275),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__1381 (
            .O(N__10272),
            .I(N__10269));
    LocalMux I__1380 (
            .O(N__10269),
            .I(N__10266));
    Odrv4 I__1379 (
            .O(N__10266),
            .I(vbuf_tx_data_3));
    InMux I__1378 (
            .O(N__10263),
            .I(N__10260));
    LocalMux I__1377 (
            .O(N__10260),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1376 (
            .O(N__10257),
            .I(N__10254));
    LocalMux I__1375 (
            .O(N__10254),
            .I(N__10251));
    Odrv12 I__1374 (
            .O(N__10251),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__1373 (
            .O(N__10248),
            .I(N__10245));
    LocalMux I__1372 (
            .O(N__10245),
            .I(N__10242));
    Odrv12 I__1371 (
            .O(N__10242),
            .I(vbuf_tx_data_4));
    InMux I__1370 (
            .O(N__10239),
            .I(N__10236));
    LocalMux I__1369 (
            .O(N__10236),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    CEMux I__1368 (
            .O(N__10233),
            .I(N__10230));
    LocalMux I__1367 (
            .O(N__10230),
            .I(N__10226));
    CEMux I__1366 (
            .O(N__10229),
            .I(N__10223));
    Odrv4 I__1365 (
            .O(N__10226),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    LocalMux I__1364 (
            .O(N__10223),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__1363 (
            .O(N__10218),
            .I(N__10215));
    LocalMux I__1362 (
            .O(N__10215),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__1361 (
            .O(N__10212),
            .I(N__10209));
    InMux I__1360 (
            .O(N__10209),
            .I(N__10206));
    LocalMux I__1359 (
            .O(N__10206),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__1358 (
            .O(N__10203),
            .I(N__10199));
    InMux I__1357 (
            .O(N__10202),
            .I(N__10196));
    InMux I__1356 (
            .O(N__10199),
            .I(N__10193));
    LocalMux I__1355 (
            .O(N__10196),
            .I(N__10190));
    LocalMux I__1354 (
            .O(N__10193),
            .I(\uu0.l_countZ0Z_13 ));
    Odrv4 I__1353 (
            .O(N__10190),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__1352 (
            .O(N__10185),
            .I(N__10179));
    InMux I__1351 (
            .O(N__10184),
            .I(N__10172));
    InMux I__1350 (
            .O(N__10183),
            .I(N__10172));
    InMux I__1349 (
            .O(N__10182),
            .I(N__10172));
    LocalMux I__1348 (
            .O(N__10179),
            .I(N__10169));
    LocalMux I__1347 (
            .O(N__10172),
            .I(\uu0.un4_l_count_0_8 ));
    Odrv4 I__1346 (
            .O(N__10169),
            .I(\uu0.un4_l_count_0_8 ));
    InMux I__1345 (
            .O(N__10164),
            .I(N__10157));
    InMux I__1344 (
            .O(N__10163),
            .I(N__10157));
    InMux I__1343 (
            .O(N__10162),
            .I(N__10154));
    LocalMux I__1342 (
            .O(N__10157),
            .I(N__10151));
    LocalMux I__1341 (
            .O(N__10154),
            .I(\uu0.l_countZ0Z_12 ));
    Odrv4 I__1340 (
            .O(N__10151),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__1339 (
            .O(N__10146),
            .I(N__10141));
    CascadeMux I__1338 (
            .O(N__10145),
            .I(N__10137));
    CascadeMux I__1337 (
            .O(N__10144),
            .I(N__10134));
    LocalMux I__1336 (
            .O(N__10141),
            .I(N__10131));
    InMux I__1335 (
            .O(N__10140),
            .I(N__10128));
    InMux I__1334 (
            .O(N__10137),
            .I(N__10123));
    InMux I__1333 (
            .O(N__10134),
            .I(N__10123));
    Odrv4 I__1332 (
            .O(N__10131),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__1331 (
            .O(N__10128),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__1330 (
            .O(N__10123),
            .I(\uu0.un154_ci_9 ));
    InMux I__1329 (
            .O(N__10116),
            .I(N__10113));
    LocalMux I__1328 (
            .O(N__10113),
            .I(N__10110));
    Odrv4 I__1327 (
            .O(N__10110),
            .I(\uu0.un165_ci_0 ));
    InMux I__1326 (
            .O(N__10107),
            .I(N__10104));
    LocalMux I__1325 (
            .O(N__10104),
            .I(N__10101));
    Odrv4 I__1324 (
            .O(N__10101),
            .I(vbuf_tx_data_0));
    InMux I__1323 (
            .O(N__10098),
            .I(N__10095));
    LocalMux I__1322 (
            .O(N__10095),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1321 (
            .O(N__10092),
            .I(N__10089));
    LocalMux I__1320 (
            .O(N__10089),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1319 (
            .O(N__10086),
            .I(N__10083));
    LocalMux I__1318 (
            .O(N__10083),
            .I(N__10080));
    Span12Mux_s1_h I__1317 (
            .O(N__10080),
            .I(N__10077));
    Odrv12 I__1316 (
            .O(N__10077),
            .I(o_serial_data_c));
    InMux I__1315 (
            .O(N__10074),
            .I(N__10071));
    LocalMux I__1314 (
            .O(N__10071),
            .I(N__10068));
    Odrv12 I__1313 (
            .O(N__10068),
            .I(vbuf_tx_data_1));
    InMux I__1312 (
            .O(N__10065),
            .I(N__10062));
    LocalMux I__1311 (
            .O(N__10062),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__1310 (
            .O(N__10059),
            .I(N__10056));
    LocalMux I__1309 (
            .O(N__10056),
            .I(N__10053));
    Odrv4 I__1308 (
            .O(N__10053),
            .I(vbuf_tx_data_2));
    InMux I__1307 (
            .O(N__10050),
            .I(N__10047));
    LocalMux I__1306 (
            .O(N__10047),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__1305 (
            .O(N__10044),
            .I(N__10041));
    LocalMux I__1304 (
            .O(N__10041),
            .I(N__10038));
    Sp12to4 I__1303 (
            .O(N__10038),
            .I(N__10035));
    Odrv12 I__1302 (
            .O(N__10035),
            .I(\uu2.r_data_wire_1 ));
    InMux I__1301 (
            .O(N__10032),
            .I(N__10029));
    LocalMux I__1300 (
            .O(N__10029),
            .I(N__10026));
    Span4Mux_v I__1299 (
            .O(N__10026),
            .I(N__10023));
    Odrv4 I__1298 (
            .O(N__10023),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1297 (
            .O(N__10020),
            .I(N__10017));
    LocalMux I__1296 (
            .O(N__10017),
            .I(N__10014));
    Span4Mux_v I__1295 (
            .O(N__10014),
            .I(N__10011));
    Odrv4 I__1294 (
            .O(N__10011),
            .I(\uu2.r_data_wire_3 ));
    InMux I__1293 (
            .O(N__10008),
            .I(N__10005));
    LocalMux I__1292 (
            .O(N__10005),
            .I(N__10002));
    Span4Mux_v I__1291 (
            .O(N__10002),
            .I(N__9999));
    Odrv4 I__1290 (
            .O(N__9999),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1289 (
            .O(N__9996),
            .I(N__9993));
    LocalMux I__1288 (
            .O(N__9993),
            .I(N__9990));
    Span4Mux_v I__1287 (
            .O(N__9990),
            .I(N__9987));
    Odrv4 I__1286 (
            .O(N__9987),
            .I(\uu2.r_data_wire_5 ));
    InMux I__1285 (
            .O(N__9984),
            .I(N__9981));
    LocalMux I__1284 (
            .O(N__9981),
            .I(vbuf_tx_data_5));
    InMux I__1283 (
            .O(N__9978),
            .I(N__9975));
    LocalMux I__1282 (
            .O(N__9975),
            .I(N__9972));
    Span4Mux_v I__1281 (
            .O(N__9972),
            .I(N__9969));
    Odrv4 I__1280 (
            .O(N__9969),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1279 (
            .O(N__9966),
            .I(N__9963));
    LocalMux I__1278 (
            .O(N__9963),
            .I(vbuf_tx_data_6));
    InMux I__1277 (
            .O(N__9960),
            .I(N__9957));
    LocalMux I__1276 (
            .O(N__9957),
            .I(N__9954));
    Span12Mux_s2_h I__1275 (
            .O(N__9954),
            .I(N__9951));
    Odrv12 I__1274 (
            .O(N__9951),
            .I(\uu2.r_data_wire_7 ));
    InMux I__1273 (
            .O(N__9948),
            .I(N__9945));
    LocalMux I__1272 (
            .O(N__9945),
            .I(vbuf_tx_data_7));
    CascadeMux I__1271 (
            .O(N__9942),
            .I(N__9938));
    InMux I__1270 (
            .O(N__9941),
            .I(N__9935));
    InMux I__1269 (
            .O(N__9938),
            .I(N__9932));
    LocalMux I__1268 (
            .O(N__9935),
            .I(N__9929));
    LocalMux I__1267 (
            .O(N__9932),
            .I(N__9923));
    Span12Mux_s5_v I__1266 (
            .O(N__9929),
            .I(N__9920));
    InMux I__1265 (
            .O(N__9928),
            .I(N__9917));
    InMux I__1264 (
            .O(N__9927),
            .I(N__9912));
    InMux I__1263 (
            .O(N__9926),
            .I(N__9912));
    Odrv4 I__1262 (
            .O(N__9923),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv12 I__1261 (
            .O(N__9920),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1260 (
            .O(N__9917),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1259 (
            .O(N__9912),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__1258 (
            .O(N__9903),
            .I(N__9900));
    LocalMux I__1257 (
            .O(N__9900),
            .I(N__9894));
    InMux I__1256 (
            .O(N__9899),
            .I(N__9891));
    InMux I__1255 (
            .O(N__9898),
            .I(N__9886));
    InMux I__1254 (
            .O(N__9897),
            .I(N__9886));
    Odrv12 I__1253 (
            .O(N__9894),
            .I(\uu2.un404_ci ));
    LocalMux I__1252 (
            .O(N__9891),
            .I(\uu2.un404_ci ));
    LocalMux I__1251 (
            .O(N__9886),
            .I(\uu2.un404_ci ));
    InMux I__1250 (
            .O(N__9879),
            .I(N__9876));
    LocalMux I__1249 (
            .O(N__9876),
            .I(N__9869));
    InMux I__1248 (
            .O(N__9875),
            .I(N__9860));
    InMux I__1247 (
            .O(N__9874),
            .I(N__9860));
    InMux I__1246 (
            .O(N__9873),
            .I(N__9860));
    InMux I__1245 (
            .O(N__9872),
            .I(N__9860));
    Odrv12 I__1244 (
            .O(N__9869),
            .I(\uu2.trig_rd_is_det ));
    LocalMux I__1243 (
            .O(N__9860),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__1242 (
            .O(N__9855),
            .I(N__9851));
    InMux I__1241 (
            .O(N__9854),
            .I(N__9848));
    InMux I__1240 (
            .O(N__9851),
            .I(N__9845));
    LocalMux I__1239 (
            .O(N__9848),
            .I(N__9841));
    LocalMux I__1238 (
            .O(N__9845),
            .I(N__9838));
    CascadeMux I__1237 (
            .O(N__9844),
            .I(N__9834));
    Span4Mux_v I__1236 (
            .O(N__9841),
            .I(N__9829));
    Span4Mux_h I__1235 (
            .O(N__9838),
            .I(N__9829));
    InMux I__1234 (
            .O(N__9837),
            .I(N__9826));
    InMux I__1233 (
            .O(N__9834),
            .I(N__9823));
    Span4Mux_v I__1232 (
            .O(N__9829),
            .I(N__9820));
    LocalMux I__1231 (
            .O(N__9826),
            .I(N__9817));
    LocalMux I__1230 (
            .O(N__9823),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__1229 (
            .O(N__9820),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv12 I__1228 (
            .O(N__9817),
            .I(\uu2.r_addrZ0Z_5 ));
    CEMux I__1227 (
            .O(N__9810),
            .I(N__9807));
    LocalMux I__1226 (
            .O(N__9807),
            .I(N__9804));
    Span4Mux_v I__1225 (
            .O(N__9804),
            .I(N__9801));
    Odrv4 I__1224 (
            .O(N__9801),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    InMux I__1223 (
            .O(N__9798),
            .I(N__9795));
    LocalMux I__1222 (
            .O(N__9795),
            .I(N__9788));
    InMux I__1221 (
            .O(N__9794),
            .I(N__9779));
    InMux I__1220 (
            .O(N__9793),
            .I(N__9779));
    InMux I__1219 (
            .O(N__9792),
            .I(N__9779));
    InMux I__1218 (
            .O(N__9791),
            .I(N__9779));
    Odrv4 I__1217 (
            .O(N__9788),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1216 (
            .O(N__9779),
            .I(\uu2.w_addr_userZ0Z_2 ));
    CascadeMux I__1215 (
            .O(N__9774),
            .I(\uu2.N_115_cascade_ ));
    InMux I__1214 (
            .O(N__9771),
            .I(N__9765));
    CascadeMux I__1213 (
            .O(N__9770),
            .I(N__9761));
    InMux I__1212 (
            .O(N__9769),
            .I(N__9756));
    InMux I__1211 (
            .O(N__9768),
            .I(N__9756));
    LocalMux I__1210 (
            .O(N__9765),
            .I(N__9753));
    InMux I__1209 (
            .O(N__9764),
            .I(N__9748));
    InMux I__1208 (
            .O(N__9761),
            .I(N__9748));
    LocalMux I__1207 (
            .O(N__9756),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv12 I__1206 (
            .O(N__9753),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__1205 (
            .O(N__9748),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CEMux I__1204 (
            .O(N__9741),
            .I(N__9738));
    LocalMux I__1203 (
            .O(N__9738),
            .I(N__9735));
    Span4Mux_v I__1202 (
            .O(N__9735),
            .I(N__9731));
    CEMux I__1201 (
            .O(N__9734),
            .I(N__9728));
    Span4Mux_s1_h I__1200 (
            .O(N__9731),
            .I(N__9725));
    LocalMux I__1199 (
            .O(N__9728),
            .I(N__9722));
    Odrv4 I__1198 (
            .O(N__9725),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    Odrv12 I__1197 (
            .O(N__9722),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    InMux I__1196 (
            .O(N__9717),
            .I(N__9714));
    LocalMux I__1195 (
            .O(N__9714),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__1194 (
            .O(N__9711),
            .I(N__9708));
    LocalMux I__1193 (
            .O(N__9708),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__1192 (
            .O(N__9705),
            .I(N__9701));
    InMux I__1191 (
            .O(N__9704),
            .I(N__9696));
    InMux I__1190 (
            .O(N__9701),
            .I(N__9689));
    InMux I__1189 (
            .O(N__9700),
            .I(N__9689));
    InMux I__1188 (
            .O(N__9699),
            .I(N__9689));
    LocalMux I__1187 (
            .O(N__9696),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1186 (
            .O(N__9689),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__1185 (
            .O(N__9684),
            .I(N__9681));
    InMux I__1184 (
            .O(N__9681),
            .I(N__9678));
    LocalMux I__1183 (
            .O(N__9678),
            .I(N__9675));
    Span4Mux_h I__1182 (
            .O(N__9675),
            .I(N__9672));
    Span4Mux_v I__1181 (
            .O(N__9672),
            .I(N__9669));
    Odrv4 I__1180 (
            .O(N__9669),
            .I(\uu2.mem0.N_78_i ));
    CascadeMux I__1179 (
            .O(N__9666),
            .I(N__9663));
    InMux I__1178 (
            .O(N__9663),
            .I(N__9660));
    LocalMux I__1177 (
            .O(N__9660),
            .I(N__9657));
    Span4Mux_v I__1176 (
            .O(N__9657),
            .I(N__9654));
    Odrv4 I__1175 (
            .O(N__9654),
            .I(\uu2.mem0.N_77_i ));
    InMux I__1174 (
            .O(N__9651),
            .I(N__9648));
    LocalMux I__1173 (
            .O(N__9648),
            .I(N__9645));
    Sp12to4 I__1172 (
            .O(N__9645),
            .I(N__9642));
    Odrv12 I__1171 (
            .O(N__9642),
            .I(\uu2.r_data_wire_0 ));
    CascadeMux I__1170 (
            .O(N__9639),
            .I(N__9636));
    InMux I__1169 (
            .O(N__9636),
            .I(N__9633));
    LocalMux I__1168 (
            .O(N__9633),
            .I(N__9630));
    Span4Mux_v I__1167 (
            .O(N__9630),
            .I(N__9627));
    Odrv4 I__1166 (
            .O(N__9627),
            .I(\uu2.mem0.N_75_i ));
    CascadeMux I__1165 (
            .O(N__9624),
            .I(N__9621));
    InMux I__1164 (
            .O(N__9621),
            .I(N__9618));
    LocalMux I__1163 (
            .O(N__9618),
            .I(N__9615));
    Span4Mux_v I__1162 (
            .O(N__9615),
            .I(N__9612));
    Odrv4 I__1161 (
            .O(N__9612),
            .I(\uu2.mem0.N_74_i ));
    CascadeMux I__1160 (
            .O(N__9609),
            .I(N__9605));
    InMux I__1159 (
            .O(N__9608),
            .I(N__9600));
    InMux I__1158 (
            .O(N__9605),
            .I(N__9595));
    InMux I__1157 (
            .O(N__9604),
            .I(N__9595));
    InMux I__1156 (
            .O(N__9603),
            .I(N__9592));
    LocalMux I__1155 (
            .O(N__9600),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1154 (
            .O(N__9595),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__1153 (
            .O(N__9592),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__1152 (
            .O(N__9585),
            .I(N__9581));
    InMux I__1151 (
            .O(N__9584),
            .I(N__9577));
    LocalMux I__1150 (
            .O(N__9581),
            .I(N__9574));
    InMux I__1149 (
            .O(N__9580),
            .I(N__9571));
    LocalMux I__1148 (
            .O(N__9577),
            .I(\uu2.w_addr_userZ0Z_8 ));
    Odrv4 I__1147 (
            .O(N__9574),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__1146 (
            .O(N__9571),
            .I(\uu2.w_addr_userZ0Z_8 ));
    InMux I__1145 (
            .O(N__9564),
            .I(N__9561));
    LocalMux I__1144 (
            .O(N__9561),
            .I(\uu2.N_186 ));
    InMux I__1143 (
            .O(N__9558),
            .I(N__9555));
    LocalMux I__1142 (
            .O(N__9555),
            .I(\uu2.w_addr_user_3_i_a2_2_6 ));
    CascadeMux I__1141 (
            .O(N__9552),
            .I(\uu2.N_150_cascade_ ));
    CascadeMux I__1140 (
            .O(N__9549),
            .I(N__9546));
    InMux I__1139 (
            .O(N__9546),
            .I(N__9543));
    LocalMux I__1138 (
            .O(N__9543),
            .I(N__9540));
    Odrv4 I__1137 (
            .O(N__9540),
            .I(\uu2.mem0.N_79_i ));
    InMux I__1136 (
            .O(N__9537),
            .I(N__9533));
    InMux I__1135 (
            .O(N__9536),
            .I(N__9530));
    LocalMux I__1134 (
            .O(N__9533),
            .I(N__9527));
    LocalMux I__1133 (
            .O(N__9530),
            .I(N__9524));
    Odrv4 I__1132 (
            .O(N__9527),
            .I(\uu2.un1_l_count_1_0 ));
    Odrv4 I__1131 (
            .O(N__9524),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1130 (
            .O(N__9519),
            .I(N__9516));
    LocalMux I__1129 (
            .O(N__9516),
            .I(\uu0.sec_clkDZ0 ));
    CascadeMux I__1128 (
            .O(N__9513),
            .I(oneSecStrb_cascade_));
    CascadeMux I__1127 (
            .O(N__9510),
            .I(\uu2.N_118_cascade_ ));
    InMux I__1126 (
            .O(N__9507),
            .I(N__9504));
    LocalMux I__1125 (
            .O(N__9504),
            .I(\uu2.N_117 ));
    CascadeMux I__1124 (
            .O(N__9501),
            .I(\uu2.N_117_cascade_ ));
    CascadeMux I__1123 (
            .O(N__9498),
            .I(\uu2.un404_ci_cascade_ ));
    InMux I__1122 (
            .O(N__9495),
            .I(N__9492));
    LocalMux I__1121 (
            .O(N__9492),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__1120 (
            .O(N__9489),
            .I(N__9486));
    InMux I__1119 (
            .O(N__9486),
            .I(N__9481));
    InMux I__1118 (
            .O(N__9485),
            .I(N__9476));
    InMux I__1117 (
            .O(N__9484),
            .I(N__9476));
    LocalMux I__1116 (
            .O(N__9481),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1115 (
            .O(N__9476),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__1114 (
            .O(N__9471),
            .I(N__9468));
    LocalMux I__1113 (
            .O(N__9468),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    CascadeMux I__1112 (
            .O(N__9465),
            .I(N__9461));
    CascadeMux I__1111 (
            .O(N__9464),
            .I(N__9457));
    InMux I__1110 (
            .O(N__9461),
            .I(N__9453));
    InMux I__1109 (
            .O(N__9460),
            .I(N__9450));
    InMux I__1108 (
            .O(N__9457),
            .I(N__9445));
    InMux I__1107 (
            .O(N__9456),
            .I(N__9445));
    LocalMux I__1106 (
            .O(N__9453),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1105 (
            .O(N__9450),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1104 (
            .O(N__9445),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__1103 (
            .O(N__9438),
            .I(N__9435));
    InMux I__1102 (
            .O(N__9435),
            .I(N__9431));
    CascadeMux I__1101 (
            .O(N__9434),
            .I(N__9428));
    LocalMux I__1100 (
            .O(N__9431),
            .I(N__9425));
    InMux I__1099 (
            .O(N__9428),
            .I(N__9420));
    Span4Mux_h I__1098 (
            .O(N__9425),
            .I(N__9417));
    InMux I__1097 (
            .O(N__9424),
            .I(N__9412));
    InMux I__1096 (
            .O(N__9423),
            .I(N__9412));
    LocalMux I__1095 (
            .O(N__9420),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__1094 (
            .O(N__9417),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1093 (
            .O(N__9412),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1092 (
            .O(N__9405),
            .I(N__9402));
    InMux I__1091 (
            .O(N__9402),
            .I(N__9399));
    LocalMux I__1090 (
            .O(N__9399),
            .I(N__9392));
    InMux I__1089 (
            .O(N__9398),
            .I(N__9387));
    InMux I__1088 (
            .O(N__9397),
            .I(N__9387));
    InMux I__1087 (
            .O(N__9396),
            .I(N__9382));
    InMux I__1086 (
            .O(N__9395),
            .I(N__9382));
    Odrv4 I__1085 (
            .O(N__9392),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1084 (
            .O(N__9387),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__1083 (
            .O(N__9382),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1082 (
            .O(N__9375),
            .I(N__9372));
    InMux I__1081 (
            .O(N__9372),
            .I(N__9368));
    CascadeMux I__1080 (
            .O(N__9371),
            .I(N__9364));
    LocalMux I__1079 (
            .O(N__9368),
            .I(N__9358));
    InMux I__1078 (
            .O(N__9367),
            .I(N__9351));
    InMux I__1077 (
            .O(N__9364),
            .I(N__9351));
    InMux I__1076 (
            .O(N__9363),
            .I(N__9351));
    InMux I__1075 (
            .O(N__9362),
            .I(N__9346));
    InMux I__1074 (
            .O(N__9361),
            .I(N__9346));
    Odrv4 I__1073 (
            .O(N__9358),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1072 (
            .O(N__9351),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1071 (
            .O(N__9346),
            .I(\uu2.r_addrZ0Z_0 ));
    CascadeMux I__1070 (
            .O(N__9339),
            .I(N__9334));
    CascadeMux I__1069 (
            .O(N__9338),
            .I(N__9331));
    CascadeMux I__1068 (
            .O(N__9337),
            .I(N__9328));
    InMux I__1067 (
            .O(N__9334),
            .I(N__9325));
    InMux I__1066 (
            .O(N__9331),
            .I(N__9320));
    InMux I__1065 (
            .O(N__9328),
            .I(N__9320));
    LocalMux I__1064 (
            .O(N__9325),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1063 (
            .O(N__9320),
            .I(\uu2.r_addrZ0Z_3 ));
    CEMux I__1062 (
            .O(N__9315),
            .I(N__9312));
    LocalMux I__1061 (
            .O(N__9312),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__1060 (
            .O(N__9309),
            .I(N__9306));
    InMux I__1059 (
            .O(N__9306),
            .I(N__9303));
    LocalMux I__1058 (
            .O(N__9303),
            .I(\uu2.mem0.N_76_i ));
    CascadeMux I__1057 (
            .O(N__9300),
            .I(N__9297));
    InMux I__1056 (
            .O(N__9297),
            .I(N__9294));
    LocalMux I__1055 (
            .O(N__9294),
            .I(N__9291));
    Odrv4 I__1054 (
            .O(N__9291),
            .I(\uu2.mem0.N_73_i ));
    CascadeMux I__1053 (
            .O(N__9288),
            .I(N__9282));
    InMux I__1052 (
            .O(N__9287),
            .I(N__9275));
    InMux I__1051 (
            .O(N__9286),
            .I(N__9272));
    InMux I__1050 (
            .O(N__9285),
            .I(N__9269));
    InMux I__1049 (
            .O(N__9282),
            .I(N__9262));
    InMux I__1048 (
            .O(N__9281),
            .I(N__9262));
    InMux I__1047 (
            .O(N__9280),
            .I(N__9262));
    CascadeMux I__1046 (
            .O(N__9279),
            .I(N__9258));
    CascadeMux I__1045 (
            .O(N__9278),
            .I(N__9255));
    LocalMux I__1044 (
            .O(N__9275),
            .I(N__9245));
    LocalMux I__1043 (
            .O(N__9272),
            .I(N__9245));
    LocalMux I__1042 (
            .O(N__9269),
            .I(N__9245));
    LocalMux I__1041 (
            .O(N__9262),
            .I(N__9245));
    InMux I__1040 (
            .O(N__9261),
            .I(N__9236));
    InMux I__1039 (
            .O(N__9258),
            .I(N__9236));
    InMux I__1038 (
            .O(N__9255),
            .I(N__9236));
    InMux I__1037 (
            .O(N__9254),
            .I(N__9236));
    Odrv12 I__1036 (
            .O(N__9245),
            .I(\uu0.un110_ci ));
    LocalMux I__1035 (
            .O(N__9236),
            .I(\uu0.un110_ci ));
    CEMux I__1034 (
            .O(N__9231),
            .I(N__9213));
    CEMux I__1033 (
            .O(N__9230),
            .I(N__9213));
    CEMux I__1032 (
            .O(N__9229),
            .I(N__9213));
    CEMux I__1031 (
            .O(N__9228),
            .I(N__9213));
    CEMux I__1030 (
            .O(N__9227),
            .I(N__9213));
    CEMux I__1029 (
            .O(N__9226),
            .I(N__9213));
    GlobalMux I__1028 (
            .O(N__9213),
            .I(N__9210));
    gio2CtrlBuf I__1027 (
            .O(N__9210),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__1026 (
            .O(N__9207),
            .I(\uu2.trig_rd_is_det_cascade_ ));
    InMux I__1025 (
            .O(N__9204),
            .I(N__9198));
    InMux I__1024 (
            .O(N__9203),
            .I(N__9198));
    LocalMux I__1023 (
            .O(N__9198),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    InMux I__1022 (
            .O(N__9195),
            .I(N__9192));
    LocalMux I__1021 (
            .O(N__9192),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    CascadeMux I__1020 (
            .O(N__9189),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1019 (
            .O(N__9186),
            .I(N__9183));
    InMux I__1018 (
            .O(N__9183),
            .I(N__9179));
    InMux I__1017 (
            .O(N__9182),
            .I(N__9176));
    LocalMux I__1016 (
            .O(N__9179),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1015 (
            .O(N__9176),
            .I(\uu2.r_addrZ0Z_8 ));
    InMux I__1014 (
            .O(N__9171),
            .I(N__9166));
    InMux I__1013 (
            .O(N__9170),
            .I(N__9163));
    InMux I__1012 (
            .O(N__9169),
            .I(N__9160));
    LocalMux I__1011 (
            .O(N__9166),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__1010 (
            .O(N__9163),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__1009 (
            .O(N__9160),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__1008 (
            .O(N__9153),
            .I(\uu0.un154_ci_9_cascade_ ));
    CascadeMux I__1007 (
            .O(N__9150),
            .I(\uu0.un187_ci_1_cascade_ ));
    CascadeMux I__1006 (
            .O(N__9147),
            .I(N__9143));
    InMux I__1005 (
            .O(N__9146),
            .I(N__9140));
    InMux I__1004 (
            .O(N__9143),
            .I(N__9137));
    LocalMux I__1003 (
            .O(N__9140),
            .I(N__9129));
    LocalMux I__1002 (
            .O(N__9137),
            .I(N__9129));
    InMux I__1001 (
            .O(N__9136),
            .I(N__9122));
    InMux I__1000 (
            .O(N__9135),
            .I(N__9122));
    InMux I__999 (
            .O(N__9134),
            .I(N__9122));
    Odrv12 I__998 (
            .O(N__9129),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__997 (
            .O(N__9122),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__996 (
            .O(N__9117),
            .I(N__9105));
    InMux I__995 (
            .O(N__9116),
            .I(N__9105));
    InMux I__994 (
            .O(N__9115),
            .I(N__9105));
    InMux I__993 (
            .O(N__9114),
            .I(N__9105));
    LocalMux I__992 (
            .O(N__9105),
            .I(\uu0.l_countZ0Z_14 ));
    InMux I__991 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__990 (
            .O(N__9099),
            .I(N__9093));
    InMux I__989 (
            .O(N__9098),
            .I(N__9088));
    InMux I__988 (
            .O(N__9097),
            .I(N__9088));
    InMux I__987 (
            .O(N__9096),
            .I(N__9085));
    Odrv4 I__986 (
            .O(N__9093),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__985 (
            .O(N__9088),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__984 (
            .O(N__9085),
            .I(\uu0.l_countZ0Z_10 ));
    CascadeMux I__983 (
            .O(N__9078),
            .I(N__9073));
    InMux I__982 (
            .O(N__9077),
            .I(N__9070));
    InMux I__981 (
            .O(N__9076),
            .I(N__9065));
    InMux I__980 (
            .O(N__9073),
            .I(N__9065));
    LocalMux I__979 (
            .O(N__9070),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__978 (
            .O(N__9065),
            .I(\uu0.l_countZ0Z_15 ));
    InMux I__977 (
            .O(N__9060),
            .I(N__9057));
    LocalMux I__976 (
            .O(N__9057),
            .I(\uu0.un4_l_count_13 ));
    InMux I__975 (
            .O(N__9054),
            .I(N__9051));
    LocalMux I__974 (
            .O(N__9051),
            .I(N__9046));
    InMux I__973 (
            .O(N__9050),
            .I(N__9043));
    CascadeMux I__972 (
            .O(N__9049),
            .I(N__9039));
    Span4Mux_s2_v I__971 (
            .O(N__9046),
            .I(N__9034));
    LocalMux I__970 (
            .O(N__9043),
            .I(N__9034));
    InMux I__969 (
            .O(N__9042),
            .I(N__9031));
    InMux I__968 (
            .O(N__9039),
            .I(N__9028));
    Odrv4 I__967 (
            .O(N__9034),
            .I(\uu0.un66_ci ));
    LocalMux I__966 (
            .O(N__9031),
            .I(\uu0.un66_ci ));
    LocalMux I__965 (
            .O(N__9028),
            .I(\uu0.un66_ci ));
    InMux I__964 (
            .O(N__9021),
            .I(N__9017));
    InMux I__963 (
            .O(N__9020),
            .I(N__9012));
    LocalMux I__962 (
            .O(N__9017),
            .I(N__9009));
    InMux I__961 (
            .O(N__9016),
            .I(N__9004));
    InMux I__960 (
            .O(N__9015),
            .I(N__9004));
    LocalMux I__959 (
            .O(N__9012),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv12 I__958 (
            .O(N__9009),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__957 (
            .O(N__9004),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__956 (
            .O(N__8997),
            .I(N__8994));
    LocalMux I__955 (
            .O(N__8994),
            .I(N__8990));
    InMux I__954 (
            .O(N__8993),
            .I(N__8987));
    Span4Mux_v I__953 (
            .O(N__8990),
            .I(N__8981));
    LocalMux I__952 (
            .O(N__8987),
            .I(N__8981));
    InMux I__951 (
            .O(N__8986),
            .I(N__8978));
    Span4Mux_v I__950 (
            .O(N__8981),
            .I(N__8975));
    LocalMux I__949 (
            .O(N__8978),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv4 I__948 (
            .O(N__8975),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__947 (
            .O(N__8970),
            .I(N__8967));
    InMux I__946 (
            .O(N__8967),
            .I(N__8958));
    InMux I__945 (
            .O(N__8966),
            .I(N__8958));
    InMux I__944 (
            .O(N__8965),
            .I(N__8954));
    InMux I__943 (
            .O(N__8964),
            .I(N__8951));
    InMux I__942 (
            .O(N__8963),
            .I(N__8948));
    LocalMux I__941 (
            .O(N__8958),
            .I(N__8945));
    InMux I__940 (
            .O(N__8957),
            .I(N__8942));
    LocalMux I__939 (
            .O(N__8954),
            .I(N__8939));
    LocalMux I__938 (
            .O(N__8951),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__937 (
            .O(N__8948),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv4 I__936 (
            .O(N__8945),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__935 (
            .O(N__8942),
            .I(\uu0.l_countZ0Z_8 ));
    Odrv12 I__934 (
            .O(N__8939),
            .I(\uu0.l_countZ0Z_8 ));
    InMux I__933 (
            .O(N__8928),
            .I(N__8922));
    InMux I__932 (
            .O(N__8927),
            .I(N__8915));
    InMux I__931 (
            .O(N__8926),
            .I(N__8915));
    InMux I__930 (
            .O(N__8925),
            .I(N__8915));
    LocalMux I__929 (
            .O(N__8922),
            .I(N__8912));
    LocalMux I__928 (
            .O(N__8915),
            .I(\uu0.l_countZ0Z_16 ));
    Odrv4 I__927 (
            .O(N__8912),
            .I(\uu0.l_countZ0Z_16 ));
    InMux I__926 (
            .O(N__8907),
            .I(N__8904));
    LocalMux I__925 (
            .O(N__8904),
            .I(\uu0.un44_ci ));
    CascadeMux I__924 (
            .O(N__8901),
            .I(N__8898));
    InMux I__923 (
            .O(N__8898),
            .I(N__8895));
    LocalMux I__922 (
            .O(N__8895),
            .I(N__8889));
    InMux I__921 (
            .O(N__8894),
            .I(N__8884));
    InMux I__920 (
            .O(N__8893),
            .I(N__8884));
    InMux I__919 (
            .O(N__8892),
            .I(N__8881));
    Odrv4 I__918 (
            .O(N__8889),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__917 (
            .O(N__8884),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__916 (
            .O(N__8881),
            .I(\uu0.l_countZ0Z_2 ));
    InMux I__915 (
            .O(N__8874),
            .I(N__8869));
    InMux I__914 (
            .O(N__8873),
            .I(N__8864));
    InMux I__913 (
            .O(N__8872),
            .I(N__8864));
    LocalMux I__912 (
            .O(N__8869),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__911 (
            .O(N__8864),
            .I(\uu0.l_countZ0Z_3 ));
    CascadeMux I__910 (
            .O(N__8859),
            .I(N__8856));
    InMux I__909 (
            .O(N__8856),
            .I(N__8853));
    LocalMux I__908 (
            .O(N__8853),
            .I(N__8850));
    Odrv4 I__907 (
            .O(N__8850),
            .I(\uu0.un99_ci_0 ));
    InMux I__906 (
            .O(N__8847),
            .I(N__8842));
    InMux I__905 (
            .O(N__8846),
            .I(N__8837));
    InMux I__904 (
            .O(N__8845),
            .I(N__8837));
    LocalMux I__903 (
            .O(N__8842),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__902 (
            .O(N__8837),
            .I(\uu0.l_countZ0Z_7 ));
    InMux I__901 (
            .O(N__8832),
            .I(N__8829));
    LocalMux I__900 (
            .O(N__8829),
            .I(\uu0.un220_ci ));
    InMux I__899 (
            .O(N__8826),
            .I(N__8822));
    InMux I__898 (
            .O(N__8825),
            .I(N__8817));
    LocalMux I__897 (
            .O(N__8822),
            .I(N__8814));
    InMux I__896 (
            .O(N__8821),
            .I(N__8809));
    InMux I__895 (
            .O(N__8820),
            .I(N__8809));
    LocalMux I__894 (
            .O(N__8817),
            .I(N__8806));
    Odrv4 I__893 (
            .O(N__8814),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__892 (
            .O(N__8809),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__891 (
            .O(N__8806),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__890 (
            .O(N__8799),
            .I(N__8796));
    LocalMux I__889 (
            .O(N__8796),
            .I(\uu0.un4_l_count_11 ));
    CascadeMux I__888 (
            .O(N__8793),
            .I(N__8789));
    InMux I__887 (
            .O(N__8792),
            .I(N__8784));
    InMux I__886 (
            .O(N__8789),
            .I(N__8784));
    LocalMux I__885 (
            .O(N__8784),
            .I(\uu0.l_countZ0Z_18 ));
    InMux I__884 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__883 (
            .O(N__8778),
            .I(N__8775));
    Odrv4 I__882 (
            .O(N__8775),
            .I(\uu0.un4_l_count_18 ));
    CascadeMux I__881 (
            .O(N__8772),
            .I(\uu0.un4_l_count_16_cascade_ ));
    InMux I__880 (
            .O(N__8769),
            .I(N__8766));
    LocalMux I__879 (
            .O(N__8766),
            .I(N__8763));
    Odrv4 I__878 (
            .O(N__8763),
            .I(\uu0.un4_l_count_12 ));
    CascadeMux I__877 (
            .O(N__8760),
            .I(\uu0.un4_l_count_0_cascade_ ));
    InMux I__876 (
            .O(N__8757),
            .I(N__8754));
    LocalMux I__875 (
            .O(N__8754),
            .I(\uu0.un143_ci_0 ));
    CascadeMux I__874 (
            .O(N__8751),
            .I(N__8746));
    InMux I__873 (
            .O(N__8750),
            .I(N__8739));
    InMux I__872 (
            .O(N__8749),
            .I(N__8739));
    InMux I__871 (
            .O(N__8746),
            .I(N__8739));
    LocalMux I__870 (
            .O(N__8739),
            .I(N__8736));
    Odrv4 I__869 (
            .O(N__8736),
            .I(\uu0.un198_ci_2 ));
    InMux I__868 (
            .O(N__8733),
            .I(N__8720));
    InMux I__867 (
            .O(N__8732),
            .I(N__8720));
    InMux I__866 (
            .O(N__8731),
            .I(N__8720));
    InMux I__865 (
            .O(N__8730),
            .I(N__8720));
    InMux I__864 (
            .O(N__8729),
            .I(N__8717));
    LocalMux I__863 (
            .O(N__8720),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__862 (
            .O(N__8717),
            .I(\uu0.l_countZ0Z_0 ));
    CascadeMux I__861 (
            .O(N__8712),
            .I(N__8707));
    InMux I__860 (
            .O(N__8711),
            .I(N__8699));
    InMux I__859 (
            .O(N__8710),
            .I(N__8699));
    InMux I__858 (
            .O(N__8707),
            .I(N__8699));
    InMux I__857 (
            .O(N__8706),
            .I(N__8696));
    LocalMux I__856 (
            .O(N__8699),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__855 (
            .O(N__8696),
            .I(\uu0.l_countZ0Z_1 ));
    InMux I__854 (
            .O(N__8691),
            .I(N__8684));
    InMux I__853 (
            .O(N__8690),
            .I(N__8684));
    InMux I__852 (
            .O(N__8689),
            .I(N__8681));
    LocalMux I__851 (
            .O(N__8684),
            .I(N__8678));
    LocalMux I__850 (
            .O(N__8681),
            .I(\uu0.un88_ci_3 ));
    Odrv4 I__849 (
            .O(N__8678),
            .I(\uu0.un88_ci_3 ));
    CascadeMux I__848 (
            .O(N__8673),
            .I(\uu0.un66_ci_cascade_ ));
    CascadeMux I__847 (
            .O(N__8670),
            .I(\uu0.un110_ci_cascade_ ));
    CascadeMux I__846 (
            .O(N__8667),
            .I(N__8662));
    InMux I__845 (
            .O(N__8666),
            .I(N__8655));
    InMux I__844 (
            .O(N__8665),
            .I(N__8655));
    InMux I__843 (
            .O(N__8662),
            .I(N__8655));
    LocalMux I__842 (
            .O(N__8655),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__841 (
            .O(N__8652),
            .I(N__8647));
    CascadeMux I__840 (
            .O(N__8651),
            .I(N__8644));
    InMux I__839 (
            .O(N__8650),
            .I(N__8637));
    InMux I__838 (
            .O(N__8647),
            .I(N__8637));
    InMux I__837 (
            .O(N__8644),
            .I(N__8637));
    LocalMux I__836 (
            .O(N__8637),
            .I(\uu0.l_precountZ0Z_3 ));
    InMux I__835 (
            .O(N__8634),
            .I(N__8619));
    InMux I__834 (
            .O(N__8633),
            .I(N__8619));
    InMux I__833 (
            .O(N__8632),
            .I(N__8619));
    InMux I__832 (
            .O(N__8631),
            .I(N__8619));
    InMux I__831 (
            .O(N__8630),
            .I(N__8619));
    LocalMux I__830 (
            .O(N__8619),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__829 (
            .O(N__8616),
            .I(N__8610));
    InMux I__828 (
            .O(N__8615),
            .I(N__8601));
    InMux I__827 (
            .O(N__8614),
            .I(N__8601));
    InMux I__826 (
            .O(N__8613),
            .I(N__8601));
    InMux I__825 (
            .O(N__8610),
            .I(N__8601));
    LocalMux I__824 (
            .O(N__8601),
            .I(\uu0.l_precountZ0Z_2 ));
    CascadeMux I__823 (
            .O(N__8598),
            .I(N__8595));
    InMux I__822 (
            .O(N__8595),
            .I(N__8579));
    InMux I__821 (
            .O(N__8594),
            .I(N__8579));
    InMux I__820 (
            .O(N__8593),
            .I(N__8579));
    InMux I__819 (
            .O(N__8592),
            .I(N__8579));
    InMux I__818 (
            .O(N__8591),
            .I(N__8579));
    InMux I__817 (
            .O(N__8590),
            .I(N__8576));
    LocalMux I__816 (
            .O(N__8579),
            .I(N__8573));
    LocalMux I__815 (
            .O(N__8576),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv12 I__814 (
            .O(N__8573),
            .I(\uu0.l_precountZ0Z_0 ));
    CascadeMux I__813 (
            .O(N__8568),
            .I(\uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__812 (
            .O(N__8565),
            .I(\uu0.un44_ci_cascade_ ));
    InMux I__811 (
            .O(N__8562),
            .I(N__8557));
    CascadeMux I__810 (
            .O(N__8561),
            .I(N__8552));
    InMux I__809 (
            .O(N__8560),
            .I(N__8549));
    LocalMux I__808 (
            .O(N__8557),
            .I(N__8546));
    InMux I__807 (
            .O(N__8556),
            .I(N__8539));
    InMux I__806 (
            .O(N__8555),
            .I(N__8539));
    InMux I__805 (
            .O(N__8552),
            .I(N__8539));
    LocalMux I__804 (
            .O(N__8549),
            .I(\uu2.l_countZ0Z_1 ));
    Odrv4 I__803 (
            .O(N__8546),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__802 (
            .O(N__8539),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__801 (
            .O(N__8532),
            .I(N__8526));
    InMux I__800 (
            .O(N__8531),
            .I(N__8523));
    InMux I__799 (
            .O(N__8530),
            .I(N__8520));
    InMux I__798 (
            .O(N__8529),
            .I(N__8515));
    LocalMux I__797 (
            .O(N__8526),
            .I(N__8510));
    LocalMux I__796 (
            .O(N__8523),
            .I(N__8510));
    LocalMux I__795 (
            .O(N__8520),
            .I(N__8507));
    InMux I__794 (
            .O(N__8519),
            .I(N__8502));
    InMux I__793 (
            .O(N__8518),
            .I(N__8502));
    LocalMux I__792 (
            .O(N__8515),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv12 I__791 (
            .O(N__8510),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__790 (
            .O(N__8507),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__789 (
            .O(N__8502),
            .I(\uu2.l_countZ0Z_0 ));
    CascadeMux I__788 (
            .O(N__8493),
            .I(N__8490));
    InMux I__787 (
            .O(N__8490),
            .I(N__8484));
    InMux I__786 (
            .O(N__8489),
            .I(N__8484));
    LocalMux I__785 (
            .O(N__8484),
            .I(N__8481));
    Odrv4 I__784 (
            .O(N__8481),
            .I(\uu2.un284_ci ));
    CascadeMux I__783 (
            .O(N__8478),
            .I(N__8475));
    InMux I__782 (
            .O(N__8475),
            .I(N__8470));
    InMux I__781 (
            .O(N__8474),
            .I(N__8467));
    InMux I__780 (
            .O(N__8473),
            .I(N__8464));
    LocalMux I__779 (
            .O(N__8470),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__778 (
            .O(N__8467),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__777 (
            .O(N__8464),
            .I(\uu2.l_countZ0Z_7 ));
    CascadeMux I__776 (
            .O(N__8457),
            .I(N__8452));
    InMux I__775 (
            .O(N__8456),
            .I(N__8447));
    InMux I__774 (
            .O(N__8455),
            .I(N__8447));
    InMux I__773 (
            .O(N__8452),
            .I(N__8444));
    LocalMux I__772 (
            .O(N__8447),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__771 (
            .O(N__8444),
            .I(\uu2.l_countZ0Z_8 ));
    InMux I__770 (
            .O(N__8439),
            .I(N__8430));
    InMux I__769 (
            .O(N__8438),
            .I(N__8430));
    InMux I__768 (
            .O(N__8437),
            .I(N__8430));
    LocalMux I__767 (
            .O(N__8430),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__766 (
            .O(N__8427),
            .I(N__8424));
    InMux I__765 (
            .O(N__8424),
            .I(N__8421));
    LocalMux I__764 (
            .O(N__8421),
            .I(\uu2.un1_l_count_1_3 ));
    InMux I__763 (
            .O(N__8418),
            .I(N__8403));
    InMux I__762 (
            .O(N__8417),
            .I(N__8403));
    InMux I__761 (
            .O(N__8416),
            .I(N__8403));
    InMux I__760 (
            .O(N__8415),
            .I(N__8403));
    InMux I__759 (
            .O(N__8414),
            .I(N__8403));
    LocalMux I__758 (
            .O(N__8403),
            .I(\uu2.l_countZ0Z_2 ));
    CascadeMux I__757 (
            .O(N__8400),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    InMux I__756 (
            .O(N__8397),
            .I(N__8394));
    LocalMux I__755 (
            .O(N__8394),
            .I(\uu2.un1_l_count_2_2 ));
    InMux I__754 (
            .O(N__8391),
            .I(N__8386));
    InMux I__753 (
            .O(N__8390),
            .I(N__8383));
    InMux I__752 (
            .O(N__8389),
            .I(N__8380));
    LocalMux I__751 (
            .O(N__8386),
            .I(N__8377));
    LocalMux I__750 (
            .O(N__8383),
            .I(\uu2.un1_l_count_2_0 ));
    LocalMux I__749 (
            .O(N__8380),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__748 (
            .O(N__8377),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__747 (
            .O(N__8370),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__746 (
            .O(N__8367),
            .I(N__8358));
    InMux I__745 (
            .O(N__8366),
            .I(N__8358));
    InMux I__744 (
            .O(N__8365),
            .I(N__8351));
    InMux I__743 (
            .O(N__8364),
            .I(N__8351));
    InMux I__742 (
            .O(N__8363),
            .I(N__8351));
    LocalMux I__741 (
            .O(N__8358),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__740 (
            .O(N__8351),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__739 (
            .O(N__8346),
            .I(N__8337));
    InMux I__738 (
            .O(N__8345),
            .I(N__8337));
    InMux I__737 (
            .O(N__8344),
            .I(N__8330));
    InMux I__736 (
            .O(N__8343),
            .I(N__8330));
    InMux I__735 (
            .O(N__8342),
            .I(N__8330));
    LocalMux I__734 (
            .O(N__8337),
            .I(\uu2.un306_ci ));
    LocalMux I__733 (
            .O(N__8330),
            .I(\uu2.un306_ci ));
    CascadeMux I__732 (
            .O(N__8325),
            .I(N__8321));
    InMux I__731 (
            .O(N__8324),
            .I(N__8317));
    InMux I__730 (
            .O(N__8321),
            .I(N__8312));
    InMux I__729 (
            .O(N__8320),
            .I(N__8312));
    LocalMux I__728 (
            .O(N__8317),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__727 (
            .O(N__8312),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__726 (
            .O(N__8307),
            .I(N__8304));
    LocalMux I__725 (
            .O(N__8304),
            .I(N__8301));
    IoSpan4Mux I__724 (
            .O(N__8301),
            .I(N__8298));
    Odrv4 I__723 (
            .O(N__8298),
            .I(uart_RXD));
    CascadeMux I__722 (
            .O(N__8295),
            .I(N__8290));
    CascadeMux I__721 (
            .O(N__8294),
            .I(N__8287));
    InMux I__720 (
            .O(N__8293),
            .I(N__8280));
    InMux I__719 (
            .O(N__8290),
            .I(N__8280));
    InMux I__718 (
            .O(N__8287),
            .I(N__8280));
    LocalMux I__717 (
            .O(N__8280),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__716 (
            .O(N__8277),
            .I(N__8271));
    InMux I__715 (
            .O(N__8276),
            .I(N__8271));
    LocalMux I__714 (
            .O(N__8271),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    CascadeMux I__713 (
            .O(N__8268),
            .I(\uu2.vbuf_count.un328_ci_3_cascade_ ));
    InMux I__712 (
            .O(N__8265),
            .I(N__8250));
    InMux I__711 (
            .O(N__8264),
            .I(N__8250));
    InMux I__710 (
            .O(N__8263),
            .I(N__8250));
    InMux I__709 (
            .O(N__8262),
            .I(N__8250));
    InMux I__708 (
            .O(N__8261),
            .I(N__8250));
    LocalMux I__707 (
            .O(N__8250),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__706 (
            .O(N__8247),
            .I(N__8244));
    InMux I__705 (
            .O(N__8244),
            .I(N__8241));
    LocalMux I__704 (
            .O(N__8241),
            .I(\uu2.un350_ci ));
    CascadeMux I__703 (
            .O(N__8238),
            .I(\uu2.un350_ci_cascade_ ));
    InMux I__702 (
            .O(N__8235),
            .I(N__8232));
    LocalMux I__701 (
            .O(N__8232),
            .I(\uu2.un1_l_count_1_2_0 ));
    IoInMux I__700 (
            .O(N__8229),
            .I(N__8226));
    LocalMux I__699 (
            .O(N__8226),
            .I(N__8223));
    Span12Mux_s5_v I__698 (
            .O(N__8223),
            .I(N__8220));
    Odrv12 I__697 (
            .O(N__8220),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__696 (
            .O(N__8217),
            .I(N__8214));
    LocalMux I__695 (
            .O(N__8214),
            .I(N__8211));
    IoSpan4Mux I__694 (
            .O(N__8211),
            .I(N__8208));
    Odrv4 I__693 (
            .O(N__8208),
            .I(clk_in_c));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__22806));
    INV \INVuu2.w_addr_displaying_ness_6C  (
            .O(\INVuu2.w_addr_displaying_ness_6C_net ),
            .I(N__22814));
    INV \INVuu2.w_addr_displaying_2C  (
            .O(\INVuu2.w_addr_displaying_2C_net ),
            .I(N__22799));
    INV \INVuu2.w_addr_displaying_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .I(N__22811));
    INV \INVuu2.w_addr_displaying_8C  (
            .O(\INVuu2.w_addr_displaying_8C_net ),
            .I(N__22818));
    INV \INVuu2.bitmap_69C  (
            .O(\INVuu2.bitmap_69C_net ),
            .I(N__22822));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__22831));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__22846));
    INV \INVuu2.bitmap_40C  (
            .O(\INVuu2.bitmap_40C_net ),
            .I(N__22810));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__22830));
    INV \INVuu2.bitmap_215C  (
            .O(\INVuu2.bitmap_215C_net ),
            .I(N__22838));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__22845));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__22794));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__22802));
    INV \INVuu2.w_addr_user_nesr_7C  (
            .O(\INVuu2.w_addr_user_nesr_7C_net ),
            .I(N__22809));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_12_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_3_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__8229),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB bu_rx_data_rdy_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__22338),
            .GLOBALBUFFEROUTPUT(bu_rx_data_rdy_0_g));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__16569),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    ICE_GB \buart.Z_rx.sample_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__19218),
            .GLOBALBUFFEROUTPUT(buart__rx_sample_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__19647),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.vram_rd_clk_LC_1_3_5 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_1_3_5 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_1_3_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__12198),
            .in2(_gnd_net_),
            .in3(N__8391),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22854),
            .ce(),
            .sr(N__22516));
    defparam \uu2.l_count_0_LC_1_4_0 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_1_4_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_1_4_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8529),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22851),
            .ce(),
            .sr(N__22495));
    defparam \uu2.trig_rd_det_0_LC_1_4_1 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_1_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_1_4_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(N__12199),
            .in2(_gnd_net_),
            .in3(N__9536),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22851),
            .ce(),
            .sr(N__22495));
    defparam \uu2.l_count_6_LC_1_5_0 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_1_5_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_1_5_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_6_LC_1_5_0  (
            .in0(N__8343),
            .in1(N__8276),
            .in2(_gnd_net_),
            .in3(N__8264),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22843),
            .ce(),
            .sr(N__22512));
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_5_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_1_5_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_1_5_1  (
            .in0(N__8262),
            .in1(N__8519),
            .in2(N__8295),
            .in3(N__8364),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_1_5_2 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_1_5_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_1_5_2 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu2.l_count_9_LC_1_5_2  (
            .in0(N__8456),
            .in1(N__8293),
            .in2(N__8247),
            .in3(N__8390),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22843),
            .ce(),
            .sr(N__22512));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_5_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_1_5_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_1_5_3  (
            .in0(N__8261),
            .in1(N__8518),
            .in2(N__8294),
            .in3(N__8363),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_7_LC_1_5_4 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_1_5_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_1_5_4 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.l_count_7_LC_1_5_4  (
            .in0(N__8344),
            .in1(N__8265),
            .in2(N__8478),
            .in3(N__8277),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22843),
            .ce(),
            .sr(N__22512));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_5_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_1_5_5  (
            .in0(_gnd_net_),
            .in1(N__8324),
            .in2(_gnd_net_),
            .in3(N__8365),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(\uu2.vbuf_count.un328_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_5_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_5_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_1_5_6  (
            .in0(N__8342),
            .in1(N__8474),
            .in2(N__8268),
            .in3(N__8263),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_1_5_7 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_1_5_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_1_5_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.l_count_8_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8238),
            .in3(N__8455),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22843),
            .ce(),
            .sr(N__22512));
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_6_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_1_6_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_1_6_0  (
            .in0(N__8415),
            .in1(N__8555),
            .in2(N__8427),
            .in3(N__8235),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_1_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_1_6_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_1_6_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__8489),
            .in2(_gnd_net_),
            .in3(N__8417),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22836),
            .ce(),
            .sr(N__22510));
    defparam \uu2.l_count_3_LC_1_6_2 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_1_6_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_1_6_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu2.l_count_3_LC_1_6_2  (
            .in0(N__8418),
            .in1(N__8389),
            .in2(N__8493),
            .in3(N__8439),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22836),
            .ce(),
            .sr(N__22510));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_1_6_3  (
            .in0(N__8438),
            .in1(N__8530),
            .in2(N__8561),
            .in3(N__8414),
            .lcout(\uu2.un306_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_1_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_1_6_4  (
            .in0(N__8473),
            .in1(N__8320),
            .in2(N__8457),
            .in3(N__8437),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_1_6_5 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_1_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_1_6_5  (
            .in0(N__8556),
            .in1(N__8416),
            .in2(N__8400),
            .in3(N__8397),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_1_6_6 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_1_6_6 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_1_6_6 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \uu2.l_count_4_LC_1_6_6  (
            .in0(N__8346),
            .in1(_gnd_net_),
            .in2(N__8370),
            .in3(N__8366),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22836),
            .ce(),
            .sr(N__22510));
    defparam \uu2.l_count_5_LC_1_6_7 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_1_6_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_1_6_7 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uu2.l_count_5_LC_1_6_7  (
            .in0(N__8367),
            .in1(_gnd_net_),
            .in2(N__8325),
            .in3(N__8345),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22836),
            .ce(),
            .sr(N__22510));
    defparam \uu0.sec_clk_LC_1_7_0 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_1_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__12238),
            .in2(_gnd_net_),
            .in3(N__16637),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \uu2.l_count_1_LC_1_7_1 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_1_7_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_1_7_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_1_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__8560),
            .in2(_gnd_net_),
            .in3(N__8532),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \buart.Z_rx.hh_0_LC_1_7_4 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_7_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_7_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_7_4  (
            .in0(N__8307),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_hh_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \buart.Z_rx.hh_1_LC_1_7_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_1_7_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_1_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19487),
            .lcout(buart__rx_hh_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \uu0.delay_line_1_LC_1_7_6 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_1_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_1_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_1_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16316),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \uu0.l_precount_0_LC_1_7_7 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_1_7_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_1_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_1_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8590),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22827),
            .ce(),
            .sr(N__22508));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(N__8997),
            .in2(_gnd_net_),
            .in3(N__9021),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__8689),
            .in2(_gnd_net_),
            .in3(N__8826),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_9_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(N__8562),
            .in2(_gnd_net_),
            .in3(N__8531),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI2Q224_6_LC_1_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI2Q224_6_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI2Q224_6_LC_1_9_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_user_nesr_RNI2Q224_6_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(N__22556),
            .in2(_gnd_net_),
            .in3(N__12378),
            .lcout(\uu2.un28_w_addr_user_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_9_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_9_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_1_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__12841),
            .in2(_gnd_net_),
            .in3(N__12880),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22816),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_9_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_9_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_1_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_1_9_6  (
            .in0(N__12842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22816),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_0_LC_1_10_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_10_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_10_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_10_0  (
            .in0(N__8631),
            .in1(N__8592),
            .in2(N__8652),
            .in3(N__8613),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22808),
            .ce(),
            .sr(N__22509));
    defparam \uu0.l_precount_3_LC_1_10_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_10_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_10_1  (
            .in0(N__8615),
            .in1(N__8650),
            .in2(N__8598),
            .in3(N__8634),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22808),
            .ce(),
            .sr(N__22509));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_2 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_10_2  (
            .in0(N__8630),
            .in1(N__8993),
            .in2(N__8651),
            .in3(N__8706),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_1_LC_1_10_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_10_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_precount_1_LC_1_10_3  (
            .in0(N__8593),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8632),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22808),
            .ce(),
            .sr(N__22509));
    defparam \uu0.l_precount_2_LC_1_10_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_10_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_10_4 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_1_10_4  (
            .in0(N__8633),
            .in1(N__8594),
            .in2(_gnd_net_),
            .in3(N__8614),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22808),
            .ce(),
            .sr(N__22509));
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_10_5 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI3Q7K1_2_LC_1_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI3Q7K1_2_LC_1_10_5  (
            .in0(N__8965),
            .in1(N__8892),
            .in2(N__8616),
            .in3(N__8729),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIO2782_16_LC_1_10_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNIO2782_16_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIO2782_16_LC_1_10_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu0.l_count_RNIO2782_16_LC_1_10_6  (
            .in0(N__10185),
            .in1(N__8591),
            .in2(N__8568),
            .in3(N__8928),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_6_LC_1_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_1_11_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_1_11_0 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \uu0.l_count_6_LC_1_11_0  (
            .in0(N__8691),
            .in1(N__8821),
            .in2(N__9049),
            .in3(N__16635),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22801),
            .ce(N__9226),
            .sr(N__22511));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_11_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_11_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_11_1  (
            .in0(N__8710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8731),
            .lcout(\uu0.un44_ci ),
            .ltout(\uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_11_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_11_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_11_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu0.l_count_2_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8565),
            .in3(N__8894),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22801),
            .ce(N__9226),
            .sr(N__22511));
    defparam \uu0.l_count_1_LC_1_11_3 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_11_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_1_11_3  (
            .in0(N__8711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8733),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22801),
            .ce(N__9226),
            .sr(N__22511));
    defparam \uu0.l_count_0_LC_1_11_4 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_11_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_11_4  (
            .in0(N__8732),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16633),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22801),
            .ce(N__9226),
            .sr(N__22511));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_5  (
            .in0(N__8893),
            .in1(N__8730),
            .in2(N__8712),
            .in3(N__8874),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_11_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_11_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_11_6  (
            .in0(N__8690),
            .in1(N__8820),
            .in2(N__8673),
            .in3(N__8847),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_12_LC_1_11_7 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_11_7 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_12_LC_1_11_7  (
            .in0(N__16634),
            .in1(N__10146),
            .in2(N__8670),
            .in3(N__10162),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22801),
            .ce(N__9226),
            .sr(N__22511));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_12_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_12_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_1_12_0  (
            .in0(N__9134),
            .in1(N__8845),
            .in2(N__8667),
            .in3(N__8872),
            .lcout(\uu0.un4_l_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_1  (
            .in0(N__9102),
            .in1(N__8966),
            .in2(_gnd_net_),
            .in3(N__9135),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_9_LC_1_12_2 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_1_12_2 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu0.l_count_9_LC_1_12_2  (
            .in0(N__9136),
            .in1(_gnd_net_),
            .in2(N__8970),
            .in3(N__9261),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22797),
            .ce(N__9227),
            .sr(N__22513));
    defparam \uu0.l_count_17_LC_1_12_3 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_1_12_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_1_12_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_17_LC_1_12_3  (
            .in0(N__8927),
            .in1(N__8666),
            .in2(N__9279),
            .in3(N__8750),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22797),
            .ce(N__9227),
            .sr(N__22513));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_12_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_12_4  (
            .in0(N__8665),
            .in1(N__9254),
            .in2(N__8751),
            .in3(N__8925),
            .lcout(\uu0.un220_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_1_12_5 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_1_12_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_1_12_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_16_LC_1_12_5  (
            .in0(N__8926),
            .in1(N__8749),
            .in2(N__9278),
            .in3(N__16621),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22797),
            .ce(N__9227),
            .sr(N__22513));
    defparam \uu0.l_count_3_LC_1_12_6 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_12_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_12_6 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu0.l_count_3_LC_1_12_6  (
            .in0(N__16623),
            .in1(N__8907),
            .in2(N__8901),
            .in3(N__8873),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22797),
            .ce(N__9227),
            .sr(N__22513));
    defparam \uu0.l_count_7_LC_1_12_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_1_12_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_7_LC_1_12_7  (
            .in0(N__8846),
            .in1(N__9042),
            .in2(N__8859),
            .in3(N__16622),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22797),
            .ce(N__9227),
            .sr(N__22513));
    defparam \uu0.l_count_18_LC_1_13_0 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_1_13_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu0.l_count_18_LC_1_13_0  (
            .in0(N__8832),
            .in1(N__8792),
            .in2(_gnd_net_),
            .in3(N__16618),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22793),
            .ce(N__9228),
            .sr(N__22515));
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_13_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIOIDD2_18_LC_1_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNIOIDD2_18_LC_1_13_1  (
            .in0(N__8825),
            .in1(N__8799),
            .in2(N__8793),
            .in3(N__9169),
            .lcout(),
            .ltout(\uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_13_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_15_LC_1_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_15_LC_1_13_2  (
            .in0(N__9060),
            .in1(N__8781),
            .in2(N__8772),
            .in3(N__8769),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_11_LC_1_13_3 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_1_13_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_1_13_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \uu0.l_count_11_LC_1_13_3  (
            .in0(N__9171),
            .in1(N__9287),
            .in2(N__8760),
            .in3(N__8757),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22793),
            .ce(N__9228),
            .sr(N__22515));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_14_0 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_14_0  (
            .in0(N__9077),
            .in1(N__9115),
            .in2(N__10144),
            .in3(N__10182),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_14_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_14_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_14_1  (
            .in0(N__9097),
            .in1(N__8957),
            .in2(N__9147),
            .in3(N__9170),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_14_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_14_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__9116),
            .in2(N__9153),
            .in3(N__10183),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_14_3 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_14_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_14_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_15_LC_1_14_3  (
            .in0(N__9076),
            .in1(N__9281),
            .in2(N__9150),
            .in3(N__16619),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22789),
            .ce(N__9229),
            .sr(N__22517));
    defparam \uu0.l_count_14_LC_1_14_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_14_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_14_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_1_14_4  (
            .in0(N__9280),
            .in1(N__9117),
            .in2(N__10145),
            .in3(N__10184),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22789),
            .ce(N__9229),
            .sr(N__22517));
    defparam \uu0.l_count_4_LC_1_14_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_14_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu0.l_count_4_LC_1_14_5  (
            .in0(N__9050),
            .in1(N__9016),
            .in2(_gnd_net_),
            .in3(N__16620),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22789),
            .ce(N__9229),
            .sr(N__22517));
    defparam \uu0.l_count_10_LC_1_14_6 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_14_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_14_6 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_10_LC_1_14_6  (
            .in0(N__9146),
            .in1(N__8964),
            .in2(N__9288),
            .in3(N__9098),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22789),
            .ce(N__9229),
            .sr(N__22517));
    defparam \uu0.l_count_RNIGTCU_15_LC_1_14_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIGTCU_15_LC_1_14_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uu0.l_count_RNIGTCU_15_LC_1_14_7  (
            .in0(N__9114),
            .in1(N__9096),
            .in2(N__9078),
            .in3(N__9015),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_5_LC_1_15_0 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_1_15_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_1_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu0.l_count_5_LC_1_15_0  (
            .in0(N__9054),
            .in1(N__8986),
            .in2(_gnd_net_),
            .in3(N__9020),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22785),
            .ce(N__9230),
            .sr(N__22518));
    defparam \uu0.l_count_8_LC_1_15_1 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_15_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_count_8_LC_1_15_1  (
            .in0(_gnd_net_),
            .in1(N__9286),
            .in2(_gnd_net_),
            .in3(N__8963),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22785),
            .ce(N__9230),
            .sr(N__22518));
    defparam \uu0.l_count_13_LC_1_16_5 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_16_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_16_5 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_13_LC_1_16_5  (
            .in0(N__9285),
            .in1(N__10116),
            .in2(N__10203),
            .in3(N__16636),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22782),
            .ce(N__9231),
            .sr(N__22521));
    defparam \uu2.r_addr_2_LC_2_4_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_2_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_2_4_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_2_4_0  (
            .in0(N__9398),
            .in1(N__9367),
            .in2(N__9434),
            .in3(N__9875),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22844),
            .ce(),
            .sr(N__22497));
    defparam \uu2.r_addr_1_LC_2_4_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_2_4_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.r_addr_1_LC_2_4_1  (
            .in0(N__9873),
            .in1(_gnd_net_),
            .in2(N__9371),
            .in3(N__9397),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22844),
            .ce(),
            .sr(N__22497));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_4_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_4_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__9872),
            .in2(_gnd_net_),
            .in3(N__22559),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_4_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_4_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__9195),
            .in2(_gnd_net_),
            .in3(N__9203),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(\uu2.trig_rd_is_det_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_0_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_2_4_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu2.r_addr_0_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9207),
            .in3(N__9363),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22844),
            .ce(),
            .sr(N__22497));
    defparam \uu2.trig_rd_det_1_LC_2_4_5 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_2_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9204),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22844),
            .ce(),
            .sr(N__22497));
    defparam \uu2.r_addr_4_LC_2_4_7 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_2_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_2_4_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_4_LC_2_4_7  (
            .in0(N__9874),
            .in1(N__9928),
            .in2(_gnd_net_),
            .in3(N__9899),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22844),
            .ce(),
            .sr(N__22497));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_5_0 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__9837),
            .in2(_gnd_net_),
            .in3(N__9926),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_2_5_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_2_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_2_5_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_2_5_1  (
            .in0(N__9182),
            .in1(N__9471),
            .in2(N__9189),
            .in3(N__9898),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22837),
            .ce(N__9315),
            .sr(N__22496));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_5_2  (
            .in0(N__9423),
            .in1(N__9395),
            .in2(N__9337),
            .in3(N__9361),
            .lcout(\uu2.un404_ci ),
            .ltout(\uu2.un404_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_7_LC_2_5_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_2_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_2_5_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_7_LC_2_5_3  (
            .in0(N__9485),
            .in1(N__9460),
            .in2(N__9498),
            .in3(N__9495),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22837),
            .ce(N__9315),
            .sr(N__22496));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_5_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__9484),
            .in2(_gnd_net_),
            .in3(N__9456),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_2_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_2_5_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_6_LC_2_5_5  (
            .in0(N__9927),
            .in1(N__9854),
            .in2(N__9464),
            .in3(N__9897),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22837),
            .ce(N__9315),
            .sr(N__22496));
    defparam \uu2.r_addr_esr_3_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_2_5_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_2_5_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_2_5_6  (
            .in0(N__9424),
            .in1(N__9396),
            .in2(N__9338),
            .in3(N__9362),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22837),
            .ce(N__9315),
            .sr(N__22496));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_2_6_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_2_6_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_2_6_4  (
            .in0(N__9771),
            .in1(N__11718),
            .in2(_gnd_net_),
            .in3(N__13389),
            .lcout(\uu2.mem0.N_76_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI84IJ2_2_LC_2_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI84IJ2_2_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI84IJ2_2_LC_2_6_6 .LUT_INIT=16'b1000000000010000;
    LogicCell40 \uu2.w_addr_displaying_RNI84IJ2_2_LC_2_6_6  (
            .in0(N__11895),
            .in1(N__13171),
            .in2(N__13521),
            .in3(N__13721),
            .lcout(\uu2.bitmap_pmux_sn_N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_2_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_2_7_6  (
            .in0(N__9585),
            .in1(N__11713),
            .in2(_gnd_net_),
            .in3(N__13827),
            .lcout(\uu2.mem0.N_73_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_2_7_7 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_2_7_7 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_2_7_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uu0.sec_clkD_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__12239),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.sec_clkDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22821),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_2_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_2_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_2_8_3  (
            .in0(N__9798),
            .in1(N__11712),
            .in2(_gnd_net_),
            .in3(N__11893),
            .lcout(\uu2.mem0.N_79_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_2_8_4 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_2_8_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_2_8_4  (
            .in0(N__12207),
            .in1(N__9537),
            .in2(N__11007),
            .in3(N__22560),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22817),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_5 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_2_8_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__9519),
            .in2(_gnd_net_),
            .in3(N__12234),
            .lcout(oneSecStrb),
            .ltout(oneSecStrb_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_2_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_2_8_6 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_2_8_6  (
            .in0(N__12503),
            .in1(N__10709),
            .in2(N__9513),
            .in3(N__15090),
            .lcout(\Lab_UT.dispString.un46_dOutP_i_m_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_7_LC_2_9_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_2_9_0 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_2_9_0  (
            .in0(N__12319),
            .in1(N__9507),
            .in2(N__9609),
            .in3(N__10583),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_7C_net ),
            .ce(N__9734),
            .sr(N__22472));
    defparam \uu2.w_addr_user_nesr_RNO_0_8_LC_2_9_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_8_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_8_LC_2_9_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_8_LC_2_9_1  (
            .in0(N__10582),
            .in1(N__9769),
            .in2(N__12356),
            .in3(N__12284),
            .lcout(),
            .ltout(\uu2.N_118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_2_9_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_2_9_2 .LUT_INIT=16'b0101000100000100;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_2_9_2  (
            .in0(N__12320),
            .in1(N__9608),
            .in2(N__9510),
            .in3(N__9584),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_7C_net ),
            .ce(N__9734),
            .sr(N__22472));
    defparam \uu2.w_addr_user_nesr_RNIHSS8_5_LC_2_9_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIHSS8_5_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIHSS8_5_LC_2_9_3 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIHSS8_5_LC_2_9_3  (
            .in0(N__12348),
            .in1(N__9768),
            .in2(_gnd_net_),
            .in3(N__12283),
            .lcout(\uu2.N_117 ),
            .ltout(\uu2.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_6_LC_2_9_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_6_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_6_LC_2_9_4 .LUT_INIT=16'b0001000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_6_LC_2_9_4  (
            .in0(N__12318),
            .in1(N__10553),
            .in2(N__9501),
            .in3(N__10585),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_7C_net ),
            .ce(N__9734),
            .sr(N__22472));
    defparam \uu2.w_addr_user_nesr_0_LC_2_9_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_0_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_0_LC_2_9_5 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \uu2.w_addr_user_nesr_0_LC_2_9_5  (
            .in0(N__10584),
            .in1(N__10552),
            .in2(N__11824),
            .in3(N__12317),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_7C_net ),
            .ce(N__9734),
            .sr(N__22472));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_2_9_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_2_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_2_9_6  (
            .in0(N__10586),
            .in1(N__11710),
            .in2(_gnd_net_),
            .in3(N__13260),
            .lcout(\uu2.mem0.N_75_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_2_9_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_2_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_2_9_7  (
            .in0(N__11711),
            .in1(N__9604),
            .in2(_gnd_net_),
            .in3(N__13350),
            .lcout(\uu2.mem0.N_74_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIG9RA_1_LC_2_10_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIG9RA_1_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIG9RA_1_LC_2_10_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu2.w_addr_user_RNIG9RA_1_LC_2_10_0  (
            .in0(N__11811),
            .in1(N__9558),
            .in2(N__11779),
            .in3(N__9564),
            .lcout(\uu2.N_225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIVCU1_8_LC_2_10_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIVCU1_8_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIVCU1_8_LC_2_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uu2.w_addr_user_nesr_RNIVCU1_8_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__9603),
            .in2(_gnd_net_),
            .in3(N__9580),
            .lcout(\uu2.N_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_2_10_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_2_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNINJD5_3_LC_2_10_2  (
            .in0(N__12281),
            .in1(N__9699),
            .in2(N__9770),
            .in3(N__9791),
            .lcout(\uu2.w_addr_user_3_i_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_2_10_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_2_10_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_3_LC_2_10_3  (
            .in0(N__9793),
            .in1(N__11775),
            .in2(N__9705),
            .in3(N__11813),
            .lcout(),
            .ltout(\uu2.N_150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_2_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_2_10_4 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_2_10_4  (
            .in0(N__12329),
            .in1(_gnd_net_),
            .in2(N__9552),
            .in3(N__12352),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__9741),
            .sr(N__22473));
    defparam \uu2.w_addr_user_nesr_2_LC_2_10_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_2_LC_2_10_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_2_LC_2_10_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu2.w_addr_user_nesr_2_LC_2_10_5  (
            .in0(N__9794),
            .in1(N__11814),
            .in2(N__11781),
            .in3(N__12328),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__9741),
            .sr(N__22473));
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_2_10_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_2_10_6 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIFBD5_3_LC_2_10_6  (
            .in0(N__11812),
            .in1(N__9700),
            .in2(N__11780),
            .in3(N__9792),
            .lcout(\uu2.N_115 ),
            .ltout(\uu2.N_115_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_5_LC_2_10_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_5_LC_2_10_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_5_LC_2_10_7 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \uu2.w_addr_user_nesr_5_LC_2_10_7  (
            .in0(N__12285),
            .in1(N__9764),
            .in2(N__9774),
            .in3(N__12330),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__9741),
            .sr(N__22473));
    defparam \buart.Z_tx.shifter_6_LC_2_11_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_11_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_11_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_11_0  (
            .in0(N__10983),
            .in1(N__9717),
            .in2(_gnd_net_),
            .in3(N__9984),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22798),
            .ce(N__10229),
            .sr(N__22514));
    defparam \buart.Z_tx.shifter_7_LC_2_11_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_2_11_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_2_11_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_7_LC_2_11_1  (
            .in0(N__9711),
            .in1(N__10984),
            .in2(_gnd_net_),
            .in3(N__9966),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22798),
            .ce(N__10229),
            .sr(N__22514));
    defparam \buart.Z_tx.shifter_8_LC_2_11_2 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_2_11_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_2_11_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \buart.Z_tx.shifter_8_LC_2_11_2  (
            .in0(N__10982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9948),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22798),
            .ce(N__10229),
            .sr(N__22514));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_11_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_2_11_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__10981),
            .in2(_gnd_net_),
            .in3(N__11066),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_2_11_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_2_11_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_2_11_5  (
            .in0(N__9704),
            .in1(N__11708),
            .in2(_gnd_net_),
            .in3(N__13728),
            .lcout(\uu2.mem0.N_78_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_2_11_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_2_11_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_2_11_6  (
            .in0(N__11709),
            .in1(N__12282),
            .in2(_gnd_net_),
            .in3(N__13506),
            .lcout(\uu2.mem0.N_77_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_0_LC_2_12_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_0_LC_2_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9651),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_12_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_12_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_1_LC_2_12_1  (
            .in0(N__10044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_12_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_12_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_2_LC_2_12_2  (
            .in0(N__10032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_12_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_12_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_3_LC_2_12_3  (
            .in0(N__10020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_12_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10008),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_12_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_2_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9996),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_12_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9978),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_12_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_12_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9960),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__9810),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_5_LC_2_13_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_2_13_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_2_13_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_2_13_0  (
            .in0(N__9941),
            .in1(N__9903),
            .in2(N__9844),
            .in3(N__9879),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22790),
            .ce(),
            .sr(N__22555));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_13_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_2_13_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_2_13_1  (
            .in0(N__12156),
            .in1(N__12177),
            .in2(_gnd_net_),
            .in3(N__22554),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_0_LC_2_13_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_2_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_2_13_2  (
            .in0(N__11010),
            .in1(N__10934),
            .in2(_gnd_net_),
            .in3(N__11067),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22790),
            .ce(),
            .sr(N__22555));
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_13_3 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_2_13_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__10202),
            .in2(_gnd_net_),
            .in3(N__10163),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_13_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_13_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_2_13_4  (
            .in0(N__10164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10140),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_14_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_14_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_14_0  (
            .in0(N__11011),
            .in1(N__10065),
            .in2(_gnd_net_),
            .in3(N__10107),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.shifter_0_LC_2_14_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_14_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__10098),
            .in2(_gnd_net_),
            .in3(N__11015),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.uart_tx_LC_2_14_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_14_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_14_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__11008),
            .in2(_gnd_net_),
            .in3(N__10092),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.shifter_2_LC_2_14_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_14_3  (
            .in0(N__11009),
            .in1(N__10050),
            .in2(_gnd_net_),
            .in3(N__10074),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.shifter_3_LC_2_14_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_14_4  (
            .in0(N__11012),
            .in1(N__10263),
            .in2(_gnd_net_),
            .in3(N__10059),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.shifter_4_LC_2_14_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_14_5  (
            .in0(N__10239),
            .in1(N__11014),
            .in2(_gnd_net_),
            .in3(N__10272),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \buart.Z_tx.shifter_5_LC_2_14_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_14_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_14_6  (
            .in0(N__11013),
            .in1(N__10257),
            .in2(_gnd_net_),
            .in3(N__10248),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22786),
            .ce(N__10233),
            .sr(N__22519));
    defparam \Lab_UT.didp.regrce1.q_RNI2NVO3_1_LC_4_1_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNI2NVO3_1_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNI2NVO3_1_LC_4_1_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNI2NVO3_1_LC_4_1_0  (
            .in0(N__14973),
            .in1(N__15465),
            .in2(N__15059),
            .in3(N__14034),
            .lcout(\Lab_UT.sec2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNI4PVO3_2_LC_4_1_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNI4PVO3_2_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNI4PVO3_2_LC_4_1_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNI4PVO3_2_LC_4_1_1  (
            .in0(N__14976),
            .in1(N__15390),
            .in2(N__13995),
            .in3(N__15055),
            .lcout(\Lab_UT.sec2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNI6RVO3_3_LC_4_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNI6RVO3_3_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNI6RVO3_3_LC_4_1_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNI6RVO3_3_LC_4_1_2  (
            .in0(N__14974),
            .in1(N__15431),
            .in2(N__15060),
            .in3(N__13946),
            .lcout(\Lab_UT.sec2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI85KT3_3_LC_4_1_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI85KT3_3_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI85KT3_3_LC_4_1_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI85KT3_3_LC_4_1_3  (
            .in0(N__14636),
            .in1(N__15051),
            .in2(N__17687),
            .in3(N__14975),
            .lcout(\Lab_UT.sec1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNIK3221_3_LC_4_1_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNIK3221_3_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNIK3221_3_LC_4_1_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNIK3221_3_LC_4_1_4  (
            .in0(N__15430),
            .in1(N__14635),
            .in2(N__17688),
            .in3(N__13945),
            .lcout(\Lab_UT.didp.did_alarmMatch_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_4_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_4_2_0 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \uu2.bitmap_93_LC_4_2_0  (
            .in0(N__13044),
            .in1(N__11242),
            .in2(N__11217),
            .in3(N__11288),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__22482));
    defparam \uu2.bitmap_221_LC_4_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_4_2_1 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_221_LC_4_2_1  (
            .in0(N__11241),
            .in1(N__11208),
            .in2(N__11292),
            .in3(N__13043),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__22482));
    defparam \uu2.bitmap_RNIAE522_93_LC_4_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIAE522_93_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIAE522_93_LC_4_2_2 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.bitmap_RNIAE522_93_LC_4_2_2  (
            .in0(N__13155),
            .in1(N__10218),
            .in2(N__10212),
            .in3(N__10881),
            .lcout(),
            .ltout(\uu2.bitmap_RNIAE522Z0Z_93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIMS86A_66_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIMS86A_66_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIMS86A_66_LC_4_2_3 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.bitmap_RNIMS86A_66_LC_4_2_3  (
            .in0(N__10335),
            .in1(N__13059),
            .in2(N__10299),
            .in3(N__10284),
            .lcout(\uu2.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_4_3_0 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_215_LC_4_3_0  (
            .in0(N__11147),
            .in1(N__10389),
            .in2(N__11118),
            .in3(N__12986),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__22479));
    defparam \uu2.bitmap_RNIKL222_212_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKL222_212_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKL222_212_LC_4_3_1 .LUT_INIT=16'b0010001011111100;
    LogicCell40 \uu2.bitmap_RNIKL222_212_LC_4_3_1  (
            .in0(N__10278),
            .in1(N__13323),
            .in2(N__10296),
            .in3(N__10350),
            .lcout(),
            .ltout(\uu2.bitmap_RNIKL222Z0Z_212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI9ITA5_3_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI9ITA5_3_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI9ITA5_3_LC_4_3_2 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI9ITA5_3_LC_4_3_2  (
            .in0(N__10334),
            .in1(N__11463),
            .in2(N__10287),
            .in3(N__13720),
            .lcout(\uu2.bitmap_pmux_27_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_4_4_0 .LUT_INIT=16'b0001001100100101;
    LogicCell40 \uu2.bitmap_308_LC_4_4_0  (
            .in0(N__13002),
            .in1(N__10396),
            .in2(N__11133),
            .in3(N__11166),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_212_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_4_4_1 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \uu2.bitmap_212_LC_4_4_1  (
            .in0(N__11165),
            .in1(N__11120),
            .in2(N__10401),
            .in3(N__13001),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_84_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_4_4_2 .LUT_INIT=16'b0001000000111101;
    LogicCell40 \uu2.bitmap_84_LC_4_4_2  (
            .in0(N__13004),
            .in1(N__10398),
            .in2(N__11135),
            .in3(N__11168),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_180_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_4_4_3 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_180_LC_4_4_3  (
            .in0(N__11164),
            .in1(N__11119),
            .in2(N__10400),
            .in3(N__13000),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_52_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_4_4_4 .LUT_INIT=16'b1111011101101101;
    LogicCell40 \uu2.bitmap_52_LC_4_4_4  (
            .in0(N__13003),
            .in1(N__10397),
            .in2(N__11134),
            .in3(N__11167),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_RNIU2IS_52_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIU2IS_52_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIU2IS_52_LC_4_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIU2IS_52_LC_4_4_5  (
            .in0(N__13804),
            .in1(N__10413),
            .in2(_gnd_net_),
            .in3(N__10407),
            .lcout(\uu2.N_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_4_4_6 .LUT_INIT=16'b0010011110011111;
    LogicCell40 \uu2.bitmap_87_LC_4_4_6  (
            .in0(N__13005),
            .in1(N__10399),
            .in2(N__11136),
            .in3(N__11169),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__22477));
    defparam \uu2.bitmap_RNIC6I01_84_LC_4_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIC6I01_84_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIC6I01_84_LC_4_4_7 .LUT_INIT=16'b0100001101001111;
    LogicCell40 \uu2.bitmap_RNIC6I01_84_LC_4_4_7  (
            .in0(N__10362),
            .in1(N__13321),
            .in2(N__13151),
            .in3(N__10356),
            .lcout(\uu2.bitmap_pmux_24_i_m2_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAJJL8_8_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAJJL8_8_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAJJL8_8_LC_4_5_0 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \uu2.w_addr_displaying_RNIAJJL8_8_LC_4_5_0  (
            .in0(N__11576),
            .in1(N__10493),
            .in2(N__11733),
            .in3(N__13441),
            .lcout(\uu2.un51_w_data_displaying ),
            .ltout(\uu2.un51_w_data_displaying_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_5_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_5_1  (
            .in0(N__10803),
            .in1(_gnd_net_),
            .in2(N__10344),
            .in3(N__11699),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_5_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__11992),
            .in2(_gnd_net_),
            .in3(N__13115),
            .lcout(\uu2.w_addr_displaying_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_5_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_5_3 .LUT_INIT=16'b1111101000111010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_5_3  (
            .in0(N__10659),
            .in1(N__10317),
            .in2(N__11717),
            .in3(N__10421),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_1_LC_4_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_1_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_0_1_LC_4_5_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI25P31_0_1_LC_4_5_4  (
            .in0(N__13818),
            .in1(N__11997),
            .in2(_gnd_net_),
            .in3(N__13117),
            .lcout(\uu2.un49_w_data_displaying_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_5_5 .LUT_INIT=16'b1110111000101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_5_5  (
            .in0(N__12132),
            .in1(N__11700),
            .in2(N__10845),
            .in3(N__10422),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_1_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_1_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI25P31_1_LC_4_5_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI25P31_1_LC_4_5_6  (
            .in0(N__13817),
            .in1(N__11996),
            .in2(_gnd_net_),
            .in3(N__13116),
            .lcout(\uu2.un31_w_data_displaying_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIASLS1_1_LC_4_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIASLS1_1_LC_4_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIASLS1_1_LC_4_5_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIASLS1_1_LC_4_5_7  (
            .in0(N__13118),
            .in1(N__11575),
            .in2(N__12012),
            .in3(N__13816),
            .lcout(\uu2.un31_w_data_displaying_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_4_6_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8NSO_4_LC_4_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_RNI8NSO_4_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__13494),
            .in2(_gnd_net_),
            .in3(N__11988),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIOELE1_4_LC_4_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIOELE1_4_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIOELE1_4_LC_4_6_1 .LUT_INIT=16'b0011100100110110;
    LogicCell40 \uu2.w_addr_displaying_RNIOELE1_4_LC_4_6_1  (
            .in0(N__13160),
            .in1(N__11888),
            .in2(N__13502),
            .in3(N__13707),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI6RE03_3_LC_4_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI6RE03_3_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI6RE03_3_LC_4_6_2 .LUT_INIT=16'b0000100100100100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI6RE03_3_LC_4_6_2  (
            .in0(N__13709),
            .in1(N__11599),
            .in2(N__10440),
            .in3(N__13161),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_i5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI1U7M3_7_LC_4_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI1U7M3_7_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI1U7M3_7_LC_4_6_3 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \uu2.w_addr_displaying_RNI1U7M3_7_LC_4_6_3  (
            .in0(N__13342),
            .in1(_gnd_net_),
            .in2(N__10437),
            .in3(N__13819),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_29_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI30QB21_7_LC_4_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI30QB21_7_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI30QB21_7_LC_4_6_4 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \uu2.w_addr_displaying_RNI30QB21_7_LC_4_6_4  (
            .in0(N__11586),
            .in1(N__10434),
            .in2(N__10425),
            .in3(N__10512),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNICAPH1_2_LC_4_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNICAPH1_2_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNICAPH1_2_LC_4_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNICAPH1_2_LC_4_6_5  (
            .in0(N__13159),
            .in1(N__11889),
            .in2(N__12011),
            .in3(N__13708),
            .lcout(\uu2.un15_w_data_displaying_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_4_7_0 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_4_7_0 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_40_LC_4_7_0  (
            .in0(N__11445),
            .in1(N__11412),
            .in2(N__11370),
            .in3(N__11325),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_40C_net ),
            .ce(),
            .sr(N__22475));
    defparam \uu2.bitmap_RNI1PH82_40_LC_4_7_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI1PH82_40_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI1PH82_40_LC_4_7_1 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \uu2.bitmap_RNI1PH82_40_LC_4_7_1  (
            .in0(N__10524),
            .in1(N__13740),
            .in2(N__11496),
            .in3(N__13710),
            .lcout(),
            .ltout(\uu2.bitmap_RNI1PH82Z0Z_40_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI208E6_40_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI208E6_40_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI208E6_40_LC_4_7_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uu2.bitmap_RNI208E6_40_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__12033),
            .in2(N__10518),
            .in3(N__12024),
            .lcout(),
            .ltout(\uu2.N_401_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIKE7JD_4_LC_4_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIKE7JD_4_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIKE7JD_4_LC_4_7_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_RNIKE7JD_4_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__11622),
            .in2(N__10515),
            .in3(N__12039),
            .lcout(\uu2.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_4_8_0 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_4_8_0  (
            .in0(N__15988),
            .in1(N__12520),
            .in2(N__10710),
            .in3(N__12141),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22803),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_4_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_4_8_1 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \Lab_UT.dispString.rdy_LC_4_8_1  (
            .in0(N__12519),
            .in1(N__10704),
            .in2(_gnd_net_),
            .in3(N__15989),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22803),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNII08G4_1_LC_4_8_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNII08G4_1_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNII08G4_1_LC_4_8_2 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNII08G4_1_LC_4_8_2  (
            .in0(N__10506),
            .in1(N__13442),
            .in2(N__10497),
            .in3(N__11580),
            .lcout(\uu2.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_8_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_4_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_4_8_3  (
            .in0(N__11707),
            .in1(N__11825),
            .in2(_gnd_net_),
            .in3(N__13172),
            .lcout(\uu2.mem0.N_81_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_8_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_4_8_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_4_8_4  (
            .in0(N__11754),
            .in1(N__11706),
            .in2(_gnd_net_),
            .in3(N__12018),
            .lcout(\uu2.mem0.N_80_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_4_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_4_8_5 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_4_8_5  (
            .in0(N__12518),
            .in1(N__10708),
            .in2(N__16007),
            .in3(N__12102),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22803),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_9_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_9_0 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_4_9_0  (
            .in0(N__10737),
            .in1(N__12620),
            .in2(N__10596),
            .in3(N__10767),
            .lcout(\uu2.mem0.N_72_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_data_0_o2_0_4_LC_4_9_1 .C_ON=1'b0;
    defparam \uu2.w_data_0_o2_0_4_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_data_0_o2_0_4_LC_4_9_1 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \uu2.w_data_0_o2_0_4_LC_4_9_1  (
            .in0(N__12618),
            .in1(N__12119),
            .in2(_gnd_net_),
            .in3(N__12726),
            .lcout(\uu2.N_111 ),
            .ltout(\uu2.N_111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_4_9_2 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_4_9_2 .LUT_INIT=16'b1011101110110011;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_4_9_2  (
            .in0(N__10736),
            .in1(N__22860),
            .in2(N__10638),
            .in3(N__10766),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_9_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_4_9_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_4_9_3  (
            .in0(N__10765),
            .in1(N__12621),
            .in2(_gnd_net_),
            .in3(N__12124),
            .lcout(),
            .ltout(\uu2.mem0.w_data_i_a2_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_4 .LUT_INIT=16'b0000100010111011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_9_4  (
            .in0(N__12729),
            .in1(N__10738),
            .in2(N__10611),
            .in3(N__10837),
            .lcout(\uu2.mem0.N_82_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_4_9_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_4_9_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_4_9_5  (
            .in0(_gnd_net_),
            .in1(N__12123),
            .in2(_gnd_net_),
            .in3(N__12728),
            .lcout(\uu2.mem0.N_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_a2_LC_4_9_6 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a2_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a2_LC_4_9_6 .LUT_INIT=16'b0000000000011000;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a2_LC_4_9_6  (
            .in0(N__12727),
            .in1(N__12619),
            .in2(N__12128),
            .in3(N__10764),
            .lcout(\uu2.N_144 ),
            .ltout(\uu2.N_144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIU0804_6_LC_4_9_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIU0804_6_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIU0804_6_LC_4_9_7 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \uu2.w_addr_user_nesr_RNIU0804_6_LC_4_9_7  (
            .in0(N__10587),
            .in1(N__10554),
            .in2(N__10527),
            .in3(N__10735),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_4_10_0 .LUT_INIT=16'b1011000110111011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_4_10_0  (
            .in0(N__12596),
            .in1(N__10875),
            .in2(N__12517),
            .in3(N__13913),
            .lcout(\Lab_UT.dispString.dOut_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_10_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_17_LC_4_10_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_17_LC_4_10_1  (
            .in0(N__10752),
            .in1(N__10802),
            .in2(N__11543),
            .in3(N__10652),
            .lcout(),
            .ltout(\uu2.mem0.w_data_0_a2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_10_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_10_2 .LUT_INIT=16'b1011101000110011;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_10_2  (
            .in0(N__10779),
            .in1(N__10844),
            .in2(N__10818),
            .in3(N__10740),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_4_10_3 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_o2_0_LC_4_10_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \uu2.un28_w_addr_user_i_0_o2_0_LC_4_10_3  (
            .in0(N__10801),
            .in1(N__10778),
            .in2(N__11542),
            .in3(N__10651),
            .lcout(\uu2.N_109 ),
            .ltout(\uu2.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_i_0_tz_0_LC_4_10_4 .C_ON=1'b0;
    defparam \uu2.w_addr_i_0_tz_0_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_i_0_tz_0_LC_4_10_4 .LUT_INIT=16'b0000001111111111;
    LogicCell40 \uu2.w_addr_i_0_tz_0_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__10751),
            .in2(N__10743),
            .in3(N__10739),
            .lcout(\uu2.w_addr_i_0_tzZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIOG7L_1_LC_4_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_1_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_1_LC_4_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIOG7L_1_LC_4_11_0  (
            .in0(N__12569),
            .in1(N__12667),
            .in2(N__12521),
            .in3(N__12712),
            .lcout(\Lab_UT.dispString.dOutP_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_4_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_4_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_4_11_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_4_11_1  (
            .in0(N__12713),
            .in1(N__12697),
            .in2(N__12507),
            .in3(N__12571),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22791),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_4_11_3 .LUT_INIT=16'b0000011111110111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_4_11_3  (
            .in0(N__15994),
            .in1(N__14805),
            .in2(N__12505),
            .in3(N__14033),
            .lcout(\Lab_UT.dispString.N_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_11_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dispString.cnt_RNIFV4E_1_LC_4_11_4  (
            .in0(N__12568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12666),
            .lcout(\Lab_UT.dispString.N_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_4_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_4_11_5 .LUT_INIT=16'b1010111111101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_4_11_5  (
            .in0(N__12668),
            .in1(N__13947),
            .in2(N__12506),
            .in3(N__12570),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_4_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_4_11_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_4_11_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_4_11_6  (
            .in0(N__10866),
            .in1(N__10680),
            .in2(N__10668),
            .in3(N__10665),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22791),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_4_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_4_11_7 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_4_11_7  (
            .in0(N__15993),
            .in1(N__14841),
            .in2(N__12504),
            .in3(N__13589),
            .lcout(\Lab_UT.dispString.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_2_LC_4_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_4_12_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_4_12_0 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_4_12_0  (
            .in0(N__12574),
            .in1(_gnd_net_),
            .in2(N__12492),
            .in3(N__12687),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22787),
            .ce(),
            .sr(N__22499));
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_4_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_4_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_3_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__12441),
            .in2(_gnd_net_),
            .in3(N__12572),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_12_2 .LUT_INIT=16'b1101111110001111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_4_12_2  (
            .in0(N__12681),
            .in1(N__14643),
            .in2(N__10869),
            .in3(N__14507),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_0_LC_4_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_4_12_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_4_12_3 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_4_12_3  (
            .in0(N__12685),
            .in1(N__12442),
            .in2(N__16013),
            .in3(N__12575),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22787),
            .ce(),
            .sr(N__22499));
    defparam \Lab_UT.dispString.cnt_1_LC_4_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_4_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_4_12_4  (
            .in0(N__12573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12686),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22787),
            .ce(),
            .sr(N__22499));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_13_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_4_13_0 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_4_13_0  (
            .in0(N__10910),
            .in1(N__11081),
            .in2(N__10941),
            .in3(N__11056),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_3_LC_4_13_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_4_13_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_4_13_1 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_4_13_1  (
            .in0(N__11027),
            .in1(N__11065),
            .in2(N__10860),
            .in3(N__10857),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22783),
            .ce(),
            .sr(N__22522));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_13_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_13_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_4_13_2  (
            .in0(_gnd_net_),
            .in1(N__10856),
            .in2(_gnd_net_),
            .in3(N__10935),
            .lcout(),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_13_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_13_3 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_4_13_3  (
            .in0(N__11080),
            .in1(N__10908),
            .in2(N__11091),
            .in3(N__12798),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_13_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_4_13_4 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_4_13_4  (
            .in0(N__10909),
            .in1(_gnd_net_),
            .in2(N__11088),
            .in3(N__10936),
            .lcout(),
            .ltout(\buart.Z_tx.un1_bitcount_c2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_2_LC_4_13_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_4_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_4_13_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_4_13_5  (
            .in0(N__11026),
            .in1(N__11064),
            .in2(N__11085),
            .in3(N__11082),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22783),
            .ce(),
            .sr(N__22522));
    defparam \buart.Z_tx.bitcount_1_LC_4_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_4_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_4_13_7 .LUT_INIT=16'b1111110011110110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_4_13_7  (
            .in0(N__11057),
            .in1(N__10911),
            .in2(N__11031),
            .in3(N__10940),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22783),
            .ce(),
            .sr(N__22522));
    defparam \uu2.bitmap_314_LC_5_1_0 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_5_1_0 .LUT_INIT=16'b0000011000011011;
    LogicCell40 \uu2.bitmap_314_LC_5_1_0  (
            .in0(N__11214),
            .in1(N__11247),
            .in2(N__11290),
            .in3(N__13035),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__22485));
    defparam \uu2.bitmap_218_LC_5_1_1 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_5_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_5_1_1 .LUT_INIT=16'b0001000100000101;
    LogicCell40 \uu2.bitmap_218_LC_5_1_1  (
            .in0(N__13034),
            .in1(N__11277),
            .in2(N__11252),
            .in3(N__11213),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__22485));
    defparam \uu2.bitmap_90_LC_5_1_2 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_5_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_5_1_2 .LUT_INIT=16'b0001010000011101;
    LogicCell40 \uu2.bitmap_90_LC_5_1_2  (
            .in0(N__11216),
            .in1(N__11251),
            .in2(N__11291),
            .in3(N__13037),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__22485));
    defparam \uu2.bitmap_RNILGG61_90_LC_5_1_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNILGG61_90_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNILGG61_90_LC_5_1_3 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNILGG61_90_LC_5_1_3  (
            .in0(N__10896),
            .in1(N__13170),
            .in2(N__10890),
            .in3(N__13337),
            .lcout(\uu2.bitmap_pmux_25_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_5_1_4 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_5_1_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_186_LC_5_1_4  (
            .in0(N__11212),
            .in1(N__11243),
            .in2(N__11289),
            .in3(N__13033),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__22485));
    defparam \uu2.bitmap_58_LC_5_1_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_5_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_5_1_5 .LUT_INIT=16'b1111011101101101;
    LogicCell40 \uu2.bitmap_58_LC_5_1_5  (
            .in0(N__13036),
            .in1(N__11281),
            .in2(N__11253),
            .in3(N__11215),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__22485));
    defparam \uu2.bitmap_RNI7GKQ_58_LC_5_1_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI7GKQ_58_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI7GKQ_58_LC_5_1_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNI7GKQ_58_LC_5_1_6  (
            .in0(N__13336),
            .in1(N__11184),
            .in2(_gnd_net_),
            .in3(N__11178),
            .lcout(),
            .ltout(\uu2.N_216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIS4UH1_314_LC_5_1_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIS4UH1_314_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIS4UH1_314_LC_5_1_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.bitmap_RNIS4UH1_314_LC_5_1_7  (
            .in0(_gnd_net_),
            .in1(N__12095),
            .in2(N__11172),
            .in3(N__13823),
            .lcout(\uu2.bitmap_RNIS4UH1Z0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI41KT3_1_LC_5_2_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI41KT3_1_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI41KT3_1_LC_5_2_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI41KT3_1_LC_5_2_0  (
            .in0(N__14948),
            .in1(N__17928),
            .in2(N__15572),
            .in3(N__15024),
            .lcout(\Lab_UT.sec1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI63KT3_2_LC_5_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI63KT3_2_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI63KT3_2_LC_5_2_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI63KT3_2_LC_5_2_1  (
            .in0(N__15026),
            .in1(N__17515),
            .in2(N__15524),
            .in3(N__14950),
            .lcout(\Lab_UT.sec1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNI49824_0_LC_5_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNI49824_0_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNI49824_0_LC_5_2_2 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNI49824_0_LC_5_2_2  (
            .in0(N__13912),
            .in1(N__15025),
            .in2(N__14962),
            .in3(N__15860),
            .lcout(\Lab_UT.min2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNI6B824_1_LC_5_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNI6B824_1_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNI6B824_1_LC_5_2_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNI6B824_1_LC_5_2_3  (
            .in0(N__15021),
            .in1(N__15903),
            .in2(N__14603),
            .in3(N__14949),
            .lcout(\Lab_UT.min2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNI8D824_2_LC_5_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNI8D824_2_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNI8D824_2_LC_5_2_4 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNI8D824_2_LC_5_2_4  (
            .in0(N__14951),
            .in1(N__15824),
            .in2(N__14388),
            .in3(N__15023),
            .lcout(\Lab_UT.min2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNIAF824_3_LC_5_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNIAF824_3_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNIAF824_3_LC_5_2_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNIAF824_3_LC_5_2_5  (
            .in0(N__15022),
            .in1(N__15726),
            .in2(N__14508),
            .in3(N__14952),
            .lcout(\Lab_UT.min2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_5_3_0 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_296_LC_5_3_0  (
            .in0(N__11316),
            .in1(N__11353),
            .in2(N__11407),
            .in3(N__11436),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_200_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_5_3_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_200_LC_5_3_1  (
            .in0(N__11434),
            .in1(N__11392),
            .in2(N__11362),
            .in3(N__11314),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_72_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_5_3_2 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_72_LC_5_3_2  (
            .in0(N__11317),
            .in1(N__11354),
            .in2(N__11408),
            .in3(N__11437),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_RNIC4D61_72_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIC4D61_72_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIC4D61_72_LC_5_3_3 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \uu2.bitmap_RNIC4D61_72_LC_5_3_3  (
            .in0(N__11481),
            .in1(N__13119),
            .in2(N__11475),
            .in3(N__13322),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_24_i_m2_bm_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI1UT12_75_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI1UT12_75_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI1UT12_75_LC_5_3_4 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \uu2.bitmap_RNI1UT12_75_LC_5_3_4  (
            .in0(N__13120),
            .in1(N__11451),
            .in2(N__11466),
            .in3(N__11457),
            .lcout(\uu2.bitmap_RNI1UT12Z0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_5_3_5 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.bitmap_75_LC_5_3_5  (
            .in0(N__11438),
            .in1(N__11402),
            .in2(N__11363),
            .in3(N__11318),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_203_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_5_3_6 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \uu2.bitmap_203_LC_5_3_6  (
            .in0(N__11315),
            .in1(N__11352),
            .in2(N__11406),
            .in3(N__11435),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_168_LC_5_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_5_3_7 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_168_LC_5_3_7  (
            .in0(N__11433),
            .in1(N__11391),
            .in2(N__11361),
            .in3(N__11313),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__22483));
    defparam \uu2.bitmap_69_LC_5_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_5_4_0 .LUT_INIT=16'b0010011110011111;
    LogicCell40 \uu2.bitmap_69_LC_5_4_0  (
            .in0(N__14567),
            .in1(N__14538),
            .in2(N__13870),
            .in3(N__14875),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.bitmap_197_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_5_4_1 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_197_LC_5_4_1  (
            .in0(N__14537),
            .in1(N__13857),
            .in2(N__14887),
            .in3(N__14568),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.bitmap_RNI10J51_69_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI10J51_69_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI10J51_69_LC_5_4_2 .LUT_INIT=16'b0100010000111111;
    LogicCell40 \uu2.bitmap_RNI10J51_69_LC_5_4_2  (
            .in0(N__11562),
            .in1(N__13113),
            .in2(N__11556),
            .in3(N__13319),
            .lcout(\uu2.bitmap_pmux_25_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un437_ci_0_LC_5_4_3 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un437_ci_0_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un437_ci_0_LC_5_4_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu2.vbuf_w_addr_displaying.counter_gen_label_7__un437_ci_0_LC_5_4_3  (
            .in0(N__13250),
            .in1(N__13477),
            .in2(_gnd_net_),
            .in3(N__13384),
            .lcout(),
            .ltout(\uu2.un437_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_7_LC_5_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_5_4_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_7_LC_5_4_4  (
            .in0(N__12962),
            .in1(N__11920),
            .in2(N__11547),
            .in3(N__13320),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_5_4_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_displaying_4_LC_5_4_5  (
            .in0(N__11924),
            .in1(N__12960),
            .in2(_gnd_net_),
            .in3(N__13478),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.w_addr_displaying_5_LC_5_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_5_4_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_displaying_5_LC_5_4_6  (
            .in0(N__12961),
            .in1(N__13385),
            .in2(N__13493),
            .in3(N__11925),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.w_addr_displaying_0_LC_5_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_5_4_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_0_LC_5_4_7  (
            .in0(N__13114),
            .in1(_gnd_net_),
            .in2(N__11930),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_69C_net ),
            .ce(),
            .sr(N__22480));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_5_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_5_5_0 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_5_5_0  (
            .in0(N__11705),
            .in1(N__11544),
            .in2(_gnd_net_),
            .in3(N__11732),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_8_LC_5_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_5_5_1 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_8_LC_5_5_1  (
            .in0(N__13812),
            .in1(N__13420),
            .in2(N__11931),
            .in3(N__12941),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_8C_net ),
            .ce(),
            .sr(N__22478));
    defparam \uu2.w_addr_displaying_RNIQN495_8_LC_5_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIQN495_8_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIQN495_8_LC_5_5_2 .LUT_INIT=16'b0001111100111111;
    LogicCell40 \uu2.w_addr_displaying_RNIQN495_8_LC_5_5_2  (
            .in0(N__12939),
            .in1(N__11502),
            .in2(N__13431),
            .in3(N__13810),
            .lcout(\uu2.un33_w_data_displaying ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_5_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_5_5_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \uu2.w_addr_displaying_RNI0ES07_8_LC_5_5_3  (
            .in0(N__13811),
            .in1(N__12940),
            .in2(N__13443),
            .in3(N__11704),
            .lcout(\uu2.un21_w_addr_displaying_i ),
            .ltout(\uu2.un21_w_addr_displaying_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_5_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_5_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_5_5_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_displaying_RNI47N27_8_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11625),
            .in3(N__22557),
            .lcout(\uu2.un21_w_addr_displaying_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIS6T61_1_LC_5_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIS6T61_1_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIS6T61_1_LC_5_5_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIS6T61_1_LC_5_5_6  (
            .in0(N__11987),
            .in1(N__13702),
            .in2(_gnd_net_),
            .in3(N__13809),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_5_6_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_5_6_1  (
            .in0(N__13168),
            .in1(N__11887),
            .in2(N__12013),
            .in3(N__13706),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__13548),
            .sr(N__22476));
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_6_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_6_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_1_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__12000),
            .in2(_gnd_net_),
            .in3(N__13169),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__13548),
            .sr(N__22476));
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_5_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_5_6_4 .LUT_INIT=16'b0101100011000000;
    LogicCell40 \uu2.w_addr_displaying_RNIGEPH1_4_LC_5_6_4  (
            .in0(N__13704),
            .in1(N__13498),
            .in2(N__11894),
            .in3(N__11998),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIUNPV1_2_LC_5_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIUNPV1_2_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIUNPV1_2_LC_5_6_5 .LUT_INIT=16'b0110001101101100;
    LogicCell40 \uu2.w_addr_displaying_RNIUNPV1_2_LC_5_6_5  (
            .in0(N__11999),
            .in1(N__11886),
            .in2(N__11604),
            .in3(N__13705),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m15_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIOM1S6_2_LC_5_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIOM1S6_2_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIOM1S6_2_LC_5_6_6 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \uu2.w_addr_displaying_RNIOM1S6_2_LC_5_6_6  (
            .in0(N__13212),
            .in1(N__11616),
            .in2(N__11607),
            .in3(N__11603),
            .lcout(\uu2.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_5_6_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8NSO_2_LC_5_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI8NSO_2_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__11882),
            .in2(_gnd_net_),
            .in3(N__13703),
            .lcout(\uu2.un15_w_data_displaying_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIVKR41_180_LC_5_7_0 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIVKR41_180_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIVKR41_180_LC_5_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIVKR41_180_LC_5_7_0  (
            .in0(N__13696),
            .in1(N__12096),
            .in2(_gnd_net_),
            .in3(N__12081),
            .lcout(),
            .ltout(\uu2.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIAKAQ2_7_LC_5_7_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIAKAQ2_7_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIAKAQ2_7_LC_5_7_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.w_addr_displaying_RNIAKAQ2_7_LC_5_7_1  (
            .in0(N__13701),
            .in1(N__13338),
            .in2(N__12072),
            .in3(N__12069),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_RNIAKAQ2Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI206J5_7_LC_5_7_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI206J5_7_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI206J5_7_LC_5_7_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_RNI206J5_7_LC_5_7_2  (
            .in0(_gnd_net_),
            .in1(N__12060),
            .in2(N__12051),
            .in3(N__12048),
            .lcout(\uu2.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIJHPH1_2_LC_5_7_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIJHPH1_2_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIJHPH1_2_LC_5_7_3 .LUT_INIT=16'b0000010100001110;
    LogicCell40 \uu2.w_addr_displaying_RNIJHPH1_2_LC_5_7_3  (
            .in0(N__11860),
            .in1(N__13698),
            .in2(N__13346),
            .in3(N__11986),
            .lcout(\uu2.bitmap_pmux_sn_N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_5_7_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIM0T61_2_LC_5_7_4 .LUT_INIT=16'b1111000000000101;
    LogicCell40 \uu2.w_addr_displaying_RNIM0T61_2_LC_5_7_4  (
            .in0(N__13697),
            .in1(_gnd_net_),
            .in2(N__12010),
            .in3(N__11859),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIELSJ2_111_LC_5_7_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIELSJ2_111_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIELSJ2_111_LC_5_7_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \uu2.bitmap_RNIELSJ2_111_LC_5_7_5  (
            .in0(N__13614),
            .in1(_gnd_net_),
            .in2(N__12027),
            .in3(N__12213),
            .lcout(\uu2.bitmap_RNIELSJ2Z0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_2_LC_5_8_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_5_8_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_2_LC_5_8_0  (
            .in0(N__11881),
            .in1(N__12017),
            .in2(N__13176),
            .in3(N__11929),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \uu2.w_addr_user_1_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_5_8_1 .LUT_INIT=16'b0001001011110000;
    LogicCell40 \uu2.w_addr_user_1_LC_5_8_1  (
            .in0(N__11826),
            .in1(N__12315),
            .in2(N__11768),
            .in3(N__12376),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \uu2.w_addr_user_4_LC_5_8_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_5_8_2 .LUT_INIT=16'b0101000011010010;
    LogicCell40 \uu2.w_addr_user_4_LC_5_8_2  (
            .in0(N__12377),
            .in1(N__12360),
            .in2(N__12280),
            .in3(N__12316),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \uu2.bitmap_111_LC_5_8_3 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_5_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_5_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12243),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \uu2.vram_rd_clk_det_0_LC_5_8_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_5_8_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_5_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_5_8_4  (
            .in0(N__12206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \uu2.vram_rd_clk_det_1_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_5_8_5 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_5_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_5_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12170),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_2C_net ),
            .ce(),
            .sr(N__22474));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_0 .LUT_INIT=16'b0111011101010111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_5_9_0  (
            .in0(N__12511),
            .in1(N__12600),
            .in2(N__12698),
            .in3(N__14047),
            .lcout(\Lab_UT.dispString.dOutP_1_iv_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_2 .LUT_INIT=16'b0100111101000101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_2  (
            .in0(N__12603),
            .in1(N__12714),
            .in2(N__12525),
            .in3(N__15573),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOut_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(N__12694),
            .in2(N__12135),
            .in3(N__12384),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22795),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_5_9_4 .LUT_INIT=16'b0101111101111111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_5_LC_5_9_4  (
            .in0(N__12512),
            .in1(N__12601),
            .in2(N__12699),
            .in3(N__14048),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_9_6 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_5_9_6  (
            .in0(N__16008),
            .in1(N__14732),
            .in2(N__12524),
            .in3(N__13991),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_41_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_9_7 .LUT_INIT=16'b1101110100001111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_5_9_7  (
            .in0(N__14379),
            .in1(N__12513),
            .in2(N__12741),
            .in3(N__12602),
            .lcout(\Lab_UT.dispString.dOut_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_5_10_1 .LUT_INIT=16'b0001010100011111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_5_10_1  (
            .in0(N__12598),
            .in1(N__14159),
            .in2(N__12523),
            .in3(N__14682),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOut_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_5_10_2 .LUT_INIT=16'b0000101001011111;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_5_10_2  (
            .in0(N__12695),
            .in1(_gnd_net_),
            .in2(N__12738),
            .in3(N__12735),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22792),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_1_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_1_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_1_LC_5_10_3 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI_1_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__14221),
            .in2(_gnd_net_),
            .in3(N__14189),
            .lcout(\Lab_UT.alarmchar_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_10_4 .LUT_INIT=16'b0010001000111111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_5_10_4  (
            .in0(N__14160),
            .in1(N__12599),
            .in2(N__15528),
            .in3(N__12502),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOut_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_5_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_5_10_5 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(N__12696),
            .in2(N__12630),
            .in3(N__12627),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22792),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_5_10_7 .LUT_INIT=16'b0001101100010001;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_5_10_7  (
            .in0(N__12597),
            .in1(N__12531),
            .in2(N__12522),
            .in3(N__14607),
            .lcout(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_5_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_5_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__18666),
            .in2(_gnd_net_),
            .in3(N__17563),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m1_0_LC_5_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m1_0_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m1_0_LC_5_11_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m1_0_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(N__18667),
            .in2(_gnd_net_),
            .in3(N__17564),
            .lcout(\Lab_UT.dictrl.alarmstate8_2_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_2_LC_5_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_2_LC_5_11_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_2_LC_5_11_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_2_LC_5_11_4  (
            .in0(N__18669),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22788),
            .ce(N__15606),
            .sr(N__22520));
    defparam \Lab_UT.dictrl.shifter_ret_1_LC_5_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_1_LC_5_11_5 .SEQ_MODE=4'b1011;
    defparam \Lab_UT.dictrl.shifter_ret_1_LC_5_11_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_1_LC_5_11_5  (
            .in0(_gnd_net_),
            .in1(N__18668),
            .in2(_gnd_net_),
            .in3(N__17565),
            .lcout(\Lab_UT.dictrl.alarmstate8_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22788),
            .ce(N__15606),
            .sr(N__22520));
    defparam \buart.Z_rx.shifter_0_3_LC_5_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_3_LC_5_11_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_3_LC_5_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_3_LC_5_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21063),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22788),
            .ce(N__15606),
            .sr(N__22520));
    defparam \buart.Z_rx.shifter_ret_2_LC_5_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_2_LC_5_11_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_2_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_2_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17566),
            .lcout(bu_rx_data_i_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22788),
            .ce(N__15606),
            .sr(N__22520));
    defparam \buart.Z_rx.shifter_ret_LC_5_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_LC_5_12_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_LC_5_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_LC_5_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20799),
            .lcout(bu_rx_data_i_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22784),
            .ce(N__15604),
            .sr(N__22523));
    defparam \resetGen.escKey_4_LC_5_13_1 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_5_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \resetGen.escKey_4_LC_5_13_1  (
            .in0(N__21069),
            .in1(N__18154),
            .in2(N__20833),
            .in3(N__18695),
            .lcout(\resetGen.escKeyZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_6_rep1_LC_5_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_6_rep1_LC_5_13_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_6_rep1_LC_5_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_6_rep1_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21072),
            .lcout(bu_rx_data_i_4_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__15602),
            .sr(N__22525));
    defparam \buart.Z_rx.shifter_ret_6_fast_LC_5_13_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_6_fast_LC_5_13_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_6_fast_LC_5_13_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_6_fast_LC_5_13_3  (
            .in0(N__21071),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_4_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__15602),
            .sr(N__22525));
    defparam \buart.Z_rx.shifter_0_fast_3_LC_5_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_3_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_3_LC_5_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_3_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21073),
            .lcout(buart__rx_shifter_0_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__15602),
            .sr(N__22525));
    defparam \buart.Z_rx.shifter_ret_6_LC_5_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_6_LC_5_13_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_6_LC_5_13_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_6_LC_5_13_5  (
            .in0(N__21070),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__15602),
            .sr(N__22525));
    defparam \buart.Z_rx.shifter_0_1_LC_5_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_1_LC_5_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_1_LC_5_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_1_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17596),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__15602),
            .sr(N__22525));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_13_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_13_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_13_7  (
            .in0(N__12887),
            .in1(N__12821),
            .in2(N__12860),
            .in3(N__12912),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_5_14_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_5_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__12891),
            .in2(N__12864),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_5_14_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_5_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12924),
            .in3(N__12825),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__22776),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_5_14_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_5_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_5_14_2  (
            .in0(N__12800),
            .in1(N__12822),
            .in2(_gnd_net_),
            .in3(N__12810),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__22776),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_5_14_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_5_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12768),
            .in3(N__12807),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__22776),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_5_14_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_5_14_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_5_14_4  (
            .in0(N__12801),
            .in1(_gnd_net_),
            .in2(N__12780),
            .in3(N__12804),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__22776),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_5_14_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_5_14_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_5_14_5  (
            .in0(N__12755),
            .in1(N__12799),
            .in2(_gnd_net_),
            .in3(N__12783),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22776),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_5_14_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_5_14_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNIHV38_6_LC_5_14_6  (
            .in0(N__12776),
            .in1(N__12764),
            .in2(N__12756),
            .in3(N__12920),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNICJDT_1_LC_6_1_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNICJDT_1_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNICJDT_1_LC_6_1_1 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNICJDT_1_LC_6_1_1  (
            .in0(N__15377),
            .in1(N__14023),
            .in2(N__13987),
            .in3(N__15457),
            .lcout(\Lab_UT.didp.did_alarmMatch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14459),
            .in3(N__15378),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_1_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_1_3 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_1_3  (
            .in0(N__17834),
            .in1(N__18729),
            .in2(N__12906),
            .in3(N__15428),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_1_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_1_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_6_1_4  (
            .in0(N__15930),
            .in1(N__15429),
            .in2(N__12903),
            .in3(N__14445),
            .lcout(\Lab_UT.didp.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22835),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_6_1_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_6_1_6 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_6_1_6  (
            .in0(N__15394),
            .in1(N__17833),
            .in2(N__14460),
            .in3(N__17634),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_6_1_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_6_1_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_6_1_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_6_1_7  (
            .in0(N__14444),
            .in1(N__15929),
            .in2(N__12900),
            .in3(N__15395),
            .lcout(\Lab_UT.didp.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22835),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_2_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_6_2_0 .LUT_INIT=16'b0000111000000001;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_6_2_0  (
            .in0(N__15776),
            .in1(N__16248),
            .in2(N__16281),
            .in3(N__12897),
            .lcout(\Lab_UT.didp.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22825),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_2_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_6_2_1  (
            .in0(N__15858),
            .in1(N__15772),
            .in2(_gnd_net_),
            .in3(N__18214),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNINAVN_0_LC_6_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNINAVN_0_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNINAVN_0_LC_6_2_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNINAVN_0_LC_6_2_2  (
            .in0(_gnd_net_),
            .in1(N__13911),
            .in2(_gnd_net_),
            .in3(N__15857),
            .lcout(),
            .ltout(\Lab_UT.didp.un2_did_alarmMatch_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNIOMK62_0_LC_6_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNIOMK62_0_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNIOMK62_0_LC_6_2_3 .LUT_INIT=16'b0000100100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNIOMK62_0_LC_6_2_3  (
            .in0(N__15227),
            .in1(N__14834),
            .in2(N__13047),
            .in3(N__12969),
            .lcout(\Lab_UT.didp.regrce4.did_alarmMatch_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_6_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_6_2_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_1_LC_6_2_4  (
            .in0(N__20886),
            .in1(N__15902),
            .in2(N__15786),
            .in3(N__15859),
            .lcout(\Lab_UT.didp.countrce3.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNI0LVO3_0_LC_6_3_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNI0LVO3_0_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNI0LVO3_0_LC_6_3_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNI0LVO3_0_LC_6_3_0  (
            .in0(N__14944),
            .in1(N__17795),
            .in2(N__15048),
            .in3(N__13588),
            .lcout(\Lab_UT.sec2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIR0LH1_LC_6_3_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIR0LH1_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNIR0LH1_LC_6_3_1 .LUT_INIT=16'b1100111111011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNIR0LH1_LC_6_3_1  (
            .in0(N__16764),
            .in1(N__20345),
            .in2(N__18024),
            .in3(N__16547),
            .lcout(\Lab_UT.loadalarm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_RNIITJO1_LC_6_3_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNIITJO1_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNIITJO1_LC_6_3_2 .LUT_INIT=16'b1111010111110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNIITJO1_LC_6_3_2  (
            .in0(N__22242),
            .in1(N__14770),
            .in2(N__20368),
            .in3(N__16765),
            .lcout(\Lab_UT.loadalarm_0_0 ),
            .ltout(\Lab_UT.loadalarm_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI2VJT3_0_LC_6_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI2VJT3_0_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI2VJT3_0_LC_6_3_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI2VJT3_0_LC_6_3_3  (
            .in0(N__14664),
            .in1(N__17472),
            .in2(N__13008),
            .in3(N__15030),
            .lcout(\Lab_UT.sec1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_RNI8N121_0_LC_6_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_RNI8N121_0_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_RNI8N121_0_LC_6_3_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce1.q_RNI8N121_0_LC_6_3_4  (
            .in0(N__13587),
            .in1(N__17471),
            .in2(N__14671),
            .in3(N__17794),
            .lcout(\Lab_UT.didp.did_alarmMatch_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNIANSM3_2_LC_6_3_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNIANSM3_2_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNIANSM3_2_LC_6_3_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNIANSM3_2_LC_6_3_7  (
            .in0(N__14960),
            .in1(N__14423),
            .in2(N__14733),
            .in3(N__15031),
            .lcout(\Lab_UT.min1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_6_LC_6_4_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_6_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_6_LC_6_4_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_6_LC_6_4_0  (
            .in0(N__13380),
            .in1(N__13246),
            .in2(N__12963),
            .in3(N__13476),
            .lcout(),
            .ltout(\uu2.o_adder_vbuf_w_addr_displaying_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_6_LC_6_4_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_6_4_1 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_6_4_1 .LUT_INIT=16'b1111101011110000;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_6_4_1  (
            .in0(N__13815),
            .in1(_gnd_net_),
            .in2(N__13551),
            .in3(N__13424),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_ness_6C_net ),
            .ce(N__13547),
            .sr(N__22484));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_6_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_6_4_2 .LUT_INIT=16'b0000001101001000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_6_4_2  (
            .in0(N__13377),
            .in1(N__13311),
            .in2(N__13251),
            .in3(N__13813),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_6_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_6_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_6_4_3  (
            .in0(N__13312),
            .in1(N__13475),
            .in2(N__13253),
            .in3(N__13378),
            .lcout(\uu2.un15_w_data_displaying_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_6_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_6_4_4 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_6_4_4  (
            .in0(N__13379),
            .in1(N__13313),
            .in2(N__13252),
            .in3(N__13814),
            .lcout(\uu2.bitmap_pmux_sn_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_290_LC_6_5_0 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_6_5_0 .LUT_INIT=16'b0000011000011011;
    LogicCell40 \uu2.bitmap_290_LC_6_5_0  (
            .in0(N__14533),
            .in1(N__13862),
            .in2(N__14900),
            .in3(N__14565),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__22481));
    defparam \uu2.bitmap_194_LC_6_5_1 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_6_5_1 .LUT_INIT=16'b0001000100000101;
    LogicCell40 \uu2.bitmap_194_LC_6_5_1  (
            .in0(N__14562),
            .in1(N__14888),
            .in2(N__13871),
            .in3(N__14535),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__22481));
    defparam \uu2.bitmap_66_LC_6_5_2 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_6_5_2 .LUT_INIT=16'b0001010000011101;
    LogicCell40 \uu2.bitmap_66_LC_6_5_2  (
            .in0(N__14534),
            .in1(N__13863),
            .in2(N__14901),
            .in3(N__14566),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__22481));
    defparam \uu2.bitmap_RNIV8902_66_LC_6_5_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIV8902_66_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIV8902_66_LC_6_5_3 .LUT_INIT=16'b0011001111100010;
    LogicCell40 \uu2.bitmap_RNIV8902_66_LC_6_5_3  (
            .in0(N__13200),
            .in1(N__13194),
            .in2(N__13188),
            .in3(N__13150),
            .lcout(\uu2.bitmap_RNIV8902Z0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_6_5_4 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_6_5_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_162_LC_6_5_4  (
            .in0(N__14532),
            .in1(N__13861),
            .in2(N__14899),
            .in3(N__14564),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__22481));
    defparam \uu2.bitmap_34_LC_6_5_5 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_6_5_5 .LUT_INIT=16'b1111011101101101;
    LogicCell40 \uu2.bitmap_34_LC_6_5_5  (
            .in0(N__14563),
            .in1(N__14889),
            .in2(N__13872),
            .in3(N__14536),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__22481));
    defparam \uu2.bitmap_RNIEJM91_34_LC_6_5_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIEJM91_34_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIEJM91_34_LC_6_5_6 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \uu2.bitmap_RNIEJM91_34_LC_6_5_6  (
            .in0(N__13833),
            .in1(N__13805),
            .in2(N__13749),
            .in3(N__13700),
            .lcout(\uu2.bitmap_pmux_26_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_5_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI6RO21_162_LC_6_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNI6RO21_162_LC_6_5_7  (
            .in0(N__13699),
            .in1(N__13629),
            .in2(_gnd_net_),
            .in3(N__13620),
            .lcout(\uu2.N_217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_6_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__14690),
            .in2(_gnd_net_),
            .in3(N__14413),
            .lcout(\Lab_UT.didp.countrce4.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNIOF7P_1_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNIOF7P_1_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNIOF7P_1_LC_6_6_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNIOF7P_1_LC_6_6_3  (
            .in0(N__16159),
            .in1(N__14715),
            .in2(N__14422),
            .in3(N__14793),
            .lcout(),
            .ltout(\Lab_UT.didp.regrce4.did_alarmMatch_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNIGCKQ8_0_LC_6_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNIGCKQ8_0_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNIGCKQ8_0_LC_6_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNIGCKQ8_0_LC_6_6_4  (
            .in0(N__15099),
            .in1(N__14343),
            .in2(N__13605),
            .in3(N__13602),
            .lcout(\Lab_UT.alarmMatch ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_6_5 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_6_6_5  (
            .in0(N__14414),
            .in1(N__15173),
            .in2(N__14694),
            .in3(N__17620),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_6_6_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_6_6_6  (
            .in0(N__16086),
            .in1(N__15141),
            .in2(N__13593),
            .in3(N__14415),
            .lcout(\Lab_UT.didp.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22800),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_0_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_0_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_0_LC_6_7_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce1.q_0_LC_6_7_0  (
            .in0(N__18200),
            .in1(N__16548),
            .in2(N__13590),
            .in3(N__16436),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce1.q_1_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_1_LC_6_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_1_LC_6_7_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_1_LC_6_7_1  (
            .in0(N__16549),
            .in1(N__20878),
            .in2(N__16450),
            .in3(N__14022),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce1.q_2_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_2_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_2_LC_6_7_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce1.q_2_LC_6_7_2  (
            .in0(N__17615),
            .in1(N__16550),
            .in2(N__13986),
            .in3(N__16440),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce1.q_3_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_3_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_3_LC_6_7_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_3_LC_6_7_3  (
            .in0(N__16551),
            .in1(N__18718),
            .in2(N__16451),
            .in3(N__13936),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce3.q_0_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_0_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_0_LC_6_7_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_0_LC_6_7_4  (
            .in0(N__18201),
            .in1(N__16762),
            .in2(N__13914),
            .in3(N__16444),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce3.q_3_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_3_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_3_LC_6_7_5 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_3_LC_6_7_5  (
            .in0(N__16761),
            .in1(N__18719),
            .in2(N__16452),
            .in3(N__14493),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.didp.regrce3.q_2_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_2_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_2_LC_6_7_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_2_LC_6_7_6  (
            .in0(N__17616),
            .in1(N__16763),
            .in2(N__14387),
            .in3(N__16445),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22796),
            .ce(),
            .sr(N__22498));
    defparam \Lab_UT.dictrl.g0_9_1_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_9_1_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_9_1_LC_6_8_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.g0_9_1_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__18707),
            .in2(_gnd_net_),
            .in3(N__17600),
            .lcout(\Lab_UT.dictrl.g0_9Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIR2IE1_2_LC_6_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR2IE1_2_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR2IE1_2_LC_6_8_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIR2IE1_2_LC_6_8_7  (
            .in0(N__20175),
            .in1(N__16993),
            .in2(_gnd_net_),
            .in3(N__21386),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_0_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_0_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_0_LC_6_9_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_0_LC_6_9_0  (
            .in0(N__19645),
            .in1(N__14185),
            .in2(_gnd_net_),
            .in3(N__14214),
            .lcout(\Lab_UT.dictrl.alarmstate_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIMIM09_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIMIM09_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIMIM09_LC_6_9_1 .LUT_INIT=16'b0000010000100110;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNIMIM09_LC_6_9_1  (
            .in0(N__14186),
            .in1(N__14112),
            .in2(N__14223),
            .in3(N__14148),
            .lcout(\Lab_UT.dictrl.alarmstate_1_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIGCKQ8_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIGCKQ8_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIGCKQ8_LC_6_9_2 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNIGCKQ8_LC_6_9_2  (
            .in0(N__14147),
            .in1(N__14219),
            .in2(N__14058),
            .in3(N__14188),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIK5FS8_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIK5FS8_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIK5FS8_LC_6_9_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNIK5FS8_LC_6_9_3  (
            .in0(N__14220),
            .in1(N__14085),
            .in2(N__14097),
            .in3(N__14091),
            .lcout(\Lab_UT.shifter_ret_3_RNIK5FS8_0 ),
            .ltout(\Lab_UT.shifter_ret_3_RNIK5FS8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_LC_6_9_4 .LUT_INIT=16'b1010111111111111;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI4PQ1_LC_6_9_4  (
            .in0(N__19644),
            .in1(_gnd_net_),
            .in2(N__14094),
            .in3(N__14184),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i ),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIQBH29_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIQBH29_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNIQBH29_LC_6_9_5 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNIQBH29_LC_6_9_5  (
            .in0(N__14187),
            .in1(N__14084),
            .in2(N__14076),
            .in3(N__14073),
            .lcout(\Lab_UT.shifter_ret_3_RNIQBH29_0 ),
            .ltout(\Lab_UT.shifter_ret_3_RNIQBH29_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_2_LC_6_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_2_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_2_LC_6_9_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI_2_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14067),
            .in3(N__14218),
            .lcout(\Lab_UT.trig ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI6H8A1_2_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI6H8A1_2_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI6H8A1_2_LC_6_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI6H8A1_2_LC_6_9_7  (
            .in0(N__21387),
            .in1(N__16449),
            .in2(_gnd_net_),
            .in3(N__20176),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_6_10_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_6_10_0  (
            .in0(N__20359),
            .in1(N__14256),
            .in2(N__14247),
            .in3(N__14064),
            .lcout(\Lab_UT.dictrl.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI6626_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI6626_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI6626_LC_6_10_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI6626_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__14108),
            .in2(_gnd_net_),
            .in3(N__14231),
            .lcout(\Lab_UT.dictrl.N_127_0_0 ),
            .ltout(\Lab_UT.dictrl.N_127_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNI_LC_6_10_2 .LUT_INIT=16'b1111111110100010;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNI_LC_6_10_2  (
            .in0(N__14232),
            .in1(N__14049),
            .in2(N__14235),
            .in3(N__14127),
            .lcout(\Lab_UT.dictrl.justentered_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.m9_LC_6_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.m9_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.m9_LC_6_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dispString.m9_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__14222),
            .in2(_gnd_net_),
            .in3(N__14190),
            .lcout(\Lab_UT.armed ),
            .ltout(\Lab_UT.armed_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_10_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14151),
            .in3(N__14146),
            .lcout(G_203),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_5_LC_6_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_5_LC_6_11_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_5_LC_6_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_5_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21532),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \buart.Z_rx.shifter_0_7_LC_6_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_7_LC_6_11_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_7_LC_6_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_7_LC_6_11_1  (
            .in0(N__19473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \buart.Z_rx.shifter_0_6_LC_6_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_6_LC_6_11_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_6_LC_6_11_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_0_6_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__14271),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \Lab_UT.dictrl.shifter_ret_3_RNO_0_LC_6_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNO_0_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_3_RNO_0_LC_6_11_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_RNO_0_LC_6_11_3  (
            .in0(N__20967),
            .in1(N__21062),
            .in2(N__14274),
            .in3(N__20851),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate8_10_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_3_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_3_LC_6_11_4 .SEQ_MODE=4'b1010;
    defparam \Lab_UT.dictrl.shifter_ret_3_LC_6_11_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_3_LC_6_11_4  (
            .in0(N__14121),
            .in1(N__19472),
            .in2(N__14115),
            .in3(N__21531),
            .lcout(\Lab_UT.dictrl.alarmstate8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \buart.Z_rx.shifter_0_4_LC_6_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_4_LC_6_11_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_4_LC_6_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_4_LC_6_11_5  (
            .in0(N__20968),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \buart.Z_rx.shifter_0_fast_6_LC_6_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_6_LC_6_11_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_6_LC_6_11_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \buart.Z_rx.shifter_0_fast_6_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__14273),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \buart.Z_rx.shifter_0_6_rep1_LC_6_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_6_rep1_LC_6_11_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_6_rep1_LC_6_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_6_rep1_LC_6_11_7  (
            .in0(N__14272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22781),
            .ce(N__15605),
            .sr(N__22524));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_6_12_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_6_LC_6_12_0  (
            .in0(N__21530),
            .in1(N__20962),
            .in2(N__22269),
            .in3(N__21385),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_5_fast_LC_6_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_5_fast_LC_6_12_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_5_fast_LC_6_12_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_5_fast_LC_6_12_1  (
            .in0(N__20964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_ret_5_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22778),
            .ce(N__15603),
            .sr(N__22526));
    defparam \buart.Z_rx.shifter_0_fast_4_LC_6_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_4_LC_6_12_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_4_LC_6_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_4_LC_6_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20966),
            .lcout(bu_rx_data_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22778),
            .ce(N__15603),
            .sr(N__22526));
    defparam \buart.Z_rx.shifter_ret_5_LC_6_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_5_LC_6_12_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_5_LC_6_12_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_5_LC_6_12_3  (
            .in0(N__20963),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22778),
            .ce(N__15603),
            .sr(N__22526));
    defparam \buart.Z_rx.shifter_0_4_rep1_LC_6_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_4_rep1_LC_6_12_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_4_rep1_LC_6_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_4_rep1_LC_6_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20965),
            .lcout(bu_rx_data_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22778),
            .ce(N__15603),
            .sr(N__22526));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_6_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_7_LC_6_12_5  (
            .in0(N__21656),
            .in1(N__21430),
            .in2(N__17078),
            .in3(N__21698),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_0_LC_6_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_0_LC_6_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_0_LC_6_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_0_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20800),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22778),
            .ce(N__15603),
            .sr(N__22526));
    defparam \Lab_UT.dictrl.g0_31_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_31_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_31_LC_6_13_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_31_LC_6_13_0  (
            .in0(N__17380),
            .in1(N__17192),
            .in2(N__17277),
            .in3(N__17342),
            .lcout(\Lab_UT.dictrl.N_98_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m40_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m40_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m40_LC_6_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.m40_LC_6_13_2  (
            .in0(N__17379),
            .in1(N__17275),
            .in2(N__14313),
            .in3(N__17193),
            .lcout(\Lab_UT.dictrl.N_99_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_1_4_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_4_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_4_LC_6_13_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \Lab_UT.dictrl.g1_1_4_LC_6_13_3  (
            .in0(N__14319),
            .in1(N__17271),
            .in2(N__14312),
            .in3(N__17378),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_1_RNICGMV1_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_1_RNICGMV1_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_1_RNICGMV1_LC_6_13_4 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_1_RNICGMV1_LC_6_13_4  (
            .in0(N__17147),
            .in1(N__21544),
            .in2(N__14295),
            .in3(N__18137),
            .lcout(\Lab_UT.dictrl.g1_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_5_rep1_LC_6_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_5_rep1_LC_6_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_5_rep1_LC_6_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_5_rep1_LC_6_13_5  (
            .in0(N__21545),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22775),
            .ce(N__15601),
            .sr(N__22527));
    defparam \buart.Z_rx.shifter_0_fast_5_LC_6_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_5_LC_6_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_5_LC_6_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_fast_5_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21546),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22775),
            .ce(N__15601),
            .sr(N__22527));
    defparam \Lab_UT.dictrl.g0_43_x_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_43_x_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_43_x_LC_6_13_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_43_x_LC_6_13_7  (
            .in0(N__17311),
            .in1(N__17270),
            .in2(_gnd_net_),
            .in3(N__15344),
            .lcout(\Lab_UT.dictrl.g0_43_xZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_6_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_15_LC_6_14_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_15_LC_6_14_3  (
            .in0(N__15351),
            .in1(N__17234),
            .in2(N__15642),
            .in3(N__17307),
            .lcout(\Lab_UT.dictrl.N_98_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_20_LC_6_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_20_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_20_LC_6_14_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.g0_20_LC_6_14_4  (
            .in0(N__15677),
            .in1(N__15318),
            .in2(N__14292),
            .in3(N__20779),
            .lcout(\Lab_UT.dictrl.N_88_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_6_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_14_LC_6_14_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_14_LC_6_14_6  (
            .in0(N__17306),
            .in1(N__15350),
            .in2(_gnd_net_),
            .in3(N__20641),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_6_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_11_LC_6_14_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_11_LC_6_14_7  (
            .in0(N__20780),
            .in1(N__14283),
            .in2(N__14277),
            .in3(N__15678),
            .lcout(\Lab_UT.dictrl.N_88_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_1_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_1_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_1_1  (
            .in0(N__20887),
            .in1(N__15462),
            .in2(N__17835),
            .in3(N__17791),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_1_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_7_1_2  (
            .in0(N__15463),
            .in1(N__15923),
            .in2(N__14463),
            .in3(N__14443),
            .lcout(\Lab_UT.didp.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22847),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNIVHJJ_1_LC_7_1_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNIVHJJ_1_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNIVHJJ_1_LC_7_1_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNIVHJJ_1_LC_7_1_3  (
            .in0(_gnd_net_),
            .in1(N__15461),
            .in2(_gnd_net_),
            .in3(N__17790),
            .lcout(\Lab_UT.didp.countrce1.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI65GA_0_LC_7_1_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI65GA_0_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI65GA_0_LC_7_1_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI65GA_0_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(N__14853),
            .in2(_gnd_net_),
            .in3(N__17709),
            .lcout(\Lab_UT.didp.un1_dicLdSones_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdSones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_1_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_1_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_1_6 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_7_1_6  (
            .in0(N__17792),
            .in1(N__15922),
            .in2(N__14430),
            .in3(N__17760),
            .lcout(\Lab_UT.didp.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22847),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_7_2_1  (
            .in0(N__15228),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14427),
            .lcout(\Lab_UT.didp.reset_12_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_7_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_7_2_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_7_2_3  (
            .in0(N__15895),
            .in1(N__14383),
            .in2(N__15823),
            .in3(N__14584),
            .lcout(\Lab_UT.didp.did_alarmMatch_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI14UL1_2_LC_7_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI14UL1_2_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI14UL1_2_LC_7_2_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.didp.ce_RNI14UL1_2_LC_7_2_4  (
            .in0(N__16241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15789),
            .lcout(\Lab_UT.didp.un1_dicLdMones_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_2_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_7_2_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_7_2_5  (
            .in0(N__15896),
            .in1(N__16270),
            .in2(N__14331),
            .in3(N__14328),
            .lcout(\Lab_UT.didp.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22839),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_0_LC_7_3_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_0_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_0_LC_7_3_0 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_0_LC_7_3_0  (
            .in0(N__18215),
            .in1(N__16768),
            .in2(N__14681),
            .in3(N__17026),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce2.q_1_LC_7_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_1_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_1_LC_7_3_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_1_LC_7_3_1  (
            .in0(N__16766),
            .in1(N__20876),
            .in2(N__17036),
            .in3(N__15558),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce2.q_2_LC_7_3_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_2_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_2_LC_7_3_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_2_LC_7_3_2  (
            .in0(N__17635),
            .in1(N__16769),
            .in2(N__15516),
            .in3(N__17030),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce2.q_3_LC_7_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_3_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_3_LC_7_3_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_3_LC_7_3_3  (
            .in0(N__16767),
            .in1(N__18740),
            .in2(N__17037),
            .in3(N__14626),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce3.q_1_LC_7_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_1_LC_7_3_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_1_LC_7_3_4 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_1_LC_7_3_4  (
            .in0(N__20875),
            .in1(N__16770),
            .in2(N__16417),
            .in3(N__14590),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce4.q_3_LC_7_3_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_3_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_3_LC_7_3_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \Lab_UT.didp.regrce4.q_3_LC_7_3_5  (
            .in0(N__17025),
            .in1(N__14771),
            .in2(N__15089),
            .in3(N__18741),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22504));
    defparam \Lab_UT.didp.regrce4.q_RNI6JSM3_0_LC_7_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNI6JSM3_0_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNI6JSM3_0_LC_7_4_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNI6JSM3_0_LC_7_4_0  (
            .in0(N__15225),
            .in1(N__14953),
            .in2(N__15049),
            .in3(N__14829),
            .lcout(\Lab_UT.min1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNI8LSM3_1_LC_7_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNI8LSM3_1_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNI8LSM3_1_LC_7_4_1 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNI8LSM3_1_LC_7_4_1  (
            .in0(N__14954),
            .in1(N__16171),
            .in2(N__15050),
            .in3(N__14794),
            .lcout(\Lab_UT.min1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNISBJ41_3_LC_7_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNISBJ41_3_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNISBJ41_3_LC_7_4_2 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNISBJ41_3_LC_7_4_2  (
            .in0(N__14503),
            .in1(N__15725),
            .in2(N__16129),
            .in3(N__15078),
            .lcout(),
            .ltout(\Lab_UT.didp.regrce4.did_alarmMatch_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNICAPA4_3_LC_7_4_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNICAPA4_3_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNICAPA4_3_LC_7_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNICAPA4_3_LC_7_4_3  (
            .in0(N__15477),
            .in1(N__15126),
            .in2(N__15114),
            .in3(N__15111),
            .lcout(\Lab_UT.didp.regrce4.did_alarmMatch_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_RNICPSM3_3_LC_7_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_RNICPSM3_3_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_RNICPSM3_3_LC_7_4_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_RNICPSM3_3_LC_7_4_5  (
            .in0(N__15079),
            .in1(N__15035),
            .in2(N__16130),
            .in3(N__14961),
            .lcout(\Lab_UT.min1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_5_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_5_0 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_7_5_0  (
            .in0(N__14763),
            .in1(N__17722),
            .in2(N__22596),
            .in3(N__19947),
            .lcout(\Lab_UT.dicRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22819),
            .ce(),
            .sr(N__22501));
    defparam \Lab_UT.didp.ce_0_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_7_5_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_7_5_1  (
            .in0(N__16012),
            .in1(N__14766),
            .in2(_gnd_net_),
            .in3(N__16407),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22819),
            .ce(),
            .sr(N__22501));
    defparam \Lab_UT.didp.regrce4.q_0_LC_7_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_0_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_0_LC_7_5_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_0_LC_7_5_2  (
            .in0(N__14764),
            .in1(N__18226),
            .in2(N__17034),
            .in3(N__14833),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22819),
            .ce(),
            .sr(N__22501));
    defparam \Lab_UT.didp.regrce4.q_1_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_1_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_1_LC_7_5_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_1_LC_7_5_3  (
            .in0(N__14798),
            .in1(N__20877),
            .in2(N__14772),
            .in3(N__17021),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22819),
            .ce(),
            .sr(N__22501));
    defparam \Lab_UT.didp.regrce4.q_2_LC_7_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_2_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_2_LC_7_5_4 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_2_LC_7_5_4  (
            .in0(N__14765),
            .in1(N__17633),
            .in2(N__17035),
            .in3(N__14722),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22819),
            .ce(),
            .sr(N__22501));
    defparam \Lab_UT.didp.countrce4.q_RNI5GGH_0_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNI5GGH_0_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNI5GGH_0_LC_7_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNI5GGH_0_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__15214),
            .in2(_gnd_net_),
            .in3(N__16163),
            .lcout(\Lab_UT.didp.countrce4.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_6_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_6_1  (
            .in0(N__15215),
            .in1(N__15170),
            .in2(_gnd_net_),
            .in3(N__18225),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_7_6_2 .LUT_INIT=16'b0000000011100001;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_7_6_2  (
            .in0(N__15696),
            .in1(N__15174),
            .in2(N__15231),
            .in3(N__16080),
            .lcout(\Lab_UT.didp.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22812),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_6_3 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_6_3  (
            .in0(N__16164),
            .in1(N__15171),
            .in2(N__15226),
            .in3(N__20888),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_6_4 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_7_6_4  (
            .in0(N__16175),
            .in1(N__15139),
            .in2(N__15186),
            .in3(N__16081),
            .lcout(\Lab_UT.didp.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22812),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_6_5 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_7_6_5  (
            .in0(N__15183),
            .in1(N__18720),
            .in2(N__16128),
            .in3(N__15172),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_7_6_6 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_7_6_6  (
            .in0(N__16118),
            .in1(N__16082),
            .in2(N__15177),
            .in3(N__15140),
            .lcout(\Lab_UT.didp.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22812),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_7_6_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNIDJKH1_3_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__15695),
            .in2(_gnd_net_),
            .in3(N__15169),
            .lcout(\Lab_UT.didp.un1_dicLdMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_7_7_0 .C_ON=1'b0;
    defparam \resetGen.rst_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_7_7_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16481),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22804),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIE8RP4_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIE8RP4_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIE8RP4_LC_7_7_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIE8RP4_LC_7_7_1  (
            .in0(N__19889),
            .in1(N__16881),
            .in2(_gnd_net_),
            .in3(N__22093),
            .lcout(\Lab_UT.dictrl.N_121_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_0_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_0_LC_7_7_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_0_LC_7_7_4  (
            .in0(N__18882),
            .in1(N__19888),
            .in2(_gnd_net_),
            .in3(N__21120),
            .lcout(\Lab_UT.dictrl.g1_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_LC_7_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_LC_7_7_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNI31Q21_LC_7_7_7  (
            .in0(N__21121),
            .in1(_gnd_net_),
            .in2(N__19901),
            .in3(N__18883),
            .lcout(\Lab_UT.dictrl.g3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_27_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_27_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_27_LC_7_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_27_LC_7_8_0  (
            .in0(N__18536),
            .in1(N__16837),
            .in2(N__18223),
            .in3(N__18076),
            .lcout(\Lab_UT.dictrl.N_116_mux_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_LC_7_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_LC_7_8_1  (
            .in0(N__18077),
            .in1(N__16848),
            .in2(N__18224),
            .in3(N__18537),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_116_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_3_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_3_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_3_LC_7_8_2 .LUT_INIT=16'b0101010100011101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI4N0L4_3_LC_7_8_2  (
            .in0(N__20352),
            .in1(N__22201),
            .in2(N__15249),
            .in3(N__21359),
            .lcout(\Lab_UT.dictrl.N_1304_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI24TF4_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI24TF4_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI24TF4_LC_7_8_3 .LUT_INIT=16'b0010001101110011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNI24TF4_LC_7_8_3  (
            .in0(N__21357),
            .in1(N__20351),
            .in2(N__21146),
            .in3(N__15246),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1304_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_0_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_0_LC_7_8_4 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIQ1339_0_LC_7_8_4  (
            .in0(N__22199),
            .in1(N__22095),
            .in2(N__15240),
            .in3(N__21358),
            .lcout(\Lab_UT.dictrl.N_94_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNISK689_0_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNISK689_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNISK689_0_LC_7_8_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNISK689_0_LC_7_8_5  (
            .in0(N__22096),
            .in1(N__15237),
            .in2(N__21383),
            .in3(N__22200),
            .lcout(\Lab_UT.dictrl.N_94_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0_3_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0_3_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0_3_LC_7_9_1 .LUT_INIT=16'b0000101101001111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI4N0L4_0_3_LC_7_9_1  (
            .in0(N__21366),
            .in1(N__22262),
            .in2(N__20370),
            .in3(N__20469),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNI4N0L4_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_7_9_2 .LUT_INIT=16'b1100000001000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_7_9_2  (
            .in0(N__20879),
            .in1(N__21363),
            .in2(N__22268),
            .in3(N__20656),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNICSUJ_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNICSUJ_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNICSUJ_LC_7_9_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNICSUJ_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__19883),
            .in2(_gnd_net_),
            .in3(N__21149),
            .lcout(\Lab_UT.dicLdMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_7_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_7_LC_7_9_4 .LUT_INIT=16'b0011001101010011;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_7_LC_7_9_4  (
            .in0(N__20468),
            .in1(N__18288),
            .in2(N__21158),
            .in3(N__21364),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1304_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_7_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_5_LC_7_9_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_5_LC_7_9_5  (
            .in0(N__21365),
            .in1(N__21153),
            .in2(N__15273),
            .in3(N__22094),
            .lcout(\Lab_UT.dictrl.N_94_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIBHFL_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIBHFL_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIBHFL_LC_7_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIBHFL_LC_7_10_0  (
            .in0(N__21148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21355),
            .lcout(\Lab_UT.dictrl.m36_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIAUDM_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIAUDM_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIAUDM_LC_7_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIAUDM_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__18286),
            .in2(_gnd_net_),
            .in3(N__21722),
            .lcout(\Lab_UT.dictrl.m45_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_10_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_10_LC_7_10_3  (
            .in0(N__17112),
            .in1(N__18854),
            .in2(_gnd_net_),
            .in3(N__18287),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_8_LC_7_10_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_8_LC_7_10_4  (
            .in0(N__15270),
            .in1(N__15255),
            .in2(N__15258),
            .in3(N__21356),
            .lcout(\Lab_UT.dictrl.i9_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_9_LC_7_10_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_9_LC_7_10_7  (
            .in0(N__17049),
            .in1(N__15651),
            .in2(_gnd_net_),
            .in3(N__16828),
            .lcout(\Lab_UT.dictrl.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m25_4_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m25_4_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m25_4_LC_7_11_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m25_4_LC_7_11_0  (
            .in0(N__21699),
            .in1(N__17176),
            .in2(N__21431),
            .in3(N__15640),
            .lcout(\Lab_UT.dictrl.m25Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m25_0_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m25_0_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m25_0_LC_7_11_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.dictrl.m25_0_LC_7_11_1  (
            .in0(N__16943),
            .in1(_gnd_net_),
            .in2(N__17428),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.m25Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_fast_RNI13PI1_2_LC_7_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_RNI13PI1_2_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_0_fast_RNI13PI1_2_LC_7_11_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \buart.Z_rx.shifter_0_fast_RNI13PI1_2_LC_7_11_2  (
            .in0(N__18136),
            .in1(N__17420),
            .in2(N__18544),
            .in3(N__16944),
            .lcout(g0_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m25_x1_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m25_x1_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m25_x1_LC_7_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.m25_x1_LC_7_11_3  (
            .in0(N__16942),
            .in1(N__18532),
            .in2(N__17427),
            .in3(N__18135),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m25_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m25_ns_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m25_ns_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m25_ns_LC_7_11_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.m25_ns_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15294),
            .in3(N__18067),
            .lcout(\Lab_UT.dictrl.N_116_mux ),
            .ltout(\Lab_UT.dictrl.N_116_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNIB8OC4_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNIB8OC4_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_RNIB8OC4_LC_7_11_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_RNIB8OC4_LC_7_11_5  (
            .in0(N__19882),
            .in1(N__17973),
            .in2(N__15291),
            .in3(N__21354),
            .lcout(\Lab_UT.dictrl.N_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_11_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_11_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_11_LC_7_12_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_11_LC_7_12_0  (
            .in0(N__20946),
            .in1(N__21037),
            .in2(N__21540),
            .in3(N__21630),
            .lcout(\Lab_UT.dictrl.N_98_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_1_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_1_LC_7_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_1_LC_7_12_1  (
            .in0(N__20637),
            .in1(N__20945),
            .in2(_gnd_net_),
            .in3(N__21038),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_35_LC_7_12_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Lab_UT.dictrl.g0_35_LC_7_12_2  (
            .in0(N__20856),
            .in1(N__15680),
            .in2(N__15288),
            .in3(N__18561),
            .lcout(\Lab_UT.dictrl.g1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_7_12_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_7_12_3  (
            .in0(N__15285),
            .in1(N__20371),
            .in2(N__18576),
            .in3(N__21502),
            .lcout(\Lab_UT.dictrl.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_46_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_46_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_46_LC_7_12_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_46_LC_7_12_4  (
            .in0(N__20944),
            .in1(N__21036),
            .in2(N__21539),
            .in3(N__21629),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_98_mux_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_42_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_42_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_42_LC_7_12_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.g0_42_LC_7_12_5  (
            .in0(N__15357),
            .in1(N__15681),
            .in2(N__15276),
            .in3(N__20857),
            .lcout(\Lab_UT.dictrl.g1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_1_0_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_0_LC_7_12_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.g1_1_0_LC_7_12_6  (
            .in0(N__20943),
            .in1(N__21035),
            .in2(_gnd_net_),
            .in3(N__20636),
            .lcout(\Lab_UT.dictrl.g1_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_2_1_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_2_1_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_2_1_LC_7_12_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.g1_2_1_LC_7_12_7  (
            .in0(N__21631),
            .in1(N__20947),
            .in2(N__21560),
            .in3(N__21039),
            .lcout(\Lab_UT.dictrl.g1_2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_28_1_0_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_28_1_0_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_28_1_0_LC_7_13_0 .LUT_INIT=16'b0101111100110011;
    LogicCell40 \Lab_UT.dictrl.g0_28_1_0_LC_7_13_0  (
            .in0(N__17336),
            .in1(N__15343),
            .in2(N__15312),
            .in3(N__20801),
            .lcout(\Lab_UT.dictrl.g0_28_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_3_0_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_3_0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_3_0_LC_7_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_3_0_LC_7_13_1  (
            .in0(N__15311),
            .in1(N__17377),
            .in2(_gnd_net_),
            .in3(N__17338),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_3_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_3_LC_7_13_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.dictrl.g0_3_LC_7_13_2  (
            .in0(N__15327),
            .in1(N__15679),
            .in2(N__15321),
            .in3(N__20802),
            .lcout(\Lab_UT.dictrl.N_88_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_4_1_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_4_1_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_4_1_LC_7_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_4_1_LC_7_13_3  (
            .in0(N__15310),
            .in1(N__17376),
            .in2(_gnd_net_),
            .in3(N__17337),
            .lcout(\Lab_UT.dictrl.g0_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_13_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_1_fast_LC_7_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_1_fast_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18716),
            .lcout(buart__rx_shifter_ret_1_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22780),
            .ce(N__15600),
            .sr(N__22529));
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_fast_2_LC_7_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_fast_2_LC_7_13_5  (
            .in0(N__18717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buart__rx_shifter_0_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22780),
            .ce(N__15600),
            .sr(N__22529));
    defparam \buart.Z_rx.shifter_ret_1_LC_7_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_1_LC_7_13_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_1_LC_7_13_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_1_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18715),
            .lcout(bu_rx_data_i_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22780),
            .ce(N__15600),
            .sr(N__22529));
    defparam \Lab_UT.dictrl.m31_x0_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m31_x0_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m31_x0_LC_7_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.m31_x0_LC_7_13_7  (
            .in0(N__20632),
            .in1(N__17375),
            .in2(N__15641),
            .in3(N__17335),
            .lcout(\Lab_UT.dictrl.m31_xZ0Z0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m19_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m19_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m19_LC_7_14_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.m19_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__17232),
            .in2(_gnd_net_),
            .in3(N__15635),
            .lcout(\Lab_UT.dictrl.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_12_LC_7_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_12_LC_7_14_4  (
            .in0(N__15636),
            .in1(N__17233),
            .in2(N__17312),
            .in3(N__21436),
            .lcout(\Lab_UT.dictrl.g0_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_3_fast_LC_7_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_fast_LC_7_14_5 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_3_fast_LC_7_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_3_fast_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19470),
            .lcout(bu_rx_data_i_4_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22777),
            .ce(N__15599),
            .sr(N__22531));
    defparam \buart.Z_rx.shifter_ret_3_rep1_LC_7_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_rep1_LC_7_14_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_3_rep1_LC_7_14_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_3_rep1_LC_7_14_6  (
            .in0(N__19471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_i_4_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22777),
            .ce(N__15599),
            .sr(N__22531));
    defparam \buart.Z_rx.shifter_ret_3_LC_7_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_LC_7_14_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_3_LC_7_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_3_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19469),
            .lcout(bu_rx_data_i_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22777),
            .ce(N__15599),
            .sr(N__22531));
    defparam \buart.Z_rx.shifter_ret_4_LC_7_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_4_LC_7_15_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.shifter_ret_4_LC_7_15_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_rx.shifter_ret_4_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21571),
            .lcout(bu_rx_data_i_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22774),
            .ce(N__15598),
            .sr(N__22533));
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_1_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_1_1 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_1_1  (
            .in0(N__17503),
            .in1(N__15559),
            .in2(N__15517),
            .in3(N__17920),
            .lcout(\Lab_UT.didp.did_alarmMatch_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_1_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_1_2  (
            .in0(N__15464),
            .in1(N__15432),
            .in2(N__15396),
            .in3(N__17793),
            .lcout(\Lab_UT.didp.un18_ce ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_1_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_1_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_1_6  (
            .in0(N__17921),
            .in1(N__17675),
            .in2(N__17516),
            .in3(N__17470),
            .lcout(\Lab_UT.didp.un24_ce_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_2_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_2_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_2_0  (
            .in0(N__15867),
            .in1(N__15901),
            .in2(N__15825),
            .in3(N__15722),
            .lcout(\Lab_UT.didp.countrce3.ce_12_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_0_LC_8_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_0_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNI36SS_0_LC_8_2_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNI36SS_0_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__15900),
            .in2(_gnd_net_),
            .in3(N__15866),
            .lcout(\Lab_UT.didp.countrce3.un13_qPone ),
            .ltout(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_8_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_8_2_2 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_8_2_2  (
            .in0(N__15821),
            .in1(N__15787),
            .in2(N__15837),
            .in3(N__17636),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_8_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_8_2_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_8_2_3  (
            .in0(N__16280),
            .in1(N__15734),
            .in2(N__15834),
            .in3(N__15822),
            .lcout(\Lab_UT.didp.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22848),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_2_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_2_5  (
            .in0(_gnd_net_),
            .in1(N__15831),
            .in2(_gnd_net_),
            .in3(N__15820),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_2_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_2_6 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_2_6  (
            .in0(N__15788),
            .in1(N__18739),
            .in2(N__15741),
            .in3(N__15723),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_8_2_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_8_2_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_8_2_7  (
            .in0(N__15724),
            .in1(N__16269),
            .in2(N__15738),
            .in3(N__15735),
            .lcout(\Lab_UT.didp.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22848),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_1_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_8_3_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_8_3_0  (
            .in0(N__16030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16057),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.ce_3_LC_8_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_8_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_8_3_1  (
            .in0(N__16061),
            .in1(N__16229),
            .in2(N__16214),
            .in3(N__16035),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.reset_2_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_8_3_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_8_3_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_8_3_2  (
            .in0(N__16032),
            .in1(N__16062),
            .in2(N__16215),
            .in3(N__16230),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.ce_2_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_8_3_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_8_3_3  (
            .in0(N__16058),
            .in1(N__16209),
            .in2(_gnd_net_),
            .in3(N__16034),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.reset_1_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_8_3_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_8_3_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_8_3_4  (
            .in0(N__16031),
            .in1(N__16205),
            .in2(_gnd_net_),
            .in3(N__16060),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_3_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_3_5  (
            .in0(N__16056),
            .in1(N__16228),
            .in2(N__16213),
            .in3(N__16029),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_8_3_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_8_3_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_8_3_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_8_3_6  (
            .in0(N__16182),
            .in1(N__16176),
            .in2(N__16134),
            .in3(N__16131),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \Lab_UT.didp.reset_0_LC_8_3_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_8_3_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_8_3_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_8_3_7  (
            .in0(N__16059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16033),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22840),
            .ce(),
            .sr(N__22505));
    defparam \resetGen.reset_count_1_LC_8_4_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_8_4_0 .LUT_INIT=16'b0100010000010100;
    LogicCell40 \resetGen.reset_count_1_LC_8_4_0  (
            .in0(N__18480),
            .in1(N__16383),
            .in2(N__16368),
            .in3(N__16480),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_8_4_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_8_4_1 .LUT_INIT=16'b0000000010100101;
    LogicCell40 \resetGen.reset_count_0_LC_8_4_1  (
            .in0(N__16363),
            .in1(_gnd_net_),
            .in2(N__16482),
            .in3(N__18479),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_4_2 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__16382),
            .in2(_gnd_net_),
            .in3(N__16362),
            .lcout(\resetGen.un241_ci ),
            .ltout(\resetGen.un241_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_8_4_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_8_4_3 .LUT_INIT=16'b0000000010011100;
    LogicCell40 \resetGen.reset_count_2_LC_8_4_3  (
            .in0(N__16478),
            .in1(N__16340),
            .in2(N__16506),
            .in3(N__18481),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_8_4_4 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_8_4_4 .LUT_INIT=16'b0100000101010000;
    LogicCell40 \resetGen.reset_count_3_LC_8_4_4  (
            .in0(N__18482),
            .in1(N__16479),
            .in2(N__16503),
            .in3(N__16326),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_8_4_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_8_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__16499),
            .in2(_gnd_net_),
            .in3(N__16339),
            .lcout(),
            .ltout(\resetGen.reset_count_2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_8_4_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_8_4_6 .LUT_INIT=16'b0101010001000100;
    LogicCell40 \resetGen.reset_count_4_LC_8_4_6  (
            .in0(N__18483),
            .in1(N__16474),
            .in2(N__16491),
            .in3(N__16488),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNINALF_LC_8_4_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNINALF_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNINALF_LC_8_4_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNINALF_LC_8_4_7  (
            .in0(N__18020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20347),
            .lcout(\Lab_UT.dicRun_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_1_LC_8_5_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_8_5_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_8_5_0 .LUT_INIT=16'b0100011101110100;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_8_5_0  (
            .in0(N__22988),
            .in1(N__19404),
            .in2(N__19166),
            .in3(N__18048),
            .lcout(buart__rx_bitcount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22823),
            .ce(N__19349),
            .sr(N__22528));
    defparam \buart.Z_rx.bitcount_es_2_LC_8_5_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_8_5_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_8_5_1 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_8_5_1  (
            .in0(N__19403),
            .in1(N__22989),
            .in2(N__19200),
            .in3(N__18039),
            .lcout(buart__rx_bitcount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22823),
            .ce(N__19349),
            .sr(N__22528));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_8_5_2  (
            .in0(N__16381),
            .in1(N__16367),
            .in2(_gnd_net_),
            .in3(N__16341),
            .lcout(\resetGen.un252_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_RNILLLG7_1_LC_8_5_5 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_8_5_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_8_5_5  (
            .in0(N__16320),
            .in1(N__16296),
            .in2(_gnd_net_),
            .in3(N__16644),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_5_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_5_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_5_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_5_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ3CG_2_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ3CG_2_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ3CG_2_LC_8_6_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIQ3CG_2_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21951),
            .in3(N__20129),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIQ3CGZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJT2J_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJT2J_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJT2J_LC_8_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIJT2J_LC_8_6_2  (
            .in0(N__18000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20095),
            .lcout(\Lab_UT.dicLdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_1_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_1_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_1_LC_8_6_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUQEL8_1_LC_8_6_4  (
            .in0(N__16698),
            .in1(N__16683),
            .in2(N__16521),
            .in3(N__21298),
            .lcout(),
            .ltout(\Lab_UT.dictrl.i9_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIU0079_2_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIU0079_2_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIU0079_2_LC_8_6_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIU0079_2_LC_8_6_5  (
            .in0(N__21937),
            .in1(_gnd_net_),
            .in2(N__16512),
            .in3(N__19547),
            .lcout(\Lab_UT.dictrl.N_2000_0 ),
            .ltout(\Lab_UT.dictrl.N_2000_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKPIVI_2_LC_8_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKPIVI_2_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKPIVI_2_LC_8_6_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKPIVI_2_LC_8_6_6  (
            .in0(N__20128),
            .in1(N__16722),
            .in2(N__16509),
            .in3(N__21941),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIGJHP81_2_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIGJHP81_2_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIGJHP81_2_LC_8_7_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIGJHP81_2_LC_8_7_0  (
            .in0(N__18453),
            .in1(N__18432),
            .in2(N__21943),
            .in3(N__20130),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_7_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_7_1  (
            .in0(N__20132),
            .in1(N__21912),
            .in2(N__18441),
            .in3(N__18456),
            .lcout(\Lab_UT.dictrl.state_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22813),
            .ce(N__18249),
            .sr(N__22500));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_7_2 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_7_2  (
            .in0(N__18454),
            .in1(N__18433),
            .in2(N__21944),
            .in3(N__20133),
            .lcout(\Lab_UT.dictrl.state_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22813),
            .ce(N__18249),
            .sr(N__22500));
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_7_3 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_0_LC_8_7_3  (
            .in0(N__20131),
            .in1(N__21910),
            .in2(N__18440),
            .in3(N__18455),
            .lcout(\Lab_UT.dictrl.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22813),
            .ce(N__18249),
            .sr(N__22500));
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_7_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_7_4 .LUT_INIT=16'b0001101100001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_LC_8_7_4  (
            .in0(N__21913),
            .in1(N__19572),
            .in2(N__16788),
            .in3(N__20134),
            .lcout(\Lab_UT.dictrl.state_i_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22813),
            .ce(N__18249),
            .sr(N__22500));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIHOSE_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIHOSE_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIHOSE_LC_8_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNIHOSE_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__16776),
            .in2(_gnd_net_),
            .in3(N__21254),
            .lcout(\Lab_UT.dicLdAMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_7_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_2_LC_8_7_6  (
            .in0(N__21911),
            .in1(N__16718),
            .in2(N__20174),
            .in3(N__16704),
            .lcout(\Lab_UT.dictrl.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22813),
            .ce(N__18249),
            .sr(N__22500));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_LC_8_8_0 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_LC_8_8_0  (
            .in0(N__16847),
            .in1(_gnd_net_),
            .in2(N__20034),
            .in3(N__16866),
            .lcout(\Lab_UT.dictrl.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_0_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_0_LC_8_8_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIV6AH3_0_0_LC_8_8_1  (
            .in0(N__16865),
            .in1(N__20030),
            .in2(_gnd_net_),
            .in3(N__16846),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_0_1_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_0_1_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUQEL8_0_1_LC_8_8_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUQEL8_0_1_LC_8_8_2  (
            .in0(N__16689),
            .in1(N__16682),
            .in2(N__16659),
            .in3(N__21295),
            .lcout(),
            .ltout(\Lab_UT.dictrl.i9_mux_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIU0079_0_2_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIU0079_0_2_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIU0079_0_2_LC_8_8_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIU0079_0_2_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__19546),
            .in2(N__16656),
            .in3(N__21929),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_2000_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNII6FQI_2_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNII6FQI_2_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNII6FQI_2_LC_8_8_4 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNII6FQI_2_LC_8_8_4  (
            .in0(N__21930),
            .in1(N__16653),
            .in2(N__16647),
            .in3(N__20118),
            .lcout(Lab_UT_dictrl_next_state_0_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU5J2B_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU5J2B_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU5J2B_LC_8_9_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU5J2B_LC_8_9_0  (
            .in0(N__16994),
            .in1(N__16899),
            .in2(_gnd_net_),
            .in3(N__19026),
            .lcout(\Lab_UT.dictrl.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TO6_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TO6_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TO6_LC_8_9_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TO6_LC_8_9_3  (
            .in0(N__21157),
            .in1(N__19586),
            .in2(_gnd_net_),
            .in3(N__22091),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6 ),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIR1TOZ0Z6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIHF8LB_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIHF8LB_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIHF8LB_LC_8_9_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIHF8LB_LC_8_9_4  (
            .in0(N__18786),
            .in1(N__17006),
            .in2(N__16893),
            .in3(N__18893),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_96_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNICE00K_1_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNICE00K_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNICE00K_1_LC_8_9_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNICE00K_1_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__18374),
            .in2(N__16890),
            .in3(N__21343),
            .lcout(\Lab_UT.dictrl.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_3_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_3_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIQ1339_3_LC_8_9_6 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIQ1339_3_LC_8_9_6  (
            .in0(N__22092),
            .in1(N__16887),
            .in2(_gnd_net_),
            .in3(N__16880),
            .lcout(\Lab_UT.dictrl.N_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIFKL21_0_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIFKL21_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIFKL21_0_LC_8_10_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIFKL21_0_LC_8_10_0  (
            .in0(N__21724),
            .in1(N__17082),
            .in2(N__17111),
            .in3(N__18282),
            .lcout(\Lab_UT.dictrl.g1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIS94O2_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIS94O2_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIS94O2_LC_8_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIS94O2_LC_8_10_1  (
            .in0(N__18981),
            .in1(N__16854),
            .in2(N__17088),
            .in3(N__16827),
            .lcout(\Lab_UT.dictrl.N_119_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_8_10_3 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_8_10_3  (
            .in0(N__16806),
            .in1(N__16797),
            .in2(N__19554),
            .in3(N__21945),
            .lcout(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI0DI21_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI0DI21_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI0DI21_LC_8_10_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNI0DI21_LC_8_10_4  (
            .in0(N__17086),
            .in1(N__18281),
            .in2(N__21579),
            .in3(N__17391),
            .lcout(\Lab_UT.dictrl.g0_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_13_LC_8_10_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_13_LC_8_10_5  (
            .in0(N__18300),
            .in1(N__17104),
            .in2(N__17087),
            .in3(N__21723),
            .lcout(\Lab_UT.dictrl.g1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIEIOO8_0_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIEIOO8_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIEIOO8_0_LC_8_11_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIEIOO8_0_LC_8_11_0  (
            .in0(N__21949),
            .in1(N__16905),
            .in2(N__21975),
            .in3(N__16917),
            .lcout(\Lab_UT.dictrl.next_state_RNIEIOO8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIPHQ67_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIPHQ67_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIPHQ67_LC_8_11_1 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIPHQ67_LC_8_11_1  (
            .in0(N__17043),
            .in1(N__16923),
            .in2(N__21147),
            .in3(N__22056),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_1300_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOH1FC_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOH1FC_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOH1FC_LC_8_11_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOH1FC_LC_8_11_2  (
            .in0(N__16998),
            .in1(N__18889),
            .in2(N__16956),
            .in3(N__16953),
            .lcout(\Lab_UT.dictrl.N_96_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOJ371_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOJ371_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOJ371_LC_8_11_3 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIOJ371_LC_8_11_3  (
            .in0(N__21125),
            .in1(N__20855),
            .in2(N__21946),
            .in3(N__20652),
            .lcout(\Lab_UT.dictrl.g0_4_a4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_5_x1_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_5_x1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_5_x1_LC_8_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_5_x1_LC_8_12_0  (
            .in0(N__21432),
            .in1(N__17429),
            .in2(N__21648),
            .in3(N__21720),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_5_5_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_5_ns_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_5_ns_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_5_ns_LC_8_12_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.g0_5_5_ns_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16947),
            .in3(N__16941),
            .lcout(\Lab_UT.dictrl.g0_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIP5KF4_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIP5KF4_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIP5KF4_LC_8_12_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIP5KF4_LC_8_12_2  (
            .in0(N__21947),
            .in1(N__21145),
            .in2(N__19902),
            .in3(N__22040),
            .lcout(\Lab_UT.dictrl.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIN8JN3_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIN8JN3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIN8JN3_LC_8_12_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIN8JN3_LC_8_12_3  (
            .in0(N__19899),
            .in1(N__17121),
            .in2(N__18888),
            .in3(N__16911),
            .lcout(\Lab_UT.dictrl.N_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_3_RNI9ARR_LC_8_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_3_RNI9ARR_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_ret_3_RNI9ARR_LC_8_12_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \buart.Z_rx.shifter_ret_3_RNI9ARR_LC_8_12_6  (
            .in0(N__21628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21561),
            .lcout(N_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m33_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m33_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m33_LC_8_13_0 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \Lab_UT.dictrl.m33_LC_8_13_0  (
            .in0(N__17430),
            .in1(N__21721),
            .in2(N__19077),
            .in3(N__19044),
            .lcout(\Lab_UT.dictrl.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m30_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m30_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m30_LC_8_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m30_LC_8_13_1  (
            .in0(N__17194),
            .in1(N__17387),
            .in2(N__17276),
            .in3(N__17346),
            .lcout(\Lab_UT.dictrl.N_98_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_28_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_28_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_28_LC_8_13_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.g0_28_LC_8_13_2  (
            .in0(N__17313),
            .in1(N__17269),
            .in2(N__17244),
            .in3(N__17196),
            .lcout(\Lab_UT.dictrl.g1_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m31_ns_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m31_ns_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m31_ns_LC_8_13_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.m31_ns_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__17235),
            .in2(_gnd_net_),
            .in3(N__17202),
            .lcout(\Lab_UT.dictrl.N_84 ),
            .ltout(\Lab_UT.dictrl.N_84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_1_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_LC_8_13_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \Lab_UT.dictrl.g1_1_LC_8_13_5  (
            .in0(N__17195),
            .in1(N__17163),
            .in2(N__17154),
            .in3(N__20853),
            .lcout(\Lab_UT.dictrl.g1_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.shifter_ret_1_RNI1OGT_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.shifter_ret_1_RNI1OGT_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.shifter_ret_1_RNI1OGT_LC_8_14_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.shifter_ret_1_RNI1OGT_LC_8_14_1  (
            .in0(N__20702),
            .in1(N__17151),
            .in2(_gnd_net_),
            .in3(N__18191),
            .lcout(\Lab_UT.dictrl.m68_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIG3207_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIG3207_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIG3207_LC_8_14_2 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIG3207_LC_8_14_2  (
            .in0(N__19900),
            .in1(N__20703),
            .in2(N__17130),
            .in3(N__22020),
            .lcout(\Lab_UT.dictrl.N_95_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_4_a4_5_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_4_a4_5_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_4_a4_5_LC_8_14_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_4_a4_5_LC_8_14_3  (
            .in0(N__20984),
            .in1(N__21077),
            .in2(N__21580),
            .in3(N__21621),
            .lcout(\Lab_UT.dictrl.g0_4_a4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_9_1_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_9_1_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_9_1_0  (
            .in0(N__17461),
            .in1(N__17858),
            .in2(N__17958),
            .in3(N__17643),
            .lcout(\Lab_UT.didp.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22855),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_1_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI1S78_1_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(N__17460),
            .in2(_gnd_net_),
            .in3(N__17925),
            .lcout(\Lab_UT.didp.countrce2.un13_qPone ),
            .ltout(\Lab_UT.didp.countrce2.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_9_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_9_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_3_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17697),
            .in3(N__17510),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_1_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_1_3 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_9_1_3  (
            .in0(N__17895),
            .in1(N__18738),
            .in2(N__17694),
            .in3(N__17676),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_9_1_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_9_1_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_9_1_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_9_1_4  (
            .in0(N__17957),
            .in1(N__17677),
            .in2(N__17691),
            .in3(N__17859),
            .lcout(\Lab_UT.didp.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22855),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_9_2_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_9_2_0 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_0_LC_9_2_0  (
            .in0(N__17886),
            .in1(N__18231),
            .in2(_gnd_net_),
            .in3(N__17462),
            .lcout(\Lab_UT.didp.countrce2.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_9_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_9_2_1 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_9_2_1  (
            .in0(N__17637),
            .in1(N__17526),
            .in2(N__17517),
            .in3(N__17890),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_9_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_9_2_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_9_2_2  (
            .in0(N__17514),
            .in1(N__17948),
            .in2(N__17520),
            .in3(N__17852),
            .lcout(\Lab_UT.didp.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22852),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_9_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_9_2_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_1_LC_9_2_4  (
            .in0(N__20892),
            .in1(N__17463),
            .in2(N__17894),
            .in3(N__17926),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_9_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_9_2_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_9_2_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_9_2_5  (
            .in0(N__17927),
            .in1(N__17947),
            .in2(N__17931),
            .in3(N__17851),
            .lcout(\Lab_UT.didp.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22852),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_9_3_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_9_3_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_LC_9_3_0  (
            .in0(N__19702),
            .in1(N__19981),
            .in2(N__17748),
            .in3(N__19944),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22849),
            .ce(N__18252),
            .sr(N__22507));
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_3_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_3_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_9_3_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_LC_9_3_1  (
            .in0(N__19946),
            .in1(N__17746),
            .in2(N__19989),
            .in3(N__19704),
            .lcout(\Lab_UT.LdStens_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22849),
            .ce(N__18252),
            .sr(N__22507));
    defparam \Lab_UT.dictrl.state_ret_7_esr_LC_9_3_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_esr_LC_9_3_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_7_esr_LC_9_3_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_esr_LC_9_3_3  (
            .in0(N__19945),
            .in1(N__17745),
            .in2(N__19988),
            .in3(N__19703),
            .lcout(\Lab_UT.LdStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22849),
            .ce(N__18252),
            .sr(N__22507));
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_9_3_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI62AM_1_LC_9_3_4  (
            .in0(N__17871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17865),
            .lcout(\Lab_UT.didp.un1_dicLdStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_3_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_3_6 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_9_3_6  (
            .in0(N__18227),
            .in1(N__17815),
            .in2(_gnd_net_),
            .in3(N__17799),
            .lcout(\Lab_UT.didp.countrce1.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_ess_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_ess_LC_9_4_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_9_ess_LC_9_4_4 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_ess_LC_9_4_4  (
            .in0(N__19701),
            .in1(N__19973),
            .in2(N__17747),
            .in3(N__19943),
            .lcout(\Lab_UT.LdSones_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22841),
            .ce(N__18251),
            .sr(N__22506));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_5_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_9_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__19377),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_5_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__19147),
            .in2(_gnd_net_),
            .in3(N__18042),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_5_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__19186),
            .in2(_gnd_net_),
            .in3(N__18033),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_5_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__19799),
            .in2(_gnd_net_),
            .in3(N__18030),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_9_5_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_9_5_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_9_5_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_9_5_4  (
            .in0(N__19402),
            .in1(N__22981),
            .in2(N__19122),
            .in3(N__18027),
            .lcout(buart__rx_bitcount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22834),
            .ce(N__19350),
            .sr(N__22530));
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_9_6_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_9_6_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_LC_9_6_0  (
            .in0(N__17989),
            .in1(N__18401),
            .in2(_gnd_net_),
            .in3(N__20509),
            .lcout(\Lab_UT.dictrl.state_i_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__18250),
            .sr(N__22503));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_9_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_9_6_2  (
            .in0(N__17988),
            .in1(N__18363),
            .in2(_gnd_net_),
            .in3(N__20414),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_6_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_6_3 .LUT_INIT=16'b0010011100001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_LC_9_6_3  (
            .in0(N__17993),
            .in1(N__18378),
            .in2(N__18003),
            .in3(N__21299),
            .lcout(\Lab_UT.dictrl.state_i_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__18250),
            .sr(N__22503));
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_9_6_4 .LUT_INIT=16'b0011010100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_LC_9_6_4  (
            .in0(N__18402),
            .in1(N__20510),
            .in2(N__17994),
            .in3(N__19700),
            .lcout(\Lab_UT.dictrl.dicLdStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__18250),
            .sr(N__22503));
    defparam \Lab_UT.dictrl.state_0_esr_RNI9CU3Q_2_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI9CU3Q_2_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI9CU3Q_2_LC_9_7_0 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI9CU3Q_2_LC_9_7_0  (
            .in0(N__20413),
            .in1(N__18317),
            .in2(N__20177),
            .in3(N__21880),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI4L025_3_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4L025_3_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4L025_3_LC_9_7_1 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI4L025_3_LC_9_7_1  (
            .in0(N__22198),
            .in1(N__18609),
            .in2(N__20332),
            .in3(N__21294),
            .lcout(\Lab_UT.dictrl.N_101 ),
            .ltout(\Lab_UT.dictrl.N_101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI3QHJ5_1_LC_9_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI3QHJ5_1_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI3QHJ5_1_LC_9_7_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI3QHJ5_1_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__18333),
            .in2(N__18321),
            .in3(N__21879),
            .lcout(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_state_RNI3QHJ5Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_9_7_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_1_LC_9_7_3  (
            .in0(N__21885),
            .in1(N__18318),
            .in2(N__18303),
            .in3(N__20151),
            .lcout(\Lab_UT.dictrl.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22820),
            .ce(N__18248),
            .sr(N__22502));
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_9_7_4 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_3_LC_9_7_4  (
            .in0(N__19259),
            .in1(N__19291),
            .in2(N__20179),
            .in3(N__21886),
            .lcout(\Lab_UT.dictrl.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22820),
            .ce(N__18248),
            .sr(N__22502));
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_9_7_5 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_3_LC_9_7_5  (
            .in0(N__20159),
            .in1(N__19293),
            .in2(N__21936),
            .in3(N__19260),
            .lcout(\Lab_UT.dictrl.state_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22820),
            .ce(N__18248),
            .sr(N__22502));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_9_7_6 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_LC_9_7_6  (
            .in0(N__19257),
            .in1(N__19290),
            .in2(N__20178),
            .in3(N__21881),
            .lcout(\Lab_UT.dictrl.state_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22820),
            .ce(N__18248),
            .sr(N__22502));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_9_7_7 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_LC_9_7_7  (
            .in0(N__20158),
            .in1(N__19292),
            .in2(N__21935),
            .in3(N__19258),
            .lcout(\Lab_UT.dictrl.state_3_rep2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22820),
            .ce(N__18248),
            .sr(N__22502));
    defparam \Lab_UT.dictrl.g0_30_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_30_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_30_LC_9_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_30_LC_9_8_0  (
            .in0(N__18549),
            .in1(N__18216),
            .in2(N__18093),
            .in3(N__18081),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_116_mux_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIU2C38_3_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIU2C38_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIU2C38_3_LC_9_8_1 .LUT_INIT=16'b1110001011110011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIU2C38_3_LC_9_8_1  (
            .in0(N__20337),
            .in1(N__22202),
            .in2(N__18051),
            .in3(N__22104),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_120_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNI5OGCH_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNI5OGCH_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNI5OGCH_LC_9_8_2 .LUT_INIT=16'b1110111100000001;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNI5OGCH_LC_9_8_2  (
            .in0(N__21296),
            .in1(N__21931),
            .in2(N__18459),
            .in3(N__18420),
            .lcout(\Lab_UT.dictrl.N_1302_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIHNKSM_3_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIHNKSM_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIHNKSM_3_LC_9_8_3 .LUT_INIT=16'b0000110001010101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIHNKSM_3_LC_9_8_3  (
            .in0(N__18807),
            .in1(N__18585),
            .in2(N__20367),
            .in3(N__21297),
            .lcout(\Lab_UT.dictrl.N_119_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNIVIE9H_LC_9_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNIVIE9H_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNIVIE9H_LC_9_9_0 .LUT_INIT=16'b1100110011000101;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNIVIE9H_LC_9_9_0  (
            .in0(N__18387),
            .in1(N__18419),
            .in2(N__21950),
            .in3(N__21344),
            .lcout(\Lab_UT.dictrl.state_ret_12_RNIVIE9HZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIOT908_3_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIOT908_3_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIOT908_3_LC_9_9_1 .LUT_INIT=16'b1010110010101111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIOT908_3_LC_9_9_1  (
            .in0(N__20486),
            .in1(N__20336),
            .in2(N__22249),
            .in3(N__22105),
            .lcout(\Lab_UT.dictrl.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_3_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_3_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_3_LC_9_9_2 .LUT_INIT=16'b0001010100011111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI4CET7_3_LC_9_9_2  (
            .in0(N__22220),
            .in1(N__20485),
            .in2(N__20366),
            .in3(N__19024),
            .lcout(\Lab_UT.dictrl.N_99 ),
            .ltout(\Lab_UT.dictrl.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_1_LC_9_9_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_1_LC_9_9_3  (
            .in0(N__21345),
            .in1(N__18359),
            .in2(N__18348),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_9_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_1_LC_9_9_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__18345),
            .in2(N__18336),
            .in3(N__20168),
            .lcout(\Lab_UT.dictrl.next_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22805),
            .ce(N__22295),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIH7T88_3_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH7T88_3_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH7T88_3_LC_9_10_0 .LUT_INIT=16'b0000001100100010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIH7T88_3_LC_9_10_0  (
            .in0(N__22090),
            .in1(N__20305),
            .in2(N__19025),
            .in3(N__22219),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI51E3N_1_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI51E3N_1_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI51E3N_1_LC_9_10_1 .LUT_INIT=16'b1010000011110101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI51E3N_1_LC_9_10_1  (
            .in0(N__21342),
            .in1(_gnd_net_),
            .in2(N__18324),
            .in3(N__18750),
            .lcout(\Lab_UT.dictrl.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI48008_3_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI48008_3_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI48008_3_LC_9_10_2 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI48008_3_LC_9_10_2  (
            .in0(N__22089),
            .in1(N__20304),
            .in2(N__18899),
            .in3(N__18777),
            .lcout(\Lab_UT.dictrl.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI89VA1_3_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI89VA1_3_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI89VA1_3_LC_9_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI89VA1_3_LC_9_10_4  (
            .in0(N__20300),
            .in1(N__22216),
            .in2(N__21948),
            .in3(N__21340),
            .lcout(\Lab_UT.dictrl.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_0_3_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_0_3_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI4CET7_0_3_LC_9_10_5 .LUT_INIT=16'b0001010100011111;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI4CET7_0_3_LC_9_10_5  (
            .in0(N__22217),
            .in1(N__20481),
            .in2(N__20346),
            .in3(N__19016),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_99_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIJGPPK_1_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIJGPPK_1_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIJGPPK_1_LC_9_10_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIJGPPK_1_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__21341),
            .in2(N__18594),
            .in3(N__18591),
            .lcout(\Lab_UT.dictrl.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIOIJR7_0_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIOIJR7_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIOIJR7_0_LC_9_10_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIOIJR7_0_LC_9_10_7  (
            .in0(N__22218),
            .in1(N__19017),
            .in2(_gnd_net_),
            .in3(N__22088),
            .lcout(\Lab_UT.dictrl.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIPED74_3_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIPED74_3_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIPED74_3_LC_9_11_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIPED74_3_LC_9_11_0  (
            .in0(N__20341),
            .in1(N__18897),
            .in2(_gnd_net_),
            .in3(N__18776),
            .lcout(\Lab_UT.dictrl.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_1  (
            .in0(N__20970),
            .in1(N__21065),
            .in2(N__18900),
            .in3(N__21650),
            .lcout(\Lab_UT.dictrl.g0_0_0_a3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_37_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_37_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_37_LC_9_11_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.g0_37_LC_9_11_3  (
            .in0(N__20969),
            .in1(N__21064),
            .in2(N__21572),
            .in3(N__21649),
            .lcout(\Lab_UT.dictrl.N_98_mux_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_5_LC_9_11_4 .C_ON=1'b0;
    defparam \resetGen.escKey_5_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_5_LC_9_11_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \resetGen.escKey_5_LC_9_11_4  (
            .in0(N__21651),
            .in1(N__18548),
            .in2(N__20664),
            .in3(N__21556),
            .lcout(),
            .ltout(\resetGen.escKeyZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_9_11_5 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_9_11_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \resetGen.escKey_LC_9_11_5  (
            .in0(N__18498),
            .in1(N__19800),
            .in2(N__18486),
            .in3(N__19740),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKE4Q8_0_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKE4Q8_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKE4Q8_0_LC_9_12_0 .LUT_INIT=16'b0011101011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKE4Q8_0_LC_9_12_0  (
            .in0(N__22039),
            .in1(N__18887),
            .in2(N__22263),
            .in3(N__18921),
            .lcout(\Lab_UT.dictrl.g2_0_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIGU6P7_LC_9_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIGU6P7_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIGU6P7_LC_9_12_1 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIGU6P7_LC_9_12_1  (
            .in0(N__19894),
            .in1(N__18912),
            .in2(N__18898),
            .in3(N__22038),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_95_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI9TD6E_0_LC_9_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI9TD6E_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI9TD6E_0_LC_9_12_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI9TD6E_0_LC_9_12_2  (
            .in0(N__22247),
            .in1(_gnd_net_),
            .in2(N__18810),
            .in3(N__18959),
            .lcout(\Lab_UT.dictrl.N_103_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_2_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_2_LC_9_12_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \Lab_UT.dictrl.g1_2_LC_9_12_3  (
            .in0(N__20865),
            .in1(N__19080),
            .in2(N__18798),
            .in3(N__20660),
            .lcout(\Lab_UT.dictrl.g1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m47_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m47_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m47_LC_9_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.m47_LC_9_12_4  (
            .in0(N__19079),
            .in1(N__20864),
            .in2(_gnd_net_),
            .in3(N__19047),
            .lcout(\Lab_UT.dictrl.N_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIT67DE_0_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIT67DE_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIT67DE_0_LC_9_12_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIT67DE_0_LC_9_12_7  (
            .in0(N__18960),
            .in1(_gnd_net_),
            .in2(N__18762),
            .in3(N__22248),
            .lcout(\Lab_UT.dictrl.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m63_0_1_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m63_0_1_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m63_0_1_LC_9_13_0 .LUT_INIT=16'b0100011111001111;
    LogicCell40 \Lab_UT.dictrl.m63_0_1_LC_9_13_0  (
            .in0(N__19046),
            .in1(N__18714),
            .in2(N__19078),
            .in3(N__21728),
            .lcout(\Lab_UT.dictrl.m63_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIVHJND_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIVHJND_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIVHJND_0_LC_9_13_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIVHJND_0_LC_9_13_2  (
            .in0(N__22243),
            .in1(N__18933),
            .in2(_gnd_net_),
            .in3(N__18600),
            .lcout(\Lab_UT.dictrl.N_103_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m48_LC_9_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m48_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m48_LC_9_13_5 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \Lab_UT.dictrl.m48_LC_9_13_5  (
            .in0(N__20854),
            .in1(N__19068),
            .in2(N__20706),
            .in3(N__19045),
            .lcout(\Lab_UT.dictrl.N_89 ),
            .ltout(\Lab_UT.dictrl.N_89_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI3DTV5_LC_9_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI3DTV5_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI3DTV5_LC_9_13_6 .LUT_INIT=16'b0001101101011111;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNI3DTV5_LC_9_13_6  (
            .in0(N__19895),
            .in1(N__18990),
            .in2(N__18984),
            .in3(N__18980),
            .lcout(\Lab_UT.dictrl.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIPS7A6_LC_9_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIPS7A6_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIPS7A6_LC_9_14_2 .LUT_INIT=16'b0011101011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIPS7A6_LC_9_14_2  (
            .in0(N__18951),
            .in1(N__20704),
            .in2(N__19893),
            .in3(N__18939),
            .lcout(\Lab_UT.dictrl.N_102_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_11_3_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_11_3_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3HE3_5_LC_11_3_0  (
            .in0(N__23063),
            .in1(N__20545),
            .in2(N__22929),
            .in3(N__20581),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_11_3_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_11_3_1 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_4_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__23047),
            .in2(N__18927),
            .in3(N__20562),
            .lcout(buart__rx_ser_clk),
            .ltout(buart__rx_ser_clk_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_11_3_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_11_3_2 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_11_3_2  (
            .in0(N__23073),
            .in1(N__22983),
            .in2(N__18924),
            .in3(N__20546),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22853),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_11_3_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_11_3_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_11_3_3 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_11_3_3  (
            .in0(N__20582),
            .in1(_gnd_net_),
            .in2(N__22994),
            .in3(N__20564),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22853),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_11_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_11_3_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_11_3_4  (
            .in0(N__23048),
            .in1(N__23021),
            .in2(N__23034),
            .in3(N__22987),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22853),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_11_3_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_11_3_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_11_3_5  (
            .in0(N__22982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20563),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22853),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNICF9U4_3_LC_11_3_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNICF9U4_3_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNICF9U4_3_LC_11_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNICF9U4_3_LC_11_3_6  (
            .in0(N__22869),
            .in1(N__21897),
            .in2(_gnd_net_),
            .in3(N__19236),
            .lcout(\Lab_UT.dictrl.next_state_RNICF9U4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m91_LC_11_4_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m91_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m91_LC_11_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.m91_LC_11_4_0  (
            .in0(N__19371),
            .in1(N__19126),
            .in2(N__19167),
            .in3(N__19198),
            .lcout(\Lab_UT.dictrl.N_102_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m81_e_LC_11_4_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m81_e_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m81_e_LC_11_4_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dictrl.m81_e_LC_11_4_1  (
            .in0(N__19127),
            .in1(N__19165),
            .in2(_gnd_net_),
            .in3(N__19774),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m82_LC_11_4_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m82_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m82_LC_11_4_2 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \Lab_UT.dictrl.m82_LC_11_4_2  (
            .in0(N__19372),
            .in1(N__23016),
            .in2(N__19221),
            .in3(N__19199),
            .lcout(buart__rx_sample),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_11_4_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_11_4_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIFSPI1_4_LC_11_4_3  (
            .in0(N__19197),
            .in1(N__19161),
            .in2(N__19128),
            .in3(N__19370),
            .lcout(buart__rx_valid_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_11_5_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_11_5_0 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_11_5_0  (
            .in0(N__19098),
            .in1(N__23022),
            .in2(_gnd_net_),
            .in3(N__19509),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m89_bm_LC_11_5_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m89_bm_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m89_bm_LC_11_5_1 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \Lab_UT.dictrl.m89_bm_LC_11_5_1  (
            .in0(N__19417),
            .in1(N__19452),
            .in2(N__19503),
            .in3(N__19776),
            .lcout(m89_bm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.N_27_0_i_LC_11_5_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.N_27_0_i_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.N_27_0_i_LC_11_5_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Lab_UT.dictrl.N_27_0_i_LC_11_5_2  (
            .in0(N__19726),
            .in1(_gnd_net_),
            .in2(N__19789),
            .in3(N__19418),
            .lcout(buart__rx_N_27_0_i),
            .ltout(buart__rx_N_27_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_11_5_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_11_5_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_11_5_3 .LUT_INIT=16'b0011010100111010;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_11_5_3  (
            .in0(N__19092),
            .in1(N__22980),
            .in2(N__19083),
            .in3(N__19781),
            .lcout(buart__rx_bitcount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22842),
            .ce(N__19345),
            .sr(N__22532));
    defparam \Lab_UT.dictrl.m9_LC_11_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m9_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m9_LC_11_5_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.dictrl.m9_LC_11_5_4  (
            .in0(N__19451),
            .in1(N__19498),
            .in2(_gnd_net_),
            .in3(N__19416),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_107_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m89_am_LC_11_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m89_am_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m89_am_LC_11_5_5 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \Lab_UT.dictrl.m89_am_LC_11_5_5  (
            .in0(_gnd_net_),
            .in1(N__19775),
            .in2(N__19512),
            .in3(N__19725),
            .lcout(m89_am),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m10_LC_11_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m10_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m10_LC_11_5_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m10_LC_11_5_6  (
            .in0(N__19777),
            .in1(N__19502),
            .in2(N__19468),
            .in3(N__19419),
            .lcout(buart__rx_startbit),
            .ltout(buart__rx_startbit_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_11_5_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_11_5_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_11_5_7 .LUT_INIT=16'b0001110100101110;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_11_5_7  (
            .in0(N__22899),
            .in1(N__19401),
            .in2(N__19380),
            .in3(N__19376),
            .lcout(buart__rx_bitcount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22842),
            .ce(N__19345),
            .sr(N__22532));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_11_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_6_LC_11_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_6_LC_11_6_5  (
            .in0(N__19545),
            .in1(N__21837),
            .in2(_gnd_net_),
            .in3(N__19320),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_2000_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_11_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_2_LC_11_6_6 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_2_LC_11_6_6  (
            .in0(N__21838),
            .in1(N__19308),
            .in2(N__19296),
            .in3(N__20182),
            .lcout(\Lab_UT.dictrl.next_state_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_11_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_3_LC_11_7_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_3_LC_11_7_0  (
            .in0(N__22580),
            .in1(N__21835),
            .in2(_gnd_net_),
            .in3(N__19638),
            .lcout(\Lab_UT.dictrl.state_ret_12_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_11_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_1_LC_11_7_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_1_LC_11_7_2  (
            .in0(N__22582),
            .in1(N__19677),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\Lab_UT.dictrl.state_ret_12and_a0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKRG8A_2_LC_11_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKRG8A_2_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKRG8A_2_LC_11_7_3 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKRG8A_2_LC_11_7_3  (
            .in0(N__19279),
            .in1(N__19256),
            .in2(N__21903),
            .in3(N__20141),
            .lcout(Lab_UT_dictrl_next_state_3),
            .ltout(Lab_UT_dictrl_next_state_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_11_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_4_LC_11_7_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_4_LC_11_7_4  (
            .in0(N__22581),
            .in1(N__21836),
            .in2(N__20016),
            .in3(N__19639),
            .lcout(\Lab_UT.dictrl.state_ret_12_RNOZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_RNO_0_LC_11_7_6  (
            .in0(N__20013),
            .in1(N__20007),
            .in2(_gnd_net_),
            .in3(N__20001),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_12and_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_12_LC_11_7_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_12_LC_11_7_7  (
            .in0(N__19995),
            .in1(N__19972),
            .in2(N__19950),
            .in3(N__19942),
            .lcout(Lab_UT_dictrl_un1_next_state66_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22826),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIH05S_LC_11_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIH05S_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIH05S_LC_11_8_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIH05S_LC_11_8_1  (
            .in0(N__21367),
            .in1(N__19887),
            .in2(_gnd_net_),
            .in3(N__21820),
            .lcout(\Lab_UT.dictrl.m46_i_0_a5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m3_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m3_LC_11_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.m3_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__19788),
            .in2(_gnd_net_),
            .in3(N__19736),
            .lcout(bu_rx_data_rdy),
            .ltout(bu_rx_data_rdy_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_RNIMHUCC_LC_11_8_5 .C_ON=1'b0;
    defparam \resetGen.rst_RNIMHUCC_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.rst_RNIMHUCC_LC_11_8_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \resetGen.rst_RNIMHUCC_LC_11_8_5  (
            .in0(N__21839),
            .in1(N__19676),
            .in2(N__19650),
            .in3(N__19646),
            .lcout(\resetGen.r_m3_i_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_11_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_2_LC_11_9_0 .LUT_INIT=16'b1000010110000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_2_LC_11_9_0  (
            .in0(N__21369),
            .in1(N__20532),
            .in2(N__22264),
            .in3(N__19593),
            .lcout(),
            .ltout(\Lab_UT.dictrl.i9_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_2_LC_11_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_2_LC_11_9_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__20183),
            .in2(N__19575),
            .in3(N__19571),
            .lcout(\Lab_UT.dictrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22815),
            .ce(N__22282),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_11_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_11_9_2 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_0_LC_11_9_2  (
            .in0(N__22252),
            .in1(N__20531),
            .in2(N__20373),
            .in3(N__22107),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_11_9_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_0_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__21370),
            .in2(N__20517),
            .in3(N__20439),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_0_LC_11_9_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_11_9_4  (
            .in0(N__20184),
            .in1(N__20514),
            .in2(N__20490),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.next_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22815),
            .ce(N__22282),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_11_9_5 .LUT_INIT=16'b0000001011001110;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_0_LC_11_9_5  (
            .in0(N__22106),
            .in1(N__22251),
            .in2(N__20372),
            .in3(N__20487),
            .lcout(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIL2ATH_0_LC_11_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIL2ATH_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIL2ATH_0_LC_11_10_0 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIL2ATH_0_LC_11_10_0  (
            .in0(N__21735),
            .in1(N__21981),
            .in2(N__20433),
            .in3(N__22097),
            .lcout(\Lab_UT.dictrl.N_1302_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIGENTQ_2_LC_11_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIGENTQ_2_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIGENTQ_2_LC_11_10_3 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIGENTQ_2_LC_11_10_3  (
            .in0(N__20418),
            .in1(N__20180),
            .in2(N__21942),
            .in3(N__20394),
            .lcout(N_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI38BCN_3_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI38BCN_3_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI38BCN_3_LC_11_10_6 .LUT_INIT=16'b0000100000111011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI38BCN_3_LC_11_10_6  (
            .in0(N__20385),
            .in1(N__21368),
            .in2(N__20369),
            .in3(N__20205),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_119_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIIE1Q91_2_LC_11_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIE1Q91_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIE1Q91_2_LC_11_10_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIIE1Q91_2_LC_11_10_7  (
            .in0(N__21899),
            .in1(N__20193),
            .in2(N__20187),
            .in3(N__20181),
            .lcout(Lab_UT_dictrl_next_state_0_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_4_LC_11_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_4_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_4_LC_11_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g1_4_LC_11_11_0  (
            .in0(N__21652),
            .in1(N__20980),
            .in2(N__21581),
            .in3(N__21441),
            .lcout(\Lab_UT.dictrl.g1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI6KC68_0_LC_11_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI6KC68_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI6KC68_0_LC_11_11_2 .LUT_INIT=16'b1100000011100000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI6KC68_0_LC_11_11_2  (
            .in0(N__22250),
            .in1(N__20991),
            .in2(N__22119),
            .in3(N__22103),
            .lcout(\Lab_UT.dictrl.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNISBBJ4_0_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNISBBJ4_0_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNISBBJ4_0_LC_11_11_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNISBBJ4_0_LC_11_11_3  (
            .in0(N__21968),
            .in1(N__21898),
            .in2(_gnd_net_),
            .in3(N__21183),
            .lcout(\Lab_UT.dictrl.m46_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_5_RNIIJHP1_LC_11_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_5_RNIIJHP1_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_ret_5_RNIIJHP1_LC_11_12_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \buart.Z_rx.shifter_ret_5_RNIIJHP1_LC_11_12_0  (
            .in0(N__21729),
            .in1(N__21657),
            .in2(N__21582),
            .in3(N__21440),
            .lcout(),
            .ltout(g0_3_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU7Q14_LC_11_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU7Q14_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU7Q14_LC_11_12_1 .LUT_INIT=16'b0010001000100000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIU7Q14_LC_11_12_1  (
            .in0(N__21167),
            .in1(N__21384),
            .in2(N__21198),
            .in3(N__21195),
            .lcout(\Lab_UT.dictrl.g1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIK8B43_LC_11_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIK8B43_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIK8B43_LC_11_12_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIK8B43_LC_11_12_7  (
            .in0(N__20589),
            .in1(N__21177),
            .in2(N__21168),
            .in3(N__21081),
            .lcout(\Lab_UT.dictrl.N_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_ret_6_rep1_RNI4S9J1_LC_11_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_ret_6_rep1_RNI4S9J1_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_ret_6_rep1_RNI4S9J1_LC_11_13_2 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \buart.Z_rx.shifter_ret_6_rep1_RNI4S9J1_LC_11_13_2  (
            .in0(N__20985),
            .in1(N__20852),
            .in2(N__20705),
            .in3(N__20651),
            .lcout(m46_i_0_a3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_12_3_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_12_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(N__20583),
            .in2(N__20568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_3_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_12_3_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_12_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(N__20547),
            .in2(_gnd_net_),
            .in3(N__23067),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_12_3_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_12_3_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_12_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_12_3_2  (
            .in0(N__22990),
            .in1(N__23064),
            .in2(_gnd_net_),
            .in3(N__23052),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__22856),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_12_3_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_12_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_12_3_3  (
            .in0(_gnd_net_),
            .in1(N__23049),
            .in2(_gnd_net_),
            .in3(N__23025),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_12_3_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_12_3_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_12_3_4 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_12_3_4  (
            .in0(N__22928),
            .in1(N__23020),
            .in2(N__22995),
            .in3(N__22932),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22856),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_12_5_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_12_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_3_LC_12_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22900),
            .lcout(\Lab_UT.dictrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22850),
            .ce(N__22299),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_ctle_LC_12_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_ctle_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_ctle_LC_12_8_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_ctle_LC_12_8_6  (
            .in0(_gnd_net_),
            .in1(N__22583),
            .in2(_gnd_net_),
            .in3(N__22558),
            .lcout(bu_rx_data_rdy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_RNIAL6V33_LC_12_9_2 .C_ON=1'b0;
    defparam \resetGen.rst_RNIAL6V33_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.rst_RNIAL6V33_LC_12_9_2 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \resetGen.rst_RNIAL6V33_LC_12_9_2  (
            .in0(N__22332),
            .in1(N__22326),
            .in2(N__22320),
            .in3(N__22305),
            .lcout(rst_RNIAL6V33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
