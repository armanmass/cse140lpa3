// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 21 2019 00:07:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__22396;
    wire N__22395;
    wire N__22394;
    wire N__22387;
    wire N__22386;
    wire N__22385;
    wire N__22378;
    wire N__22377;
    wire N__22376;
    wire N__22369;
    wire N__22368;
    wire N__22367;
    wire N__22360;
    wire N__22359;
    wire N__22358;
    wire N__22351;
    wire N__22350;
    wire N__22349;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22324;
    wire N__22323;
    wire N__22322;
    wire N__22315;
    wire N__22314;
    wire N__22313;
    wire N__22296;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22281;
    wire N__22278;
    wire N__22275;
    wire N__22274;
    wire N__22273;
    wire N__22272;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22268;
    wire N__22267;
    wire N__22266;
    wire N__22265;
    wire N__22264;
    wire N__22263;
    wire N__22262;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22251;
    wire N__22250;
    wire N__22249;
    wire N__22248;
    wire N__22247;
    wire N__22246;
    wire N__22245;
    wire N__22244;
    wire N__22243;
    wire N__22242;
    wire N__22241;
    wire N__22240;
    wire N__22239;
    wire N__22238;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22230;
    wire N__22229;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22215;
    wire N__22214;
    wire N__22213;
    wire N__22212;
    wire N__22211;
    wire N__22210;
    wire N__22209;
    wire N__22208;
    wire N__22207;
    wire N__22206;
    wire N__22205;
    wire N__22204;
    wire N__22203;
    wire N__22202;
    wire N__22201;
    wire N__22200;
    wire N__22199;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22185;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21998;
    wire N__21993;
    wire N__21990;
    wire N__21987;
    wire N__21986;
    wire N__21981;
    wire N__21978;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21963;
    wire N__21962;
    wire N__21957;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21949;
    wire N__21944;
    wire N__21939;
    wire N__21938;
    wire N__21937;
    wire N__21934;
    wire N__21933;
    wire N__21928;
    wire N__21923;
    wire N__21918;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21887;
    wire N__21884;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21869;
    wire N__21868;
    wire N__21865;
    wire N__21860;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21839;
    wire N__21838;
    wire N__21837;
    wire N__21836;
    wire N__21833;
    wire N__21830;
    wire N__21825;
    wire N__21822;
    wire N__21819;
    wire N__21814;
    wire N__21807;
    wire N__21806;
    wire N__21805;
    wire N__21804;
    wire N__21803;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21789;
    wire N__21788;
    wire N__21787;
    wire N__21786;
    wire N__21785;
    wire N__21782;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21768;
    wire N__21767;
    wire N__21766;
    wire N__21765;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21748;
    wire N__21735;
    wire N__21730;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21708;
    wire N__21705;
    wire N__21700;
    wire N__21693;
    wire N__21692;
    wire N__21689;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21678;
    wire N__21677;
    wire N__21676;
    wire N__21675;
    wire N__21674;
    wire N__21673;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21655;
    wire N__21650;
    wire N__21641;
    wire N__21638;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21581;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21565;
    wire N__21558;
    wire N__21557;
    wire N__21556;
    wire N__21555;
    wire N__21552;
    wire N__21545;
    wire N__21540;
    wire N__21539;
    wire N__21538;
    wire N__21535;
    wire N__21530;
    wire N__21525;
    wire N__21522;
    wire N__21521;
    wire N__21520;
    wire N__21519;
    wire N__21518;
    wire N__21513;
    wire N__21506;
    wire N__21501;
    wire N__21498;
    wire N__21495;
    wire N__21494;
    wire N__21493;
    wire N__21492;
    wire N__21487;
    wire N__21486;
    wire N__21483;
    wire N__21482;
    wire N__21481;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21449;
    wire N__21446;
    wire N__21439;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21424;
    wire N__21419;
    wire N__21410;
    wire N__21407;
    wire N__21396;
    wire N__21395;
    wire N__21392;
    wire N__21391;
    wire N__21390;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21379;
    wire N__21378;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21353;
    wire N__21352;
    wire N__21349;
    wire N__21340;
    wire N__21337;
    wire N__21336;
    wire N__21335;
    wire N__21330;
    wire N__21327;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21315;
    wire N__21314;
    wire N__21313;
    wire N__21312;
    wire N__21309;
    wire N__21308;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21292;
    wire N__21287;
    wire N__21282;
    wire N__21279;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21263;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21237;
    wire N__21236;
    wire N__21235;
    wire N__21234;
    wire N__21233;
    wire N__21232;
    wire N__21231;
    wire N__21230;
    wire N__21229;
    wire N__21224;
    wire N__21223;
    wire N__21218;
    wire N__21215;
    wire N__21214;
    wire N__21213;
    wire N__21212;
    wire N__21207;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21181;
    wire N__21176;
    wire N__21165;
    wire N__21162;
    wire N__21153;
    wire N__21152;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21140;
    wire N__21137;
    wire N__21136;
    wire N__21135;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21122;
    wire N__21121;
    wire N__21118;
    wire N__21117;
    wire N__21116;
    wire N__21115;
    wire N__21108;
    wire N__21105;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21095;
    wire N__21094;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21044;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21025;
    wire N__21022;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20988;
    wire N__20985;
    wire N__20980;
    wire N__20971;
    wire N__20958;
    wire N__20957;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20946;
    wire N__20945;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20909;
    wire N__20908;
    wire N__20905;
    wire N__20904;
    wire N__20901;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20875;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20861;
    wire N__20858;
    wire N__20849;
    wire N__20848;
    wire N__20847;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20828;
    wire N__20823;
    wire N__20816;
    wire N__20811;
    wire N__20796;
    wire N__20795;
    wire N__20794;
    wire N__20793;
    wire N__20792;
    wire N__20791;
    wire N__20790;
    wire N__20789;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20762;
    wire N__20761;
    wire N__20758;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20748;
    wire N__20747;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20723;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20711;
    wire N__20708;
    wire N__20703;
    wire N__20700;
    wire N__20699;
    wire N__20698;
    wire N__20697;
    wire N__20696;
    wire N__20695;
    wire N__20694;
    wire N__20693;
    wire N__20692;
    wire N__20691;
    wire N__20690;
    wire N__20689;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20684;
    wire N__20683;
    wire N__20682;
    wire N__20681;
    wire N__20680;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20669;
    wire N__20668;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20660;
    wire N__20659;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20627;
    wire N__20626;
    wire N__20625;
    wire N__20624;
    wire N__20623;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20618;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20453;
    wire N__20452;
    wire N__20451;
    wire N__20446;
    wire N__20439;
    wire N__20438;
    wire N__20433;
    wire N__20428;
    wire N__20425;
    wire N__20424;
    wire N__20423;
    wire N__20422;
    wire N__20421;
    wire N__20420;
    wire N__20419;
    wire N__20418;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20376;
    wire N__20373;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20354;
    wire N__20351;
    wire N__20348;
    wire N__20343;
    wire N__20342;
    wire N__20341;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20333;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20318;
    wire N__20313;
    wire N__20306;
    wire N__20301;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20291;
    wire N__20282;
    wire N__20279;
    wire N__20278;
    wire N__20277;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20204;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20196;
    wire N__20193;
    wire N__20192;
    wire N__20189;
    wire N__20184;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20157;
    wire N__20156;
    wire N__20153;
    wire N__20152;
    wire N__20149;
    wire N__20144;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20136;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20128;
    wire N__20127;
    wire N__20126;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20099;
    wire N__20096;
    wire N__20095;
    wire N__20094;
    wire N__20079;
    wire N__20076;
    wire N__20071;
    wire N__20068;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20051;
    wire N__20050;
    wire N__20047;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20031;
    wire N__20030;
    wire N__20027;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20007;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19991;
    wire N__19990;
    wire N__19989;
    wire N__19986;
    wire N__19985;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19928;
    wire N__19927;
    wire N__19924;
    wire N__19923;
    wire N__19922;
    wire N__19921;
    wire N__19920;
    wire N__19919;
    wire N__19918;
    wire N__19917;
    wire N__19916;
    wire N__19911;
    wire N__19910;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19886;
    wire N__19885;
    wire N__19884;
    wire N__19883;
    wire N__19882;
    wire N__19877;
    wire N__19874;
    wire N__19869;
    wire N__19866;
    wire N__19865;
    wire N__19864;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19850;
    wire N__19845;
    wire N__19842;
    wire N__19837;
    wire N__19832;
    wire N__19831;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19779;
    wire N__19778;
    wire N__19777;
    wire N__19776;
    wire N__19775;
    wire N__19774;
    wire N__19773;
    wire N__19770;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19740;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19712;
    wire N__19709;
    wire N__19698;
    wire N__19697;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19691;
    wire N__19688;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19675;
    wire N__19672;
    wire N__19669;
    wire N__19668;
    wire N__19663;
    wire N__19660;
    wire N__19653;
    wire N__19650;
    wire N__19641;
    wire N__19640;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19628;
    wire N__19627;
    wire N__19626;
    wire N__19623;
    wire N__19622;
    wire N__19619;
    wire N__19618;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19607;
    wire N__19606;
    wire N__19605;
    wire N__19602;
    wire N__19601;
    wire N__19600;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19590;
    wire N__19585;
    wire N__19582;
    wire N__19581;
    wire N__19578;
    wire N__19575;
    wire N__19570;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19549;
    wire N__19542;
    wire N__19539;
    wire N__19528;
    wire N__19515;
    wire N__19512;
    wire N__19511;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19507;
    wire N__19506;
    wire N__19503;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19497;
    wire N__19496;
    wire N__19491;
    wire N__19488;
    wire N__19485;
    wire N__19482;
    wire N__19479;
    wire N__19472;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19461;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19445;
    wire N__19442;
    wire N__19435;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19393;
    wire N__19392;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19359;
    wire N__19352;
    wire N__19349;
    wire N__19348;
    wire N__19347;
    wire N__19346;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19338;
    wire N__19333;
    wire N__19330;
    wire N__19327;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19305;
    wire N__19304;
    wire N__19301;
    wire N__19298;
    wire N__19293;
    wire N__19292;
    wire N__19291;
    wire N__19290;
    wire N__19289;
    wire N__19288;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19282;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19265;
    wire N__19258;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19254;
    wire N__19253;
    wire N__19252;
    wire N__19249;
    wire N__19248;
    wire N__19247;
    wire N__19242;
    wire N__19235;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19224;
    wire N__19217;
    wire N__19214;
    wire N__19211;
    wire N__19206;
    wire N__19201;
    wire N__19198;
    wire N__19191;
    wire N__19184;
    wire N__19167;
    wire N__19164;
    wire N__19163;
    wire N__19160;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19148;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19136;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19107;
    wire N__19104;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19094;
    wire N__19091;
    wire N__19088;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19062;
    wire N__19059;
    wire N__19056;
    wire N__19055;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19040;
    wire N__19037;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19024;
    wire N__19019;
    wire N__19016;
    wire N__19011;
    wire N__19008;
    wire N__18999;
    wire N__18998;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18986;
    wire N__18983;
    wire N__18982;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18970;
    wire N__18963;
    wire N__18962;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18950;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18931;
    wire N__18930;
    wire N__18925;
    wire N__18920;
    wire N__18915;
    wire N__18914;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18906;
    wire N__18905;
    wire N__18904;
    wire N__18903;
    wire N__18902;
    wire N__18901;
    wire N__18898;
    wire N__18891;
    wire N__18888;
    wire N__18887;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18872;
    wire N__18869;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18846;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18824;
    wire N__18823;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18807;
    wire N__18804;
    wire N__18803;
    wire N__18800;
    wire N__18799;
    wire N__18794;
    wire N__18791;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18779;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18749;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18704;
    wire N__18701;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18671;
    wire N__18670;
    wire N__18667;
    wire N__18662;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18630;
    wire N__18629;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18612;
    wire N__18611;
    wire N__18608;
    wire N__18607;
    wire N__18604;
    wire N__18603;
    wire N__18602;
    wire N__18593;
    wire N__18592;
    wire N__18591;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18568;
    wire N__18561;
    wire N__18558;
    wire N__18557;
    wire N__18554;
    wire N__18551;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18538;
    wire N__18535;
    wire N__18530;
    wire N__18527;
    wire N__18524;
    wire N__18519;
    wire N__18516;
    wire N__18515;
    wire N__18514;
    wire N__18511;
    wire N__18508;
    wire N__18507;
    wire N__18504;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18488;
    wire N__18483;
    wire N__18480;
    wire N__18479;
    wire N__18478;
    wire N__18477;
    wire N__18474;
    wire N__18473;
    wire N__18470;
    wire N__18469;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18445;
    wire N__18442;
    wire N__18441;
    wire N__18438;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18423;
    wire N__18422;
    wire N__18421;
    wire N__18420;
    wire N__18419;
    wire N__18418;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18396;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18348;
    wire N__18347;
    wire N__18346;
    wire N__18345;
    wire N__18342;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18338;
    wire N__18337;
    wire N__18336;
    wire N__18335;
    wire N__18334;
    wire N__18331;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18311;
    wire N__18302;
    wire N__18301;
    wire N__18300;
    wire N__18299;
    wire N__18298;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18278;
    wire N__18275;
    wire N__18270;
    wire N__18263;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18228;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18222;
    wire N__18221;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18207;
    wire N__18206;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18189;
    wire N__18184;
    wire N__18181;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18167;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18145;
    wire N__18140;
    wire N__18123;
    wire N__18122;
    wire N__18121;
    wire N__18120;
    wire N__18119;
    wire N__18118;
    wire N__18117;
    wire N__18116;
    wire N__18115;
    wire N__18114;
    wire N__18113;
    wire N__18112;
    wire N__18107;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18093;
    wire N__18092;
    wire N__18087;
    wire N__18082;
    wire N__18081;
    wire N__18080;
    wire N__18079;
    wire N__18078;
    wire N__18077;
    wire N__18074;
    wire N__18069;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18053;
    wire N__18048;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18028;
    wire N__18025;
    wire N__18012;
    wire N__18009;
    wire N__18008;
    wire N__18007;
    wire N__18004;
    wire N__18003;
    wire N__18002;
    wire N__17999;
    wire N__17998;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17986;
    wire N__17983;
    wire N__17982;
    wire N__17981;
    wire N__17980;
    wire N__17977;
    wire N__17976;
    wire N__17975;
    wire N__17972;
    wire N__17963;
    wire N__17958;
    wire N__17955;
    wire N__17950;
    wire N__17947;
    wire N__17940;
    wire N__17935;
    wire N__17928;
    wire N__17925;
    wire N__17922;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17909;
    wire N__17908;
    wire N__17907;
    wire N__17902;
    wire N__17897;
    wire N__17892;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17883;
    wire N__17882;
    wire N__17881;
    wire N__17878;
    wire N__17877;
    wire N__17870;
    wire N__17867;
    wire N__17866;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17845;
    wire N__17832;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17802;
    wire N__17801;
    wire N__17800;
    wire N__17799;
    wire N__17798;
    wire N__17797;
    wire N__17796;
    wire N__17795;
    wire N__17794;
    wire N__17793;
    wire N__17792;
    wire N__17791;
    wire N__17790;
    wire N__17787;
    wire N__17786;
    wire N__17775;
    wire N__17774;
    wire N__17773;
    wire N__17766;
    wire N__17757;
    wire N__17752;
    wire N__17749;
    wire N__17746;
    wire N__17743;
    wire N__17740;
    wire N__17733;
    wire N__17724;
    wire N__17721;
    wire N__17720;
    wire N__17719;
    wire N__17718;
    wire N__17713;
    wire N__17712;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17704;
    wire N__17701;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17679;
    wire N__17678;
    wire N__17677;
    wire N__17676;
    wire N__17675;
    wire N__17674;
    wire N__17671;
    wire N__17666;
    wire N__17663;
    wire N__17658;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17611;
    wire N__17610;
    wire N__17609;
    wire N__17604;
    wire N__17603;
    wire N__17600;
    wire N__17595;
    wire N__17592;
    wire N__17587;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17547;
    wire N__17546;
    wire N__17543;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17513;
    wire N__17512;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17493;
    wire N__17492;
    wire N__17491;
    wire N__17488;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17480;
    wire N__17477;
    wire N__17472;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17438;
    wire N__17433;
    wire N__17430;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17403;
    wire N__17400;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17359;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17334;
    wire N__17331;
    wire N__17330;
    wire N__17329;
    wire N__17328;
    wire N__17325;
    wire N__17318;
    wire N__17317;
    wire N__17316;
    wire N__17311;
    wire N__17306;
    wire N__17301;
    wire N__17300;
    wire N__17299;
    wire N__17298;
    wire N__17295;
    wire N__17294;
    wire N__17293;
    wire N__17292;
    wire N__17289;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17273;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17253;
    wire N__17252;
    wire N__17249;
    wire N__17248;
    wire N__17247;
    wire N__17244;
    wire N__17243;
    wire N__17240;
    wire N__17239;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17208;
    wire N__17205;
    wire N__17192;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17168;
    wire N__17165;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17145;
    wire N__17142;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17124;
    wire N__17123;
    wire N__17122;
    wire N__17119;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17103;
    wire N__17102;
    wire N__17101;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17087;
    wire N__17084;
    wire N__17083;
    wire N__17078;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17040;
    wire N__17037;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17008;
    wire N__17005;
    wire N__16998;
    wire N__16989;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16980;
    wire N__16979;
    wire N__16978;
    wire N__16975;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16947;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16920;
    wire N__16919;
    wire N__16914;
    wire N__16913;
    wire N__16912;
    wire N__16911;
    wire N__16910;
    wire N__16909;
    wire N__16906;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16884;
    wire N__16883;
    wire N__16882;
    wire N__16881;
    wire N__16880;
    wire N__16879;
    wire N__16878;
    wire N__16875;
    wire N__16868;
    wire N__16865;
    wire N__16860;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16838;
    wire N__16835;
    wire N__16832;
    wire N__16831;
    wire N__16830;
    wire N__16825;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16809;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16748;
    wire N__16747;
    wire N__16744;
    wire N__16743;
    wire N__16742;
    wire N__16741;
    wire N__16738;
    wire N__16735;
    wire N__16732;
    wire N__16725;
    wire N__16720;
    wire N__16717;
    wire N__16710;
    wire N__16707;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16698;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16634;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16624;
    wire N__16623;
    wire N__16618;
    wire N__16617;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16603;
    wire N__16602;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16556;
    wire N__16555;
    wire N__16554;
    wire N__16545;
    wire N__16544;
    wire N__16543;
    wire N__16542;
    wire N__16541;
    wire N__16540;
    wire N__16537;
    wire N__16530;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16481;
    wire N__16476;
    wire N__16475;
    wire N__16474;
    wire N__16473;
    wire N__16472;
    wire N__16471;
    wire N__16468;
    wire N__16457;
    wire N__16452;
    wire N__16451;
    wire N__16448;
    wire N__16447;
    wire N__16446;
    wire N__16445;
    wire N__16440;
    wire N__16437;
    wire N__16436;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16415;
    wire N__16410;
    wire N__16407;
    wire N__16406;
    wire N__16405;
    wire N__16404;
    wire N__16403;
    wire N__16400;
    wire N__16393;
    wire N__16390;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16370;
    wire N__16367;
    wire N__16364;
    wire N__16361;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16349;
    wire N__16348;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16330;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16314;
    wire N__16313;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16291;
    wire N__16290;
    wire N__16289;
    wire N__16284;
    wire N__16281;
    wire N__16276;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16259;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16238;
    wire N__16235;
    wire N__16234;
    wire N__16233;
    wire N__16232;
    wire N__16231;
    wire N__16228;
    wire N__16227;
    wire N__16224;
    wire N__16217;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16197;
    wire N__16194;
    wire N__16193;
    wire N__16192;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16181;
    wire N__16178;
    wire N__16171;
    wire N__16168;
    wire N__16161;
    wire N__16160;
    wire N__16155;
    wire N__16154;
    wire N__16153;
    wire N__16150;
    wire N__16145;
    wire N__16140;
    wire N__16139;
    wire N__16136;
    wire N__16135;
    wire N__16134;
    wire N__16125;
    wire N__16122;
    wire N__16121;
    wire N__16120;
    wire N__16117;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16099;
    wire N__16098;
    wire N__16095;
    wire N__16090;
    wire N__16085;
    wire N__16082;
    wire N__16077;
    wire N__16072;
    wire N__16069;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16040;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16025;
    wire N__16022;
    wire N__16017;
    wire N__16016;
    wire N__16013;
    wire N__16012;
    wire N__16005;
    wire N__16002;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15990;
    wire N__15987;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15975;
    wire N__15974;
    wire N__15973;
    wire N__15970;
    wire N__15965;
    wire N__15960;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15930;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15918;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15899;
    wire N__15896;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15882;
    wire N__15881;
    wire N__15880;
    wire N__15879;
    wire N__15878;
    wire N__15877;
    wire N__15876;
    wire N__15873;
    wire N__15868;
    wire N__15867;
    wire N__15866;
    wire N__15863;
    wire N__15856;
    wire N__15853;
    wire N__15850;
    wire N__15845;
    wire N__15842;
    wire N__15831;
    wire N__15828;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15816;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15806;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15773;
    wire N__15770;
    wire N__15767;
    wire N__15764;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15750;
    wire N__15747;
    wire N__15746;
    wire N__15745;
    wire N__15744;
    wire N__15743;
    wire N__15742;
    wire N__15741;
    wire N__15740;
    wire N__15739;
    wire N__15738;
    wire N__15737;
    wire N__15736;
    wire N__15731;
    wire N__15728;
    wire N__15719;
    wire N__15716;
    wire N__15711;
    wire N__15706;
    wire N__15699;
    wire N__15696;
    wire N__15691;
    wire N__15688;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15668;
    wire N__15667;
    wire N__15666;
    wire N__15665;
    wire N__15662;
    wire N__15657;
    wire N__15652;
    wire N__15645;
    wire N__15644;
    wire N__15643;
    wire N__15642;
    wire N__15641;
    wire N__15638;
    wire N__15635;
    wire N__15630;
    wire N__15625;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15611;
    wire N__15610;
    wire N__15609;
    wire N__15604;
    wire N__15603;
    wire N__15602;
    wire N__15601;
    wire N__15600;
    wire N__15597;
    wire N__15596;
    wire N__15593;
    wire N__15590;
    wire N__15589;
    wire N__15588;
    wire N__15587;
    wire N__15584;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15549;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15521;
    wire N__15520;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15508;
    wire N__15505;
    wire N__15498;
    wire N__15495;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15486;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15459;
    wire N__15458;
    wire N__15457;
    wire N__15456;
    wire N__15451;
    wire N__15446;
    wire N__15441;
    wire N__15440;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15398;
    wire N__15395;
    wire N__15388;
    wire N__15385;
    wire N__15378;
    wire N__15377;
    wire N__15376;
    wire N__15371;
    wire N__15368;
    wire N__15367;
    wire N__15364;
    wire N__15359;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15341;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15309;
    wire N__15308;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15281;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15263;
    wire N__15262;
    wire N__15259;
    wire N__15258;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15224;
    wire N__15221;
    wire N__15220;
    wire N__15217;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15195;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15164;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15113;
    wire N__15112;
    wire N__15111;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15074;
    wire N__15073;
    wire N__15072;
    wire N__15071;
    wire N__15070;
    wire N__15069;
    wire N__15064;
    wire N__15063;
    wire N__15060;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15036;
    wire N__15033;
    wire N__15032;
    wire N__15031;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15027;
    wire N__15024;
    wire N__15015;
    wire N__15010;
    wire N__15007;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14997;
    wire N__14996;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14980;
    wire N__14979;
    wire N__14978;
    wire N__14975;
    wire N__14974;
    wire N__14971;
    wire N__14968;
    wire N__14963;
    wire N__14962;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14937;
    wire N__14934;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14915;
    wire N__14914;
    wire N__14911;
    wire N__14910;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14885;
    wire N__14882;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14870;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14843;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14826;
    wire N__14823;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14724;
    wire N__14721;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14694;
    wire N__14691;
    wire N__14690;
    wire N__14685;
    wire N__14682;
    wire N__14681;
    wire N__14680;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14664;
    wire N__14661;
    wire N__14660;
    wire N__14659;
    wire N__14658;
    wire N__14657;
    wire N__14656;
    wire N__14655;
    wire N__14652;
    wire N__14639;
    wire N__14636;
    wire N__14633;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14612;
    wire N__14609;
    wire N__14604;
    wire N__14603;
    wire N__14602;
    wire N__14595;
    wire N__14592;
    wire N__14591;
    wire N__14588;
    wire N__14585;
    wire N__14580;
    wire N__14579;
    wire N__14576;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14534;
    wire N__14533;
    wire N__14528;
    wire N__14525;
    wire N__14520;
    wire N__14519;
    wire N__14516;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14493;
    wire N__14492;
    wire N__14491;
    wire N__14490;
    wire N__14487;
    wire N__14486;
    wire N__14483;
    wire N__14482;
    wire N__14479;
    wire N__14478;
    wire N__14475;
    wire N__14462;
    wire N__14457;
    wire N__14454;
    wire N__14453;
    wire N__14452;
    wire N__14451;
    wire N__14450;
    wire N__14443;
    wire N__14440;
    wire N__14439;
    wire N__14436;
    wire N__14431;
    wire N__14426;
    wire N__14421;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14410;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14391;
    wire N__14390;
    wire N__14389;
    wire N__14388;
    wire N__14387;
    wire N__14386;
    wire N__14373;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14361;
    wire N__14360;
    wire N__14357;
    wire N__14356;
    wire N__14355;
    wire N__14352;
    wire N__14351;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14317;
    wire N__14314;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14294;
    wire N__14293;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14262;
    wire N__14259;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14251;
    wire N__14246;
    wire N__14243;
    wire N__14242;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14224;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14210;
    wire N__14209;
    wire N__14208;
    wire N__14205;
    wire N__14202;
    wire N__14199;
    wire N__14196;
    wire N__14187;
    wire N__14186;
    wire N__14185;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14160;
    wire N__14159;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14151;
    wire N__14150;
    wire N__14149;
    wire N__14140;
    wire N__14137;
    wire N__14134;
    wire N__14133;
    wire N__14130;
    wire N__14123;
    wire N__14118;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14112;
    wire N__14111;
    wire N__14110;
    wire N__14109;
    wire N__14106;
    wire N__14103;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14076;
    wire N__14071;
    wire N__14064;
    wire N__14063;
    wire N__14062;
    wire N__14061;
    wire N__14060;
    wire N__14059;
    wire N__14058;
    wire N__14055;
    wire N__14042;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14018;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13976;
    wire N__13975;
    wire N__13974;
    wire N__13965;
    wire N__13964;
    wire N__13963;
    wire N__13962;
    wire N__13959;
    wire N__13952;
    wire N__13947;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13941;
    wire N__13940;
    wire N__13937;
    wire N__13936;
    wire N__13935;
    wire N__13932;
    wire N__13923;
    wire N__13916;
    wire N__13911;
    wire N__13910;
    wire N__13909;
    wire N__13908;
    wire N__13899;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13893;
    wire N__13886;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13871;
    wire N__13870;
    wire N__13869;
    wire N__13866;
    wire N__13865;
    wire N__13858;
    wire N__13855;
    wire N__13854;
    wire N__13853;
    wire N__13850;
    wire N__13845;
    wire N__13840;
    wire N__13833;
    wire N__13832;
    wire N__13831;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13818;
    wire N__13813;
    wire N__13810;
    wire N__13803;
    wire N__13800;
    wire N__13797;
    wire N__13794;
    wire N__13791;
    wire N__13790;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13782;
    wire N__13779;
    wire N__13778;
    wire N__13777;
    wire N__13774;
    wire N__13771;
    wire N__13766;
    wire N__13761;
    wire N__13758;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13727;
    wire N__13726;
    wire N__13725;
    wire N__13722;
    wire N__13721;
    wire N__13714;
    wire N__13711;
    wire N__13710;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13693;
    wire N__13686;
    wire N__13683;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13675;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13660;
    wire N__13657;
    wire N__13650;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13632;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13620;
    wire N__13619;
    wire N__13616;
    wire N__13613;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13600;
    wire N__13597;
    wire N__13590;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13579;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13563;
    wire N__13562;
    wire N__13561;
    wire N__13560;
    wire N__13559;
    wire N__13558;
    wire N__13557;
    wire N__13554;
    wire N__13541;
    wire N__13536;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13526;
    wire N__13523;
    wire N__13520;
    wire N__13517;
    wire N__13514;
    wire N__13509;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13492;
    wire N__13491;
    wire N__13486;
    wire N__13483;
    wire N__13480;
    wire N__13473;
    wire N__13470;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13464;
    wire N__13463;
    wire N__13460;
    wire N__13459;
    wire N__13456;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13436;
    wire N__13431;
    wire N__13428;
    wire N__13427;
    wire N__13426;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13418;
    wire N__13417;
    wire N__13414;
    wire N__13413;
    wire N__13410;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13383;
    wire N__13382;
    wire N__13377;
    wire N__13374;
    wire N__13373;
    wire N__13372;
    wire N__13371;
    wire N__13370;
    wire N__13369;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13350;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13336;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13297;
    wire N__13296;
    wire N__13295;
    wire N__13294;
    wire N__13293;
    wire N__13290;
    wire N__13287;
    wire N__13282;
    wire N__13275;
    wire N__13266;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13262;
    wire N__13257;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13242;
    wire N__13241;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13213;
    wire N__13208;
    wire N__13197;
    wire N__13194;
    wire N__13193;
    wire N__13190;
    wire N__13189;
    wire N__13188;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13180;
    wire N__13173;
    wire N__13168;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13112;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13104;
    wire N__13103;
    wire N__13102;
    wire N__13101;
    wire N__13100;
    wire N__13099;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13091;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13073;
    wire N__13070;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13054;
    wire N__13049;
    wire N__13042;
    wire N__13035;
    wire N__13034;
    wire N__13029;
    wire N__13028;
    wire N__13025;
    wire N__13022;
    wire N__13017;
    wire N__13016;
    wire N__13013;
    wire N__13010;
    wire N__13005;
    wire N__13002;
    wire N__13001;
    wire N__12996;
    wire N__12993;
    wire N__12992;
    wire N__12991;
    wire N__12990;
    wire N__12983;
    wire N__12982;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12968;
    wire N__12965;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12888;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12870;
    wire N__12869;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12822;
    wire N__12821;
    wire N__12818;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12790;
    wire N__12785;
    wire N__12778;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12656;
    wire N__12655;
    wire N__12648;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12642;
    wire N__12637;
    wire N__12634;
    wire N__12627;
    wire N__12626;
    wire N__12625;
    wire N__12624;
    wire N__12621;
    wire N__12620;
    wire N__12617;
    wire N__12616;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12604;
    wire N__12601;
    wire N__12598;
    wire N__12591;
    wire N__12586;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12563;
    wire N__12560;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12542;
    wire N__12539;
    wire N__12532;
    wire N__12529;
    wire N__12522;
    wire N__12519;
    wire N__12518;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12503;
    wire N__12500;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12482;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12464;
    wire N__12463;
    wire N__12460;
    wire N__12459;
    wire N__12454;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12437;
    wire N__12432;
    wire N__12431;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12401;
    wire N__12398;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12365;
    wire N__12364;
    wire N__12361;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12308;
    wire N__12307;
    wire N__12306;
    wire N__12305;
    wire N__12302;
    wire N__12299;
    wire N__12296;
    wire N__12293;
    wire N__12288;
    wire N__12279;
    wire N__12276;
    wire N__12275;
    wire N__12274;
    wire N__12273;
    wire N__12268;
    wire N__12263;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12250;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12177;
    wire N__12174;
    wire N__12173;
    wire N__12170;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12137;
    wire N__12132;
    wire N__12131;
    wire N__12128;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12111;
    wire N__12108;
    wire N__12107;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12099;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12084;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12045;
    wire N__12042;
    wire N__12033;
    wire N__12028;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12005;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11934;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11920;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11897;
    wire N__11894;
    wire N__11891;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11757;
    wire N__11754;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11708;
    wire N__11705;
    wire N__11704;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11697;
    wire N__11694;
    wire N__11693;
    wire N__11690;
    wire N__11685;
    wire N__11680;
    wire N__11671;
    wire N__11666;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11647;
    wire N__11646;
    wire N__11645;
    wire N__11638;
    wire N__11633;
    wire N__11630;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11591;
    wire N__11588;
    wire N__11587;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11553;
    wire N__11552;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11493;
    wire N__11490;
    wire N__11483;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11435;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11425;
    wire N__11420;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11389;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11371;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11311;
    wire N__11306;
    wire N__11303;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11291;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11216;
    wire N__11215;
    wire N__11210;
    wire N__11207;
    wire N__11202;
    wire N__11199;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11184;
    wire N__11183;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11175;
    wire N__11172;
    wire N__11165;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11100;
    wire N__11097;
    wire N__11096;
    wire N__11095;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11049;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11008;
    wire N__11003;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10957;
    wire N__10954;
    wire N__10949;
    wire N__10944;
    wire N__10943;
    wire N__10940;
    wire N__10939;
    wire N__10936;
    wire N__10931;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10898;
    wire N__10897;
    wire N__10894;
    wire N__10889;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10873;
    wire N__10868;
    wire N__10863;
    wire N__10862;
    wire N__10861;
    wire N__10858;
    wire N__10853;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10835;
    wire N__10834;
    wire N__10831;
    wire N__10826;
    wire N__10821;
    wire N__10820;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10808;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10700;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10658;
    wire N__10657;
    wire N__10654;
    wire N__10649;
    wire N__10644;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10632;
    wire N__10629;
    wire N__10628;
    wire N__10623;
    wire N__10620;
    wire N__10619;
    wire N__10618;
    wire N__10617;
    wire N__10616;
    wire N__10611;
    wire N__10606;
    wire N__10603;
    wire N__10600;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10582;
    wire N__10579;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10500;
    wire N__10497;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10485;
    wire N__10482;
    wire N__10479;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10451;
    wire N__10446;
    wire N__10443;
    wire N__10442;
    wire N__10441;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10426;
    wire N__10419;
    wire N__10416;
    wire N__10415;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10391;
    wire N__10390;
    wire N__10389;
    wire N__10388;
    wire N__10385;
    wire N__10376;
    wire N__10371;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10363;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10349;
    wire N__10344;
    wire N__10343;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10328;
    wire N__10327;
    wire N__10324;
    wire N__10323;
    wire N__10320;
    wire N__10315;
    wire N__10312;
    wire N__10311;
    wire N__10306;
    wire N__10301;
    wire N__10298;
    wire N__10293;
    wire N__10292;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10274;
    wire N__10273;
    wire N__10270;
    wire N__10269;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10248;
    wire N__10247;
    wire N__10244;
    wire N__10243;
    wire N__10242;
    wire N__10239;
    wire N__10238;
    wire N__10235;
    wire N__10230;
    wire N__10225;
    wire N__10220;
    wire N__10215;
    wire N__10214;
    wire N__10213;
    wire N__10210;
    wire N__10209;
    wire N__10208;
    wire N__10207;
    wire N__10202;
    wire N__10199;
    wire N__10192;
    wire N__10189;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10169;
    wire N__10168;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10156;
    wire N__10153;
    wire N__10146;
    wire N__10143;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10139;
    wire N__10138;
    wire N__10135;
    wire N__10124;
    wire N__10119;
    wire N__10116;
    wire N__10115;
    wire N__10114;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10106;
    wire N__10101;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10080;
    wire N__10077;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10069;
    wire N__10068;
    wire N__10063;
    wire N__10058;
    wire N__10053;
    wire N__10050;
    wire N__10047;
    wire N__10046;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10029;
    wire N__10028;
    wire N__10025;
    wire N__10024;
    wire N__10021;
    wire N__10020;
    wire N__10017;
    wire N__10010;
    wire N__10005;
    wire N__10002;
    wire N__9999;
    wire N__9996;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9984;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9932;
    wire N__9929;
    wire N__9926;
    wire N__9923;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9879;
    wire N__9872;
    wire N__9867;
    wire N__9866;
    wire N__9865;
    wire N__9864;
    wire N__9861;
    wire N__9860;
    wire N__9859;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9848;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9844;
    wire N__9841;
    wire N__9838;
    wire N__9833;
    wire N__9826;
    wire N__9815;
    wire N__9804;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9740;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9725;
    wire N__9724;
    wire N__9723;
    wire N__9720;
    wire N__9719;
    wire N__9716;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9700;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9659;
    wire N__9654;
    wire N__9653;
    wire N__9652;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9616;
    wire N__9611;
    wire N__9606;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9598;
    wire N__9597;
    wire N__9594;
    wire N__9587;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9545;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9537;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9522;
    wire N__9513;
    wire N__9510;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9500;
    wire N__9495;
    wire N__9492;
    wire N__9491;
    wire N__9490;
    wire N__9489;
    wire N__9484;
    wire N__9479;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9465;
    wire N__9462;
    wire N__9461;
    wire N__9460;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9440;
    wire N__9439;
    wire N__9438;
    wire N__9437;
    wire N__9436;
    wire N__9431;
    wire N__9424;
    wire N__9421;
    wire N__9414;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9402;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9381;
    wire N__9378;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9368;
    wire N__9365;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9350;
    wire N__9347;
    wire N__9340;
    wire N__9339;
    wire N__9336;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9318;
    wire N__9317;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9308;
    wire N__9301;
    wire N__9298;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9281;
    wire N__9280;
    wire N__9279;
    wire N__9272;
    wire N__9269;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9225;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9214;
    wire N__9213;
    wire N__9210;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9178;
    wire N__9175;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9118;
    wire N__9109;
    wire N__9100;
    wire N__9093;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9089;
    wire N__9088;
    wire N__9085;
    wire N__9074;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9066;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9050;
    wire N__9049;
    wire N__9046;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9032;
    wire N__9029;
    wire N__9024;
    wire N__9023;
    wire N__9020;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9003;
    wire N__9002;
    wire N__9001;
    wire N__9000;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8984;
    wire N__8981;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8960;
    wire N__8957;
    wire N__8956;
    wire N__8955;
    wire N__8946;
    wire N__8943;
    wire N__8942;
    wire N__8941;
    wire N__8936;
    wire N__8933;
    wire N__8928;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8913;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8900;
    wire N__8897;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8877;
    wire N__8874;
    wire N__8873;
    wire N__8872;
    wire N__8871;
    wire N__8870;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8850;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8833;
    wire N__8828;
    wire N__8823;
    wire N__8820;
    wire N__8819;
    wire N__8816;
    wire N__8815;
    wire N__8814;
    wire N__8811;
    wire N__8804;
    wire N__8801;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8779;
    wire N__8772;
    wire N__8771;
    wire N__8770;
    wire N__8769;
    wire N__8764;
    wire N__8759;
    wire N__8754;
    wire N__8751;
    wire N__8750;
    wire N__8749;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8724;
    wire N__8721;
    wire N__8720;
    wire N__8719;
    wire N__8718;
    wire N__8717;
    wire N__8710;
    wire N__8705;
    wire N__8700;
    wire N__8699;
    wire N__8698;
    wire N__8697;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8669;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8657;
    wire N__8646;
    wire N__8643;
    wire N__8642;
    wire N__8641;
    wire N__8636;
    wire N__8633;
    wire N__8628;
    wire N__8625;
    wire N__8624;
    wire N__8623;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8546;
    wire N__8545;
    wire N__8542;
    wire N__8537;
    wire N__8534;
    wire N__8529;
    wire N__8526;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8399;
    wire N__8396;
    wire N__8395;
    wire N__8394;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8380;
    wire N__8373;
    wire N__8370;
    wire N__8367;
    wire N__8364;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8313;
    wire N__8310;
    wire N__8309;
    wire N__8308;
    wire N__8307;
    wire N__8304;
    wire N__8297;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8282;
    wire N__8281;
    wire N__8278;
    wire N__8277;
    wire N__8276;
    wire N__8273;
    wire N__8264;
    wire N__8259;
    wire N__8258;
    wire N__8257;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8238;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8230;
    wire N__8229;
    wire N__8226;
    wire N__8221;
    wire N__8218;
    wire N__8213;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8203;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8186;
    wire N__8185;
    wire N__8178;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8162;
    wire N__8161;
    wire N__8158;
    wire N__8153;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8136;
    wire N__8135;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire \latticehx1k_pll_inst.clk ;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire uart_RXD;
    wire \uu0.un165_ci_0_cascade_ ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.un99_ci_0 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.un44_ci ;
    wire \uu0.un44_ci_cascade_ ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un66_ci_cascade_ ;
    wire \uu0.un66_ci ;
    wire \uu0.un88_ci_3 ;
    wire bfn_1_11_0_;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire \buart.Z_rx.valid_0_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_rx.idle_0_cascade_ ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.un350_ci ;
    wire \uu2.un350_ci_cascade_ ;
    wire \uu2.vbuf_count.un328_ci_3_cascade_ ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu2.un1_l_count_1_3_cascade_ ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.un1_l_count_1_0 ;
    wire \uu0.un198_ci_2 ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.un1_l_count_2_2 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu0.un187_ci_1 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.un143_ci_0_cascade_ ;
    wire \uu0.un110_ci ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.un4_l_count_13_cascade_ ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un4_l_count_16 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.l_precountZ0Z_1 ;
    wire CONSTANT_ONE_NET_cascade_;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un11_l_count_i ;
    wire \uu2.mem0.w_addr_0 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \resetGen.un241_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_1 ;
    wire \resetGen.reset_countZ0Z_0 ;
    wire \resetGen.un252_ci_cascade_ ;
    wire \resetGen.reset_countZ0Z_3 ;
    wire \resetGen.reset_countZ0Z_2 ;
    wire \resetGen.un241_ci ;
    wire \resetGen.reset_count_2_0_4_cascade_ ;
    wire \resetGen.reset_countZ0Z_4 ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.sample ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire bfn_2_13_0_;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.un404_ci_0_cascade_ ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.mem0.w_data_5 ;
    wire \uu2.N_34 ;
    wire \uu2.N_34_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.N_31 ;
    wire \uu2.N_31_cascade_ ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \INVuu2.vram_rd_clk_det_0C_net ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci_0 ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.un284_ci ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire G_188;
    wire G_188_cascade_;
    wire \Lab_UT.un1_rst_0_iclkZ0 ;
    wire G_182_cascade_;
    wire G_187;
    wire \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ;
    wire G_183;
    wire G_182;
    wire \uu2.l_countZ0Z_0 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \uu2.mem0.w_addr_8 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire \uu2.un28_w_addr_user_i_cascade_ ;
    wire \uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_15_cascade_ ;
    wire \INVuu2.w_addr_displaying_1_rep1_nesrC_net ;
    wire \uu2.N_401 ;
    wire \uu2.N_406_cascade_ ;
    wire \uu2.bitmap_pmux ;
    wire \uu2.N_383_cascade_ ;
    wire \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ;
    wire \uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ;
    wire \uu2.bitmap_pmux_sn_i5_mux ;
    wire \uu2.bitmap_pmux_u_1 ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ;
    wire \uu2.w_addr_displaying_RNI0NG56Z0Z_4 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \INVuu2.vram_rd_clk_det_1C_net ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ;
    wire \uu2.un20_w_addr_userZ0Z_1 ;
    wire L3_tx_data_rdy;
    wire \Lab_UT.dispString.N_124_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ;
    wire \Lab_UT.didp.regrce4.LdAMtens_0 ;
    wire \uu2.un1_w_user_lfZ0Z_4 ;
    wire L3_tx_data_5;
    wire \uu2.un1_w_user_crZ0Z_4 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_3 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_3 ;
    wire \uu2.un1_w_user_lfZ0Z_3 ;
    wire L3_tx_data_3;
    wire L3_tx_data_0;
    wire \uu2.un1_w_user_crZ0Z_3 ;
    wire \Lab_UT.dispString.dOutP_1_iv_i_1_4 ;
    wire L3_tx_data_4;
    wire \Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ;
    wire G_186;
    wire L3_tx_data_6;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.un1_armed_2_0_iso_iZ0 ;
    wire \Lab_UT.un1_idle_4_0_iclkZ0_cascade_ ;
    wire G_185;
    wire G_185_cascade_;
    wire \Lab_UT.dispString.N_117_cascade_ ;
    wire L3_tx_data_1;
    wire \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ;
    wire G_180_cascade_;
    wire G_181_cascade_;
    wire G_180;
    wire \Lab_UT.dictrl.alarmstate_1_0_cascade_ ;
    wire \Lab_UT.alarmstate_0_sqmuxa_1 ;
    wire \Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ;
    wire G_184;
    wire \resetGen.escKeyZ0Z_5_cascade_ ;
    wire \resetGen.escKeyZ0 ;
    wire \resetGen.escKeyZ0Z_4 ;
    wire \uu2.un28_w_addr_user_i ;
    wire \INVuu2.w_addr_user_2C_net ;
    wire \uu2.un51_w_data_displaying_i_a2_1 ;
    wire \uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ;
    wire \uu2.w_data_displaying_2_i_a2_i_a3_2_0 ;
    wire \INVuu2.w_addr_displaying_nesr_3C_net ;
    wire \uu2.bitmap_pmux_sn_N_33 ;
    wire \uu2.w_addr_displaying_RNI03P31Z0Z_4 ;
    wire \uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ;
    wire \uu2.bitmap_pmux_sn_i7_mux_0 ;
    wire \INVuu2.bitmap_93C_net ;
    wire \uu2.w_addr_displaying_1_repZ0Z1 ;
    wire \uu2.N_24_cascade_ ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.N_31_i ;
    wire \uu2.N_26_cascade_ ;
    wire \uu2.bitmap_pmux_27_ns_1 ;
    wire \uu2.N_404 ;
    wire \Lab_UT.didp.ce_12_1 ;
    wire \Lab_UT.didp.ce_12_1_cascade_ ;
    wire \Lab_UT.didp.ce_12_3_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_1 ;
    wire \Lab_UT.dispString.N_140 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ;
    wire \Lab_UT.didp.countrce1.un20_qPone ;
    wire \Lab_UT.didp.countrce1.q_5_3_cascade_ ;
    wire \Lab_UT.dispString.N_137 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ;
    wire \Lab_UT.didp.countrce4.q_5_3_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_2_2 ;
    wire \Lab_UT.didp.countrce4.q_5_0_cascade_ ;
    wire G_181;
    wire G_179;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0 ;
    wire \Lab_UT.dispString.un42_dOutP_1 ;
    wire \Lab_UT.dispString.N_95 ;
    wire \Lab_UT.didp.regrce2.LdAStens_0 ;
    wire \Lab_UT.dictrl.alarmstateZ0Z8 ;
    wire \Lab_UT.dictrl.m37_N_2LZ0Z1 ;
    wire \Lab_UT.dictrl.g1_0Z0Z_5 ;
    wire \Lab_UT.dictrl.g1_0_4_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_5_4_0 ;
    wire \Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.g0_5_3_0 ;
    wire \Lab_UT.dictrl.G_25_i_o3_3_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate8Z0Z_3 ;
    wire \INVuu2.w_addr_displaying_ness_6C_net ;
    wire \uu2.N_33_1 ;
    wire \uu2.mem0.w_addr_6 ;
    wire \uu2.mem0.w_addr_4 ;
    wire \uu2.mem0.w_addr_5 ;
    wire \uu2.mem0.w_addr_7 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \INVuu2.bitmap_168C_net ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.w_addr_displaying_fastZ0Z_1 ;
    wire \uu2.bitmap_pmux_sn_N_54_mux_cascade_ ;
    wire \uu2.N_14 ;
    wire \uu2.bitmap_RNI2Q8F1Z0Z_111 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \uu2.N_166 ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \INVuu2.bitmap_197C_net ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \uu2.N_149 ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.N_25 ;
    wire \Lab_UT.didp.countrce1.ce_12_1_1 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.didp.countrce4.un20_qPone ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.didp.countrce2.N_93 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ;
    wire \Lab_UT.didp.countrce2.N_96_cascade_ ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_3 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_1 ;
    wire \Lab_UT.di_Stens_3 ;
    wire \Lab_UT.didp.un24_ce_3 ;
    wire \Lab_UT.dispString.N_143 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_1_0 ;
    wire \Lab_UT.didp.un1_dicLdStens_0 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_2 ;
    wire \Lab_UT.didp.un1_dicLdStens_0_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \Lab_UT.didp.countrce1.q_5_0 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ;
    wire \Lab_UT.didp.N_90 ;
    wire \Lab_UT.LdSones_i_4 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.state_ret_8_ess ;
    wire \Lab_UT.di_Stens_0 ;
    wire \Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ;
    wire \Lab_UT.didp.countrce1.q_5_1 ;
    wire \Lab_UT.didp.regrce1.LdASones_0 ;
    wire \Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_ ;
    wire \Lab_UT.dictrl.G_25_i_a5_1_0_cascade_ ;
    wire \Lab_UT.i8_mux_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_0_sn ;
    wire \Lab_UT.dictrl.g1_1_0_1_cascade_ ;
    wire \Lab_UT.g1 ;
    wire \Lab_UT.dictrl.g0_0_rn_0 ;
    wire \Lab_UT.dictrl.G_25_i_0 ;
    wire \Lab_UT.dictrl.G_25_i_1 ;
    wire \Lab_UT.dictrl.g2Z0Z_0 ;
    wire \Lab_UT.dictrl.g0_6_3_0 ;
    wire \Lab_UT.dictrl.m13_out_cascade_ ;
    wire \Lab_UT.dictrl.N_18_0_0_cascade_ ;
    wire \Lab_UT.dictrl.G_25_i_o3_5 ;
    wire \Lab_UT.dictrl.G_25_i_o3_4 ;
    wire \Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ;
    wire \Lab_UT.dictrl.N_11 ;
    wire \Lab_UT.dictrl.m34Z0Z_1_cascade_ ;
    wire bu_rx_data_6;
    wire \Lab_UT.dictrl.m22Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.N_72_mux_1 ;
    wire \Lab_UT.dictrl.g1_1_0_0 ;
    wire \Lab_UT.dictrl.m22Z0Z_1 ;
    wire \Lab_UT.dictrl.g1_1_0 ;
    wire \Lab_UT.dictrl.g1_rn_0 ;
    wire \Lab_UT.dictrl.m34Z0Z_1 ;
    wire bu_rx_data_fast_3;
    wire bu_rx_data_fast_0;
    wire \Lab_UT.dictrl.g1_1_4_cascade_ ;
    wire \Lab_UT.dictrl.g1_1Z0Z_5 ;
    wire bu_rx_data_7;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire bu_rx_data_fast_7;
    wire \uu2.N_40 ;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ;
    wire \INVuu2.w_addr_displaying_fast_8C_net ;
    wire \uu2.N_37 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.N_45 ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.bitmap_pmux_sn_N_36 ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmap_pmux_20_ns_1 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.bitmap_pmux_26_bm_1 ;
    wire \uu2.bitmap_RNIP2JO1Z0Z_34 ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \INVuu2.bitmap_290C_net ;
    wire \Lab_UT.di_Sones_3 ;
    wire \Lab_UT.di_ASones_3 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.min1_0 ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.di_Mtens_3 ;
    wire \Lab_UT.min1_3 ;
    wire \Lab_UT.sec1_3 ;
    wire \Lab_UT.sec1_0 ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \uu2.bitmap_pmux_17_ns_1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.bitmap_pmux_16_ns_1 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \Lab_UT.min2_0 ;
    wire \Lab_UT.min2_3 ;
    wire \Lab_UT.min2_2 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \INVuu2.bitmap_215C_net ;
    wire \Lab_UT.di_Stens_1 ;
    wire \Lab_UT.sec1_1 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.min1_1 ;
    wire \Lab_UT.di_Stens_2 ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.sec1_2 ;
    wire \Lab_UT.di_Sones_0 ;
    wire \Lab_UT.LdSones ;
    wire \Lab_UT.didp.countrce1.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.didp.countrce1.q_5_2_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdSones_0 ;
    wire \Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ;
    wire \Lab_UT.min2_1 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.min1_2 ;
    wire \Lab_UT.didp.regrce3.LdAMones_0 ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.dispString.N_118_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_i_0_1 ;
    wire \Lab_UT.dispString.N_145 ;
    wire \Lab_UT.dictrl.dicLdAMones_1 ;
    wire \Lab_UT.LdAMones ;
    wire \Lab_UT.LdAMones_cascade_ ;
    wire \Lab_UT.dictrl.g0_1_mb_rn_0 ;
    wire \Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ;
    wire \Lab_UT.dictrl.N_57_1 ;
    wire \Lab_UT.dictrl.N_55_1 ;
    wire \Lab_UT.dictrl.next_state_0_2 ;
    wire \Lab_UT.dictrl.next_state_1_2_cascade_ ;
    wire \Lab_UT.dictrl.g0_1_mb_sn ;
    wire \Lab_UT.dictrl.un15_loadalarm_0_cascade_ ;
    wire \Lab_UT.dictrl.loadalarm_0_0 ;
    wire \Lab_UT.LdAStens ;
    wire \Lab_UT.dictrl.N_22 ;
    wire \Lab_UT.dictrl.next_state_0_1 ;
    wire \Lab_UT.dictrl.g2_0_0 ;
    wire \Lab_UT.dictrl.state_i_4_2 ;
    wire \Lab_UT.dictrl.N_20_0_0_cascade_ ;
    wire \Lab_UT.dictrl.N_22_0_0 ;
    wire \Lab_UT.next_state_0 ;
    wire \Lab_UT.next_state_1_0_0_1_cascade_ ;
    wire \Lab_UT.next_state_2 ;
    wire bu_rx_data_rdy;
    wire \Lab_UT.didp.g0_0_2Z0Z_1 ;
    wire rst;
    wire \Lab_UT.didp.g0_0Z0Z_2 ;
    wire \Lab_UT.dictrl.next_state6 ;
    wire \Lab_UT.dictrl.N_20_cascade_ ;
    wire \Lab_UT.dictrl.m34_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_3_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_3 ;
    wire \Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ;
    wire \Lab_UT.dictrl.N_26_0 ;
    wire \Lab_UT.dictrl.m34_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.N_60_0_0 ;
    wire \Lab_UT.dictrl.m19_1 ;
    wire N_5_cascade_;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ;
    wire \Lab_UT.dictrl.N_59_1_0 ;
    wire \Lab_UT.dictrl.i8_mux_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13 ;
    wire \Lab_UT.dictrl.m22_xZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.m22Z0Z_4 ;
    wire \Lab_UT.dictrl.N_72_mux_cascade_ ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.N_18 ;
    wire m7_a0;
    wire \Lab_UT.dictrl.state_fast_0 ;
    wire buart__rx_shifter_fast_4;
    wire bu_rx_data_5_rep1;
    wire \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_6_3 ;
    wire \Lab_UT.dictrl.gZ0Z2 ;
    wire \Lab_UT.dictrl.g0_6_3_cascade_ ;
    wire \Lab_UT.dictrl.g1_1 ;
    wire \Lab_UT.dictrl.N_57_0 ;
    wire bu_rx_data_fast_6;
    wire bu_rx_data_fast_5;
    wire \Lab_UT.dictrl.g1_0_4_cascade_ ;
    wire \Lab_UT.dictrl.g1_0_xZ0Z1 ;
    wire \Lab_UT.dictrl.g0_5Z0Z_4 ;
    wire \Lab_UT.dictrl.g0_5_3 ;
    wire \Lab_UT.dictrl.g1_0_cascade_ ;
    wire \Lab_UT.dictrl.N_55_0 ;
    wire \Lab_UT.dictrl.g0_3_4_cascade_ ;
    wire bu_rx_data_5;
    wire \Lab_UT.dictrl.N_72_mux_0 ;
    wire bu_rx_data_6_rep1;
    wire bu_rx_data_7_rep1;
    wire \Lab_UT.dictrl.g0_3_3 ;
    wire bu_rx_data_4;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.un3_w_addr_user_4_cascade_ ;
    wire \uu2.un3_w_addr_user_5 ;
    wire \uu2.un3_w_addr_user ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.un404_ci_cascade_ ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.mem0.w_addr_3 ;
    wire \uu2.un426_ci_3 ;
    wire \uu2.un404_ci ;
    wire \uu2.vbuf_w_addr_user.un448_ci_0 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \INVuu2.w_addr_user_nesr_3C_net ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.w_addr_user_RNI43E87Z0Z_4 ;
    wire \uu2.N_44 ;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_8 ;
    wire \uu2.bitmapZ0Z_111 ;
    wire \INVuu2.w_addr_displaying_7C_net ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.w_addr_displaying_0_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmap_pmux_19_ns_1 ;
    wire \Lab_UT.sec2_0 ;
    wire \Lab_UT.sec2_3 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.N_152_cascade_ ;
    wire \uu2.w_addr_displaying_fastZ0Z_8 ;
    wire \uu2.bitmap_RNIM5E21Z0Z_314 ;
    wire \Lab_UT.didp.countrce3.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_2_cascade_ ;
    wire \Lab_UT.didp.reset_12_1_3 ;
    wire \Lab_UT.di_Mones_2 ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire \Lab_UT.di_Mones_3 ;
    wire \Lab_UT.didp.countrce3.q_5_3 ;
    wire \Lab_UT.didp.un1_dicLdMones_0 ;
    wire \Lab_UT.didp.un1_dicLdMones_0_cascade_ ;
    wire \Lab_UT.dispString.N_144 ;
    wire \Lab_UT.di_Mtens_0 ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.di_Mtens_1 ;
    wire \Lab_UT.di_Sones_2 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.sec2_2 ;
    wire \Lab_UT.di_Mones_1 ;
    wire \Lab_UT.didp.countrce3.q_5_1 ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.didp.un1_dicLdMtens_0 ;
    wire \Lab_UT.di_Sones_1 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.loadalarm_0 ;
    wire \Lab_UT.sec2_1 ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.countrce4.un13_qPone ;
    wire \Lab_UT.di_Mtens_2 ;
    wire \Lab_UT.didp.countrce4.q_5_2 ;
    wire uu0_sec_clkD;
    wire o_One_Sec_Pulse;
    wire oneSecStrb;
    wire oneSecStrb_cascade_;
    wire \Lab_UT.dispString.N_102 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.di_Mones_0 ;
    wire \Lab_UT.dictrl.state_i_3_0 ;
    wire \Lab_UT.dictrl.state_ret_2_fast ;
    wire \Lab_UT.dictrl.N_20 ;
    wire \Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ;
    wire \Lab_UT.dictrl.state_i_4_1 ;
    wire \Lab_UT.dictrl.m19_1_0 ;
    wire \Lab_UT.dictrl.next_state_1_3 ;
    wire \Lab_UT.dictrl.next_state_0_3 ;
    wire \Lab_UT.next_state_1 ;
    wire \Lab_UT.dictrl.next_state66_2 ;
    wire \Lab_UT.bu_rx_data_rdy_0 ;
    wire \Lab_UT.state_i_4_3 ;
    wire \Lab_UT.dictrl.dicRun_1 ;
    wire \Lab_UT.state_2 ;
    wire \Lab_UT.LdASones ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire \Lab_UT.dictrl.g1_4_0 ;
    wire \Lab_UT.dictrl.g1_5_0_cascade_ ;
    wire \Lab_UT.dictrl.G_14_0_a2_4_2_cascade_ ;
    wire \Lab_UT.dictrl.G_14_0_0 ;
    wire shifter_1_rep1_RNI0FPF_cascade_;
    wire \Lab_UT.dictrl.N_33_0 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ;
    wire \Lab_UT.dictrl.G_14_0_1 ;
    wire bu_rx_data_3_rep1;
    wire \Lab_UT.dictrl.G_14_0_a2_1 ;
    wire N_15_cascade_;
    wire \Lab_UT.dictrl.N_20_0 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ;
    wire \Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ;
    wire \Lab_UT.g0_0 ;
    wire \Lab_UT.dictrl.N_15_0_cascade_ ;
    wire \Lab_UT.dictrl.N_60_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ;
    wire \Lab_UT.dictrl.next_state_0_0 ;
    wire \Lab_UT.un1_next_state66_0 ;
    wire \Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ;
    wire \Lab_UT.dictrl.N_60 ;
    wire \Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ;
    wire \Lab_UT.dicLdSones_1 ;
    wire G_6_0_a6_2_cascade_;
    wire \Lab_UT.dictrl.G_6_0_0_1 ;
    wire \Lab_UT.dictrl.G_6_0_0_cascade_ ;
    wire \Lab_UT.dictrl.G_6_0_1_0 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ;
    wire \Lab_UT.dictrl.m13_out ;
    wire \Lab_UT.dictrl.N_15_0 ;
    wire \Lab_UT.dictrl.N_72_mux ;
    wire \Lab_UT.dictrl.N_59 ;
    wire \Lab_UT.dictrl.N_8_0 ;
    wire \Lab_UT.dictrl.i8_mux ;
    wire bu_rx_data_fast_2;
    wire \Lab_UT.dictrl.state_0_rep1 ;
    wire \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_ ;
    wire \Lab_UT.dictrl.N_3 ;
    wire bu_rx_data_0;
    wire \Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.next_state_RNO_5Z0Z_0 ;
    wire \Lab_UT.dictrl.i9_mux ;
    wire Lab_UT_dictrl_state_1;
    wire bu_rx_data_2_rep1;
    wire bu_rx_data_0_rep1;
    wire \Lab_UT.dictrl.N_67_mux ;
    wire \Lab_UT.dictrl.stateZ0Z_3 ;
    wire G_6_0_a6_3_3_cascade_;
    wire \Lab_UT.stateZ0Z_0 ;
    wire \Lab_UT.dictrl.N_12 ;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_1_rep1;
    wire N_63_mux;
    wire bu_rx_data_1;
    wire bu_rx_data_3_rep2;
    wire N_14_0;
    wire bu_rx_data_3;
    wire bu_rx_data_2;
    wire \buart.Z_rx.sample_g ;
    wire rst_g;
    wire vbuf_tx_data_rdy;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \uu2.mem0.w_addr_1 ;
    wire L3_tx_data_2;
    wire \uu2.mem0.w_data_2 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.un4_w_user_data_rdyZ0Z_0 ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.mem0.w_addr_2 ;
    wire \buart.Z_tx.un1_bitcount_c2 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0_cascade_ ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.un1_bitcount_c3 ;
    wire bfn_12_2_0_;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire clk_g;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \buart.Z_tx.ser_clk ;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(\latticehx1k_pll_inst.clk ),
            .REFERENCECLK(N__8085),
            .RESETB(N__11095),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__9780,N__10050,N__10029,N__10482,N__10116,N__9759,N__10275,N__10248,N__10215}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__10533,N__11826,N__11865,N__11838,N__11850,N__16056,N__21627,N__20241,N__9582}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__9999,dangling_wire_31,N__9993,dangling_wire_32,N__9966,dangling_wire_33,N__9978,dangling_wire_34,N__21855,dangling_wire_35,N__9972,dangling_wire_36,N__10281}),
            .RCLKE(),
            .RCLK(N__22269),
            .RE(N__11100),
            .WCLKE(N__10517),
            .WCLK(N__22268),
            .WE(N__10521));
    IO_PAD led_obuft_3_iopad (
            .OE(N__22396),
            .DIN(N__22395),
            .DOUT(N__22394),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__22396),
            .PADOUT(N__22395),
            .PADIN(N__22394),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__22387),
            .DIN(N__22386),
            .DOUT(N__22385),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__22387),
            .PADOUT(N__22386),
            .PADIN(N__22385),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__22378),
            .DIN(N__22377),
            .DOUT(N__22376),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__22378),
            .PADOUT(N__22377),
            .PADIN(N__22376),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__22369),
            .DIN(N__22368),
            .DOUT(N__22367),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__22369),
            .PADOUT(N__22368),
            .PADIN(N__22367),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__22223),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__22360),
            .DIN(N__22359),
            .DOUT(N__22358),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__22360),
            .PADOUT(N__22359),
            .PADIN(N__22358),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__22351),
            .DIN(N__22350),
            .DOUT(N__22349),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__22351),
            .PADOUT(N__22350),
            .PADIN(N__22349),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__22342),
            .DIN(N__22341),
            .DOUT(N__22340),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__22342),
            .PADOUT(N__22341),
            .PADIN(N__22340),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__22333),
            .DIN(N__22332),
            .DOUT(N__22331),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__22333),
            .PADOUT(N__22332),
            .PADIN(N__22331),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__22324),
            .DIN(N__22323),
            .DOUT(N__22322),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__22324),
            .PADOUT(N__22323),
            .PADIN(N__22322),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__22315),
            .DIN(N__22314),
            .DOUT(N__22313),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__22315),
            .PADOUT(N__22314),
            .PADIN(N__22313),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5423 (
            .O(N__22296),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__5422 (
            .O(N__22293),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__5421 (
            .O(N__22290),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__5420 (
            .O(N__22287),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__5419 (
            .O(N__22284),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__5418 (
            .O(N__22281),
            .I(N__22278));
    InMux I__5417 (
            .O(N__22278),
            .I(N__22275));
    LocalMux I__5416 (
            .O(N__22275),
            .I(N__22185));
    ClkMux I__5415 (
            .O(N__22274),
            .I(N__22008));
    ClkMux I__5414 (
            .O(N__22273),
            .I(N__22008));
    ClkMux I__5413 (
            .O(N__22272),
            .I(N__22008));
    ClkMux I__5412 (
            .O(N__22271),
            .I(N__22008));
    ClkMux I__5411 (
            .O(N__22270),
            .I(N__22008));
    ClkMux I__5410 (
            .O(N__22269),
            .I(N__22008));
    ClkMux I__5409 (
            .O(N__22268),
            .I(N__22008));
    ClkMux I__5408 (
            .O(N__22267),
            .I(N__22008));
    ClkMux I__5407 (
            .O(N__22266),
            .I(N__22008));
    ClkMux I__5406 (
            .O(N__22265),
            .I(N__22008));
    ClkMux I__5405 (
            .O(N__22264),
            .I(N__22008));
    ClkMux I__5404 (
            .O(N__22263),
            .I(N__22008));
    ClkMux I__5403 (
            .O(N__22262),
            .I(N__22008));
    ClkMux I__5402 (
            .O(N__22261),
            .I(N__22008));
    ClkMux I__5401 (
            .O(N__22260),
            .I(N__22008));
    ClkMux I__5400 (
            .O(N__22259),
            .I(N__22008));
    ClkMux I__5399 (
            .O(N__22258),
            .I(N__22008));
    ClkMux I__5398 (
            .O(N__22257),
            .I(N__22008));
    ClkMux I__5397 (
            .O(N__22256),
            .I(N__22008));
    ClkMux I__5396 (
            .O(N__22255),
            .I(N__22008));
    ClkMux I__5395 (
            .O(N__22254),
            .I(N__22008));
    ClkMux I__5394 (
            .O(N__22253),
            .I(N__22008));
    ClkMux I__5393 (
            .O(N__22252),
            .I(N__22008));
    ClkMux I__5392 (
            .O(N__22251),
            .I(N__22008));
    ClkMux I__5391 (
            .O(N__22250),
            .I(N__22008));
    ClkMux I__5390 (
            .O(N__22249),
            .I(N__22008));
    ClkMux I__5389 (
            .O(N__22248),
            .I(N__22008));
    ClkMux I__5388 (
            .O(N__22247),
            .I(N__22008));
    ClkMux I__5387 (
            .O(N__22246),
            .I(N__22008));
    ClkMux I__5386 (
            .O(N__22245),
            .I(N__22008));
    ClkMux I__5385 (
            .O(N__22244),
            .I(N__22008));
    ClkMux I__5384 (
            .O(N__22243),
            .I(N__22008));
    ClkMux I__5383 (
            .O(N__22242),
            .I(N__22008));
    ClkMux I__5382 (
            .O(N__22241),
            .I(N__22008));
    ClkMux I__5381 (
            .O(N__22240),
            .I(N__22008));
    ClkMux I__5380 (
            .O(N__22239),
            .I(N__22008));
    ClkMux I__5379 (
            .O(N__22238),
            .I(N__22008));
    ClkMux I__5378 (
            .O(N__22237),
            .I(N__22008));
    ClkMux I__5377 (
            .O(N__22236),
            .I(N__22008));
    ClkMux I__5376 (
            .O(N__22235),
            .I(N__22008));
    ClkMux I__5375 (
            .O(N__22234),
            .I(N__22008));
    ClkMux I__5374 (
            .O(N__22233),
            .I(N__22008));
    ClkMux I__5373 (
            .O(N__22232),
            .I(N__22008));
    ClkMux I__5372 (
            .O(N__22231),
            .I(N__22008));
    ClkMux I__5371 (
            .O(N__22230),
            .I(N__22008));
    ClkMux I__5370 (
            .O(N__22229),
            .I(N__22008));
    ClkMux I__5369 (
            .O(N__22228),
            .I(N__22008));
    ClkMux I__5368 (
            .O(N__22227),
            .I(N__22008));
    ClkMux I__5367 (
            .O(N__22226),
            .I(N__22008));
    ClkMux I__5366 (
            .O(N__22225),
            .I(N__22008));
    ClkMux I__5365 (
            .O(N__22224),
            .I(N__22008));
    ClkMux I__5364 (
            .O(N__22223),
            .I(N__22008));
    ClkMux I__5363 (
            .O(N__22222),
            .I(N__22008));
    ClkMux I__5362 (
            .O(N__22221),
            .I(N__22008));
    ClkMux I__5361 (
            .O(N__22220),
            .I(N__22008));
    ClkMux I__5360 (
            .O(N__22219),
            .I(N__22008));
    ClkMux I__5359 (
            .O(N__22218),
            .I(N__22008));
    ClkMux I__5358 (
            .O(N__22217),
            .I(N__22008));
    ClkMux I__5357 (
            .O(N__22216),
            .I(N__22008));
    ClkMux I__5356 (
            .O(N__22215),
            .I(N__22008));
    ClkMux I__5355 (
            .O(N__22214),
            .I(N__22008));
    ClkMux I__5354 (
            .O(N__22213),
            .I(N__22008));
    ClkMux I__5353 (
            .O(N__22212),
            .I(N__22008));
    ClkMux I__5352 (
            .O(N__22211),
            .I(N__22008));
    ClkMux I__5351 (
            .O(N__22210),
            .I(N__22008));
    ClkMux I__5350 (
            .O(N__22209),
            .I(N__22008));
    ClkMux I__5349 (
            .O(N__22208),
            .I(N__22008));
    ClkMux I__5348 (
            .O(N__22207),
            .I(N__22008));
    ClkMux I__5347 (
            .O(N__22206),
            .I(N__22008));
    ClkMux I__5346 (
            .O(N__22205),
            .I(N__22008));
    ClkMux I__5345 (
            .O(N__22204),
            .I(N__22008));
    ClkMux I__5344 (
            .O(N__22203),
            .I(N__22008));
    ClkMux I__5343 (
            .O(N__22202),
            .I(N__22008));
    ClkMux I__5342 (
            .O(N__22201),
            .I(N__22008));
    ClkMux I__5341 (
            .O(N__22200),
            .I(N__22008));
    ClkMux I__5340 (
            .O(N__22199),
            .I(N__22008));
    ClkMux I__5339 (
            .O(N__22198),
            .I(N__22008));
    ClkMux I__5338 (
            .O(N__22197),
            .I(N__22008));
    ClkMux I__5337 (
            .O(N__22196),
            .I(N__22008));
    ClkMux I__5336 (
            .O(N__22195),
            .I(N__22008));
    ClkMux I__5335 (
            .O(N__22194),
            .I(N__22008));
    ClkMux I__5334 (
            .O(N__22193),
            .I(N__22008));
    ClkMux I__5333 (
            .O(N__22192),
            .I(N__22008));
    ClkMux I__5332 (
            .O(N__22191),
            .I(N__22008));
    ClkMux I__5331 (
            .O(N__22190),
            .I(N__22008));
    ClkMux I__5330 (
            .O(N__22189),
            .I(N__22008));
    ClkMux I__5329 (
            .O(N__22188),
            .I(N__22008));
    Glb2LocalMux I__5328 (
            .O(N__22185),
            .I(N__22008));
    GlobalMux I__5327 (
            .O(N__22008),
            .I(N__22005));
    gio2CtrlBuf I__5326 (
            .O(N__22005),
            .I(clk_g));
    CascadeMux I__5325 (
            .O(N__22002),
            .I(N__21999));
    InMux I__5324 (
            .O(N__21999),
            .I(N__21993));
    InMux I__5323 (
            .O(N__21998),
            .I(N__21993));
    LocalMux I__5322 (
            .O(N__21993),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__5321 (
            .O(N__21990),
            .I(N__21987));
    InMux I__5320 (
            .O(N__21987),
            .I(N__21981));
    InMux I__5319 (
            .O(N__21986),
            .I(N__21981));
    LocalMux I__5318 (
            .O(N__21981),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__5317 (
            .O(N__21978),
            .I(N__21974));
    InMux I__5316 (
            .O(N__21977),
            .I(N__21971));
    InMux I__5315 (
            .O(N__21974),
            .I(N__21968));
    LocalMux I__5314 (
            .O(N__21971),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__5313 (
            .O(N__21968),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__5312 (
            .O(N__21963),
            .I(N__21957));
    InMux I__5311 (
            .O(N__21962),
            .I(N__21957));
    LocalMux I__5310 (
            .O(N__21957),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__5309 (
            .O(N__21954),
            .I(N__21949));
    InMux I__5308 (
            .O(N__21953),
            .I(N__21944));
    InMux I__5307 (
            .O(N__21952),
            .I(N__21944));
    LocalMux I__5306 (
            .O(N__21949),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__5305 (
            .O(N__21944),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__5304 (
            .O(N__21939),
            .I(N__21934));
    InMux I__5303 (
            .O(N__21938),
            .I(N__21928));
    InMux I__5302 (
            .O(N__21937),
            .I(N__21928));
    InMux I__5301 (
            .O(N__21934),
            .I(N__21923));
    InMux I__5300 (
            .O(N__21933),
            .I(N__21923));
    LocalMux I__5299 (
            .O(N__21928),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__5298 (
            .O(N__21923),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__5297 (
            .O(N__21918),
            .I(N__21914));
    CascadeMux I__5296 (
            .O(N__21917),
            .I(N__21911));
    InMux I__5295 (
            .O(N__21914),
            .I(N__21906));
    InMux I__5294 (
            .O(N__21911),
            .I(N__21906));
    LocalMux I__5293 (
            .O(N__21906),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__5292 (
            .O(N__21903),
            .I(N__21900));
    LocalMux I__5291 (
            .O(N__21900),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    InMux I__5290 (
            .O(N__21897),
            .I(N__21887));
    InMux I__5289 (
            .O(N__21896),
            .I(N__21887));
    InMux I__5288 (
            .O(N__21895),
            .I(N__21887));
    InMux I__5287 (
            .O(N__21894),
            .I(N__21884));
    LocalMux I__5286 (
            .O(N__21887),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__5285 (
            .O(N__21884),
            .I(\buart.Z_tx.ser_clk ));
    InMux I__5284 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__5283 (
            .O(N__21876),
            .I(N__21873));
    Span4Mux_s3_v I__5282 (
            .O(N__21873),
            .I(N__21870));
    Span4Mux_h I__5281 (
            .O(N__21870),
            .I(N__21865));
    InMux I__5280 (
            .O(N__21869),
            .I(N__21860));
    InMux I__5279 (
            .O(N__21868),
            .I(N__21860));
    Odrv4 I__5278 (
            .O(N__21865),
            .I(L3_tx_data_2));
    LocalMux I__5277 (
            .O(N__21860),
            .I(L3_tx_data_2));
    InMux I__5276 (
            .O(N__21855),
            .I(N__21852));
    LocalMux I__5275 (
            .O(N__21852),
            .I(N__21849));
    Span4Mux_s0_v I__5274 (
            .O(N__21849),
            .I(N__21846));
    Span4Mux_h I__5273 (
            .O(N__21846),
            .I(N__21843));
    Odrv4 I__5272 (
            .O(N__21843),
            .I(\uu2.mem0.w_data_2 ));
    InMux I__5271 (
            .O(N__21840),
            .I(N__21833));
    InMux I__5270 (
            .O(N__21839),
            .I(N__21830));
    InMux I__5269 (
            .O(N__21838),
            .I(N__21825));
    InMux I__5268 (
            .O(N__21837),
            .I(N__21825));
    InMux I__5267 (
            .O(N__21836),
            .I(N__21822));
    LocalMux I__5266 (
            .O(N__21833),
            .I(N__21819));
    LocalMux I__5265 (
            .O(N__21830),
            .I(N__21814));
    LocalMux I__5264 (
            .O(N__21825),
            .I(N__21814));
    LocalMux I__5263 (
            .O(N__21822),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv12 I__5262 (
            .O(N__21819),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__5261 (
            .O(N__21814),
            .I(\uu2.w_addr_userZ0Z_2 ));
    InMux I__5260 (
            .O(N__21807),
            .I(N__21796));
    InMux I__5259 (
            .O(N__21806),
            .I(N__21796));
    InMux I__5258 (
            .O(N__21805),
            .I(N__21796));
    CascadeMux I__5257 (
            .O(N__21804),
            .I(N__21793));
    CascadeMux I__5256 (
            .O(N__21803),
            .I(N__21790));
    LocalMux I__5255 (
            .O(N__21796),
            .I(N__21782));
    InMux I__5254 (
            .O(N__21793),
            .I(N__21773));
    InMux I__5253 (
            .O(N__21790),
            .I(N__21773));
    InMux I__5252 (
            .O(N__21789),
            .I(N__21773));
    InMux I__5251 (
            .O(N__21788),
            .I(N__21773));
    CascadeMux I__5250 (
            .O(N__21787),
            .I(N__21769));
    InMux I__5249 (
            .O(N__21786),
            .I(N__21761));
    InMux I__5248 (
            .O(N__21785),
            .I(N__21758));
    Span4Mux_s2_v I__5247 (
            .O(N__21782),
            .I(N__21755));
    LocalMux I__5246 (
            .O(N__21773),
            .I(N__21752));
    InMux I__5245 (
            .O(N__21772),
            .I(N__21749));
    InMux I__5244 (
            .O(N__21769),
            .I(N__21735));
    InMux I__5243 (
            .O(N__21768),
            .I(N__21735));
    InMux I__5242 (
            .O(N__21767),
            .I(N__21735));
    InMux I__5241 (
            .O(N__21766),
            .I(N__21735));
    InMux I__5240 (
            .O(N__21765),
            .I(N__21735));
    InMux I__5239 (
            .O(N__21764),
            .I(N__21735));
    LocalMux I__5238 (
            .O(N__21761),
            .I(N__21730));
    LocalMux I__5237 (
            .O(N__21758),
            .I(N__21730));
    Span4Mux_h I__5236 (
            .O(N__21755),
            .I(N__21725));
    Span4Mux_s2_v I__5235 (
            .O(N__21752),
            .I(N__21725));
    LocalMux I__5234 (
            .O(N__21749),
            .I(N__21722));
    InMux I__5233 (
            .O(N__21748),
            .I(N__21719));
    LocalMux I__5232 (
            .O(N__21735),
            .I(N__21716));
    Span4Mux_s2_v I__5231 (
            .O(N__21730),
            .I(N__21713));
    Span4Mux_v I__5230 (
            .O(N__21725),
            .I(N__21708));
    Span4Mux_v I__5229 (
            .O(N__21722),
            .I(N__21708));
    LocalMux I__5228 (
            .O(N__21719),
            .I(N__21705));
    Span4Mux_s2_v I__5227 (
            .O(N__21716),
            .I(N__21700));
    Span4Mux_h I__5226 (
            .O(N__21713),
            .I(N__21700));
    Odrv4 I__5225 (
            .O(N__21708),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv12 I__5224 (
            .O(N__21705),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    Odrv4 I__5223 (
            .O(N__21700),
            .I(\uu2.un4_w_user_data_rdyZ0Z_0 ));
    InMux I__5222 (
            .O(N__21693),
            .I(N__21689));
    InMux I__5221 (
            .O(N__21692),
            .I(N__21685));
    LocalMux I__5220 (
            .O(N__21689),
            .I(N__21682));
    CascadeMux I__5219 (
            .O(N__21688),
            .I(N__21679));
    LocalMux I__5218 (
            .O(N__21685),
            .I(N__21667));
    Span4Mux_s2_v I__5217 (
            .O(N__21682),
            .I(N__21664));
    InMux I__5216 (
            .O(N__21679),
            .I(N__21655));
    InMux I__5215 (
            .O(N__21678),
            .I(N__21655));
    InMux I__5214 (
            .O(N__21677),
            .I(N__21655));
    InMux I__5213 (
            .O(N__21676),
            .I(N__21655));
    InMux I__5212 (
            .O(N__21675),
            .I(N__21650));
    InMux I__5211 (
            .O(N__21674),
            .I(N__21650));
    InMux I__5210 (
            .O(N__21673),
            .I(N__21641));
    InMux I__5209 (
            .O(N__21672),
            .I(N__21641));
    InMux I__5208 (
            .O(N__21671),
            .I(N__21641));
    InMux I__5207 (
            .O(N__21670),
            .I(N__21641));
    Span4Mux_h I__5206 (
            .O(N__21667),
            .I(N__21638));
    Odrv4 I__5205 (
            .O(N__21664),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5204 (
            .O(N__21655),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5203 (
            .O(N__21650),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__5202 (
            .O(N__21641),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv4 I__5201 (
            .O(N__21638),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    CascadeMux I__5200 (
            .O(N__21627),
            .I(N__21624));
    InMux I__5199 (
            .O(N__21624),
            .I(N__21621));
    LocalMux I__5198 (
            .O(N__21621),
            .I(N__21618));
    Span4Mux_h I__5197 (
            .O(N__21618),
            .I(N__21615));
    Span4Mux_h I__5196 (
            .O(N__21615),
            .I(N__21612));
    Odrv4 I__5195 (
            .O(N__21612),
            .I(\uu2.mem0.w_addr_2 ));
    InMux I__5194 (
            .O(N__21609),
            .I(N__21606));
    LocalMux I__5193 (
            .O(N__21606),
            .I(\buart.Z_tx.un1_bitcount_c2 ));
    InMux I__5192 (
            .O(N__21603),
            .I(N__21599));
    InMux I__5191 (
            .O(N__21602),
            .I(N__21596));
    LocalMux I__5190 (
            .O(N__21599),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__5189 (
            .O(N__21596),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    CascadeMux I__5188 (
            .O(N__21591),
            .I(\buart.Z_tx.uart_busy_0_0_cascade_ ));
    CascadeMux I__5187 (
            .O(N__21588),
            .I(N__21585));
    InMux I__5186 (
            .O(N__21585),
            .I(N__21577));
    InMux I__5185 (
            .O(N__21584),
            .I(N__21574));
    InMux I__5184 (
            .O(N__21583),
            .I(N__21565));
    InMux I__5183 (
            .O(N__21582),
            .I(N__21565));
    InMux I__5182 (
            .O(N__21581),
            .I(N__21565));
    InMux I__5181 (
            .O(N__21580),
            .I(N__21565));
    LocalMux I__5180 (
            .O(N__21577),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__5179 (
            .O(N__21574),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__5178 (
            .O(N__21565),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    InMux I__5177 (
            .O(N__21558),
            .I(N__21552));
    InMux I__5176 (
            .O(N__21557),
            .I(N__21545));
    InMux I__5175 (
            .O(N__21556),
            .I(N__21545));
    InMux I__5174 (
            .O(N__21555),
            .I(N__21545));
    LocalMux I__5173 (
            .O(N__21552),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__5172 (
            .O(N__21545),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__5171 (
            .O(N__21540),
            .I(N__21535));
    InMux I__5170 (
            .O(N__21539),
            .I(N__21530));
    InMux I__5169 (
            .O(N__21538),
            .I(N__21530));
    LocalMux I__5168 (
            .O(N__21535),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    LocalMux I__5167 (
            .O(N__21530),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__5166 (
            .O(N__21525),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    InMux I__5165 (
            .O(N__21522),
            .I(N__21513));
    InMux I__5164 (
            .O(N__21521),
            .I(N__21513));
    InMux I__5163 (
            .O(N__21520),
            .I(N__21506));
    InMux I__5162 (
            .O(N__21519),
            .I(N__21506));
    InMux I__5161 (
            .O(N__21518),
            .I(N__21506));
    LocalMux I__5160 (
            .O(N__21513),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__5159 (
            .O(N__21506),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    InMux I__5158 (
            .O(N__21501),
            .I(N__21498));
    LocalMux I__5157 (
            .O(N__21498),
            .I(\buart.Z_tx.un1_bitcount_c3 ));
    InMux I__5156 (
            .O(N__21495),
            .I(N__21487));
    InMux I__5155 (
            .O(N__21494),
            .I(N__21487));
    CascadeMux I__5154 (
            .O(N__21493),
            .I(N__21483));
    InMux I__5153 (
            .O(N__21492),
            .I(N__21477));
    LocalMux I__5152 (
            .O(N__21487),
            .I(N__21474));
    InMux I__5151 (
            .O(N__21486),
            .I(N__21469));
    InMux I__5150 (
            .O(N__21483),
            .I(N__21469));
    InMux I__5149 (
            .O(N__21482),
            .I(N__21462));
    InMux I__5148 (
            .O(N__21481),
            .I(N__21459));
    InMux I__5147 (
            .O(N__21480),
            .I(N__21456));
    LocalMux I__5146 (
            .O(N__21477),
            .I(N__21449));
    Span4Mux_h I__5145 (
            .O(N__21474),
            .I(N__21449));
    LocalMux I__5144 (
            .O(N__21469),
            .I(N__21449));
    InMux I__5143 (
            .O(N__21468),
            .I(N__21446));
    InMux I__5142 (
            .O(N__21467),
            .I(N__21439));
    InMux I__5141 (
            .O(N__21466),
            .I(N__21439));
    InMux I__5140 (
            .O(N__21465),
            .I(N__21439));
    LocalMux I__5139 (
            .O(N__21462),
            .I(N__21432));
    LocalMux I__5138 (
            .O(N__21459),
            .I(N__21429));
    LocalMux I__5137 (
            .O(N__21456),
            .I(N__21424));
    Span4Mux_v I__5136 (
            .O(N__21449),
            .I(N__21424));
    LocalMux I__5135 (
            .O(N__21446),
            .I(N__21419));
    LocalMux I__5134 (
            .O(N__21439),
            .I(N__21419));
    InMux I__5133 (
            .O(N__21438),
            .I(N__21410));
    InMux I__5132 (
            .O(N__21437),
            .I(N__21410));
    InMux I__5131 (
            .O(N__21436),
            .I(N__21410));
    InMux I__5130 (
            .O(N__21435),
            .I(N__21410));
    Span4Mux_h I__5129 (
            .O(N__21432),
            .I(N__21407));
    Odrv4 I__5128 (
            .O(N__21429),
            .I(N_63_mux));
    Odrv4 I__5127 (
            .O(N__21424),
            .I(N_63_mux));
    Odrv4 I__5126 (
            .O(N__21419),
            .I(N_63_mux));
    LocalMux I__5125 (
            .O(N__21410),
            .I(N_63_mux));
    Odrv4 I__5124 (
            .O(N__21407),
            .I(N_63_mux));
    CascadeMux I__5123 (
            .O(N__21396),
            .I(N__21392));
    InMux I__5122 (
            .O(N__21395),
            .I(N__21386));
    InMux I__5121 (
            .O(N__21392),
            .I(N__21383));
    CascadeMux I__5120 (
            .O(N__21391),
            .I(N__21380));
    InMux I__5119 (
            .O(N__21390),
            .I(N__21374));
    InMux I__5118 (
            .O(N__21389),
            .I(N__21371));
    LocalMux I__5117 (
            .O(N__21386),
            .I(N__21368));
    LocalMux I__5116 (
            .O(N__21383),
            .I(N__21365));
    InMux I__5115 (
            .O(N__21380),
            .I(N__21362));
    CascadeMux I__5114 (
            .O(N__21379),
            .I(N__21359));
    InMux I__5113 (
            .O(N__21378),
            .I(N__21356));
    InMux I__5112 (
            .O(N__21377),
            .I(N__21353));
    LocalMux I__5111 (
            .O(N__21374),
            .I(N__21349));
    LocalMux I__5110 (
            .O(N__21371),
            .I(N__21340));
    Span4Mux_s3_h I__5109 (
            .O(N__21368),
            .I(N__21340));
    Span4Mux_s3_h I__5108 (
            .O(N__21365),
            .I(N__21340));
    LocalMux I__5107 (
            .O(N__21362),
            .I(N__21340));
    InMux I__5106 (
            .O(N__21359),
            .I(N__21337));
    LocalMux I__5105 (
            .O(N__21356),
            .I(N__21330));
    LocalMux I__5104 (
            .O(N__21353),
            .I(N__21330));
    InMux I__5103 (
            .O(N__21352),
            .I(N__21327));
    Span4Mux_h I__5102 (
            .O(N__21349),
            .I(N__21322));
    Span4Mux_h I__5101 (
            .O(N__21340),
            .I(N__21322));
    LocalMux I__5100 (
            .O(N__21337),
            .I(N__21319));
    InMux I__5099 (
            .O(N__21336),
            .I(N__21316));
    CascadeMux I__5098 (
            .O(N__21335),
            .I(N__21309));
    Span4Mux_v I__5097 (
            .O(N__21330),
            .I(N__21303));
    LocalMux I__5096 (
            .O(N__21327),
            .I(N__21300));
    Span4Mux_v I__5095 (
            .O(N__21322),
            .I(N__21297));
    Span4Mux_v I__5094 (
            .O(N__21319),
            .I(N__21292));
    LocalMux I__5093 (
            .O(N__21316),
            .I(N__21292));
    InMux I__5092 (
            .O(N__21315),
            .I(N__21287));
    InMux I__5091 (
            .O(N__21314),
            .I(N__21287));
    InMux I__5090 (
            .O(N__21313),
            .I(N__21282));
    InMux I__5089 (
            .O(N__21312),
            .I(N__21282));
    InMux I__5088 (
            .O(N__21309),
            .I(N__21279));
    InMux I__5087 (
            .O(N__21308),
            .I(N__21274));
    InMux I__5086 (
            .O(N__21307),
            .I(N__21274));
    InMux I__5085 (
            .O(N__21306),
            .I(N__21271));
    Span4Mux_v I__5084 (
            .O(N__21303),
            .I(N__21268));
    Span4Mux_h I__5083 (
            .O(N__21300),
            .I(N__21263));
    Span4Mux_h I__5082 (
            .O(N__21297),
            .I(N__21263));
    Span4Mux_h I__5081 (
            .O(N__21292),
            .I(N__21258));
    LocalMux I__5080 (
            .O(N__21287),
            .I(N__21258));
    LocalMux I__5079 (
            .O(N__21282),
            .I(N__21255));
    LocalMux I__5078 (
            .O(N__21279),
            .I(N__21252));
    LocalMux I__5077 (
            .O(N__21274),
            .I(bu_rx_data_1));
    LocalMux I__5076 (
            .O(N__21271),
            .I(bu_rx_data_1));
    Odrv4 I__5075 (
            .O(N__21268),
            .I(bu_rx_data_1));
    Odrv4 I__5074 (
            .O(N__21263),
            .I(bu_rx_data_1));
    Odrv4 I__5073 (
            .O(N__21258),
            .I(bu_rx_data_1));
    Odrv4 I__5072 (
            .O(N__21255),
            .I(bu_rx_data_1));
    Odrv12 I__5071 (
            .O(N__21252),
            .I(bu_rx_data_1));
    InMux I__5070 (
            .O(N__21237),
            .I(N__21224));
    InMux I__5069 (
            .O(N__21236),
            .I(N__21224));
    InMux I__5068 (
            .O(N__21235),
            .I(N__21218));
    InMux I__5067 (
            .O(N__21234),
            .I(N__21218));
    InMux I__5066 (
            .O(N__21233),
            .I(N__21215));
    InMux I__5065 (
            .O(N__21232),
            .I(N__21207));
    InMux I__5064 (
            .O(N__21231),
            .I(N__21207));
    InMux I__5063 (
            .O(N__21230),
            .I(N__21202));
    InMux I__5062 (
            .O(N__21229),
            .I(N__21202));
    LocalMux I__5061 (
            .O(N__21224),
            .I(N__21199));
    InMux I__5060 (
            .O(N__21223),
            .I(N__21196));
    LocalMux I__5059 (
            .O(N__21218),
            .I(N__21193));
    LocalMux I__5058 (
            .O(N__21215),
            .I(N__21190));
    InMux I__5057 (
            .O(N__21214),
            .I(N__21187));
    CascadeMux I__5056 (
            .O(N__21213),
            .I(N__21184));
    InMux I__5055 (
            .O(N__21212),
            .I(N__21181));
    LocalMux I__5054 (
            .O(N__21207),
            .I(N__21176));
    LocalMux I__5053 (
            .O(N__21202),
            .I(N__21176));
    Span4Mux_v I__5052 (
            .O(N__21199),
            .I(N__21165));
    LocalMux I__5051 (
            .O(N__21196),
            .I(N__21165));
    Span4Mux_s3_h I__5050 (
            .O(N__21193),
            .I(N__21165));
    Span4Mux_s3_v I__5049 (
            .O(N__21190),
            .I(N__21165));
    LocalMux I__5048 (
            .O(N__21187),
            .I(N__21165));
    InMux I__5047 (
            .O(N__21184),
            .I(N__21162));
    LocalMux I__5046 (
            .O(N__21181),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5045 (
            .O(N__21176),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5044 (
            .O(N__21165),
            .I(bu_rx_data_3_rep2));
    LocalMux I__5043 (
            .O(N__21162),
            .I(bu_rx_data_3_rep2));
    InMux I__5042 (
            .O(N__21153),
            .I(N__21147));
    InMux I__5041 (
            .O(N__21152),
            .I(N__21147));
    LocalMux I__5040 (
            .O(N__21147),
            .I(N__21144));
    Odrv12 I__5039 (
            .O(N__21144),
            .I(N_14_0));
    InMux I__5038 (
            .O(N__21141),
            .I(N__21137));
    InMux I__5037 (
            .O(N__21140),
            .I(N__21131));
    LocalMux I__5036 (
            .O(N__21137),
            .I(N__21128));
    InMux I__5035 (
            .O(N__21136),
            .I(N__21125));
    CascadeMux I__5034 (
            .O(N__21135),
            .I(N__21122));
    InMux I__5033 (
            .O(N__21134),
            .I(N__21118));
    LocalMux I__5032 (
            .O(N__21131),
            .I(N__21108));
    Span4Mux_v I__5031 (
            .O(N__21128),
            .I(N__21108));
    LocalMux I__5030 (
            .O(N__21125),
            .I(N__21108));
    InMux I__5029 (
            .O(N__21122),
            .I(N__21105));
    InMux I__5028 (
            .O(N__21121),
            .I(N__21101));
    LocalMux I__5027 (
            .O(N__21118),
            .I(N__21098));
    InMux I__5026 (
            .O(N__21117),
            .I(N__21088));
    InMux I__5025 (
            .O(N__21116),
            .I(N__21085));
    InMux I__5024 (
            .O(N__21115),
            .I(N__21081));
    Span4Mux_h I__5023 (
            .O(N__21108),
            .I(N__21078));
    LocalMux I__5022 (
            .O(N__21105),
            .I(N__21075));
    InMux I__5021 (
            .O(N__21104),
            .I(N__21072));
    LocalMux I__5020 (
            .O(N__21101),
            .I(N__21069));
    Span4Mux_v I__5019 (
            .O(N__21098),
            .I(N__21066));
    InMux I__5018 (
            .O(N__21097),
            .I(N__21061));
    InMux I__5017 (
            .O(N__21096),
            .I(N__21061));
    InMux I__5016 (
            .O(N__21095),
            .I(N__21058));
    InMux I__5015 (
            .O(N__21094),
            .I(N__21055));
    InMux I__5014 (
            .O(N__21093),
            .I(N__21051));
    InMux I__5013 (
            .O(N__21092),
            .I(N__21048));
    InMux I__5012 (
            .O(N__21091),
            .I(N__21045));
    LocalMux I__5011 (
            .O(N__21088),
            .I(N__21039));
    LocalMux I__5010 (
            .O(N__21085),
            .I(N__21039));
    InMux I__5009 (
            .O(N__21084),
            .I(N__21036));
    LocalMux I__5008 (
            .O(N__21081),
            .I(N__21033));
    Span4Mux_v I__5007 (
            .O(N__21078),
            .I(N__21030));
    Span4Mux_v I__5006 (
            .O(N__21075),
            .I(N__21025));
    LocalMux I__5005 (
            .O(N__21072),
            .I(N__21025));
    Span4Mux_v I__5004 (
            .O(N__21069),
            .I(N__21022));
    Span4Mux_v I__5003 (
            .O(N__21066),
            .I(N__21015));
    LocalMux I__5002 (
            .O(N__21061),
            .I(N__21015));
    LocalMux I__5001 (
            .O(N__21058),
            .I(N__21015));
    LocalMux I__5000 (
            .O(N__21055),
            .I(N__21012));
    InMux I__4999 (
            .O(N__21054),
            .I(N__21009));
    LocalMux I__4998 (
            .O(N__21051),
            .I(N__21004));
    LocalMux I__4997 (
            .O(N__21048),
            .I(N__21004));
    LocalMux I__4996 (
            .O(N__21045),
            .I(N__21001));
    InMux I__4995 (
            .O(N__21044),
            .I(N__20998));
    Span12Mux_v I__4994 (
            .O(N__21039),
            .I(N__20995));
    LocalMux I__4993 (
            .O(N__21036),
            .I(N__20988));
    Span4Mux_h I__4992 (
            .O(N__21033),
            .I(N__20988));
    Span4Mux_v I__4991 (
            .O(N__21030),
            .I(N__20988));
    Span4Mux_h I__4990 (
            .O(N__21025),
            .I(N__20985));
    Span4Mux_v I__4989 (
            .O(N__21022),
            .I(N__20980));
    Span4Mux_h I__4988 (
            .O(N__21015),
            .I(N__20980));
    Span4Mux_v I__4987 (
            .O(N__21012),
            .I(N__20971));
    LocalMux I__4986 (
            .O(N__21009),
            .I(N__20971));
    Span4Mux_h I__4985 (
            .O(N__21004),
            .I(N__20971));
    Span4Mux_h I__4984 (
            .O(N__21001),
            .I(N__20971));
    LocalMux I__4983 (
            .O(N__20998),
            .I(bu_rx_data_3));
    Odrv12 I__4982 (
            .O(N__20995),
            .I(bu_rx_data_3));
    Odrv4 I__4981 (
            .O(N__20988),
            .I(bu_rx_data_3));
    Odrv4 I__4980 (
            .O(N__20985),
            .I(bu_rx_data_3));
    Odrv4 I__4979 (
            .O(N__20980),
            .I(bu_rx_data_3));
    Odrv4 I__4978 (
            .O(N__20971),
            .I(bu_rx_data_3));
    InMux I__4977 (
            .O(N__20958),
            .I(N__20953));
    InMux I__4976 (
            .O(N__20957),
            .I(N__20950));
    InMux I__4975 (
            .O(N__20956),
            .I(N__20947));
    LocalMux I__4974 (
            .O(N__20953),
            .I(N__20940));
    LocalMux I__4973 (
            .O(N__20950),
            .I(N__20940));
    LocalMux I__4972 (
            .O(N__20947),
            .I(N__20937));
    InMux I__4971 (
            .O(N__20946),
            .I(N__20934));
    InMux I__4970 (
            .O(N__20945),
            .I(N__20929));
    Span4Mux_v I__4969 (
            .O(N__20940),
            .I(N__20919));
    Span4Mux_h I__4968 (
            .O(N__20937),
            .I(N__20919));
    LocalMux I__4967 (
            .O(N__20934),
            .I(N__20919));
    InMux I__4966 (
            .O(N__20933),
            .I(N__20916));
    InMux I__4965 (
            .O(N__20932),
            .I(N__20913));
    LocalMux I__4964 (
            .O(N__20929),
            .I(N__20910));
    CascadeMux I__4963 (
            .O(N__20928),
            .I(N__20905));
    CascadeMux I__4962 (
            .O(N__20927),
            .I(N__20901));
    InMux I__4961 (
            .O(N__20926),
            .I(N__20897));
    Span4Mux_h I__4960 (
            .O(N__20919),
            .I(N__20894));
    LocalMux I__4959 (
            .O(N__20916),
            .I(N__20889));
    LocalMux I__4958 (
            .O(N__20913),
            .I(N__20889));
    Span4Mux_v I__4957 (
            .O(N__20910),
            .I(N__20886));
    InMux I__4956 (
            .O(N__20909),
            .I(N__20883));
    InMux I__4955 (
            .O(N__20908),
            .I(N__20880));
    InMux I__4954 (
            .O(N__20905),
            .I(N__20875));
    InMux I__4953 (
            .O(N__20904),
            .I(N__20875));
    InMux I__4952 (
            .O(N__20901),
            .I(N__20871));
    InMux I__4951 (
            .O(N__20900),
            .I(N__20868));
    LocalMux I__4950 (
            .O(N__20897),
            .I(N__20865));
    Span4Mux_v I__4949 (
            .O(N__20894),
            .I(N__20862));
    Span4Mux_v I__4948 (
            .O(N__20889),
            .I(N__20858));
    Span4Mux_v I__4947 (
            .O(N__20886),
            .I(N__20849));
    LocalMux I__4946 (
            .O(N__20883),
            .I(N__20849));
    LocalMux I__4945 (
            .O(N__20880),
            .I(N__20849));
    LocalMux I__4944 (
            .O(N__20875),
            .I(N__20849));
    InMux I__4943 (
            .O(N__20874),
            .I(N__20843));
    LocalMux I__4942 (
            .O(N__20871),
            .I(N__20840));
    LocalMux I__4941 (
            .O(N__20868),
            .I(N__20837));
    Span12Mux_s8_v I__4940 (
            .O(N__20865),
            .I(N__20834));
    Span4Mux_v I__4939 (
            .O(N__20862),
            .I(N__20831));
    InMux I__4938 (
            .O(N__20861),
            .I(N__20828));
    Span4Mux_v I__4937 (
            .O(N__20858),
            .I(N__20823));
    Span4Mux_h I__4936 (
            .O(N__20849),
            .I(N__20823));
    InMux I__4935 (
            .O(N__20848),
            .I(N__20816));
    InMux I__4934 (
            .O(N__20847),
            .I(N__20816));
    InMux I__4933 (
            .O(N__20846),
            .I(N__20816));
    LocalMux I__4932 (
            .O(N__20843),
            .I(N__20811));
    Span4Mux_h I__4931 (
            .O(N__20840),
            .I(N__20811));
    Odrv12 I__4930 (
            .O(N__20837),
            .I(bu_rx_data_2));
    Odrv12 I__4929 (
            .O(N__20834),
            .I(bu_rx_data_2));
    Odrv4 I__4928 (
            .O(N__20831),
            .I(bu_rx_data_2));
    LocalMux I__4927 (
            .O(N__20828),
            .I(bu_rx_data_2));
    Odrv4 I__4926 (
            .O(N__20823),
            .I(bu_rx_data_2));
    LocalMux I__4925 (
            .O(N__20816),
            .I(bu_rx_data_2));
    Odrv4 I__4924 (
            .O(N__20811),
            .I(bu_rx_data_2));
    CEMux I__4923 (
            .O(N__20796),
            .I(N__20772));
    CEMux I__4922 (
            .O(N__20795),
            .I(N__20772));
    CEMux I__4921 (
            .O(N__20794),
            .I(N__20772));
    CEMux I__4920 (
            .O(N__20793),
            .I(N__20772));
    CEMux I__4919 (
            .O(N__20792),
            .I(N__20772));
    CEMux I__4918 (
            .O(N__20791),
            .I(N__20772));
    CEMux I__4917 (
            .O(N__20790),
            .I(N__20772));
    CEMux I__4916 (
            .O(N__20789),
            .I(N__20772));
    GlobalMux I__4915 (
            .O(N__20772),
            .I(N__20769));
    gio2CtrlBuf I__4914 (
            .O(N__20769),
            .I(\buart.Z_rx.sample_g ));
    CascadeMux I__4913 (
            .O(N__20766),
            .I(N__20758));
    CascadeMux I__4912 (
            .O(N__20765),
            .I(N__20751));
    InMux I__4911 (
            .O(N__20764),
            .I(N__20743));
    InMux I__4910 (
            .O(N__20763),
            .I(N__20740));
    InMux I__4909 (
            .O(N__20762),
            .I(N__20737));
    InMux I__4908 (
            .O(N__20761),
            .I(N__20734));
    InMux I__4907 (
            .O(N__20758),
            .I(N__20731));
    InMux I__4906 (
            .O(N__20757),
            .I(N__20728));
    InMux I__4905 (
            .O(N__20756),
            .I(N__20723));
    InMux I__4904 (
            .O(N__20755),
            .I(N__20723));
    InMux I__4903 (
            .O(N__20754),
            .I(N__20720));
    InMux I__4902 (
            .O(N__20751),
            .I(N__20717));
    InMux I__4901 (
            .O(N__20750),
            .I(N__20714));
    InMux I__4900 (
            .O(N__20749),
            .I(N__20711));
    InMux I__4899 (
            .O(N__20748),
            .I(N__20708));
    InMux I__4898 (
            .O(N__20747),
            .I(N__20703));
    InMux I__4897 (
            .O(N__20746),
            .I(N__20703));
    LocalMux I__4896 (
            .O(N__20743),
            .I(N__20700));
    LocalMux I__4895 (
            .O(N__20740),
            .I(N__20655));
    LocalMux I__4894 (
            .O(N__20737),
            .I(N__20652));
    LocalMux I__4893 (
            .O(N__20734),
            .I(N__20649));
    LocalMux I__4892 (
            .O(N__20731),
            .I(N__20646));
    LocalMux I__4891 (
            .O(N__20728),
            .I(N__20643));
    LocalMux I__4890 (
            .O(N__20723),
            .I(N__20640));
    LocalMux I__4889 (
            .O(N__20720),
            .I(N__20637));
    LocalMux I__4888 (
            .O(N__20717),
            .I(N__20634));
    LocalMux I__4887 (
            .O(N__20714),
            .I(N__20631));
    LocalMux I__4886 (
            .O(N__20711),
            .I(N__20614));
    LocalMux I__4885 (
            .O(N__20708),
            .I(N__20611));
    LocalMux I__4884 (
            .O(N__20703),
            .I(N__20608));
    Glb2LocalMux I__4883 (
            .O(N__20700),
            .I(N__20469));
    SRMux I__4882 (
            .O(N__20699),
            .I(N__20469));
    SRMux I__4881 (
            .O(N__20698),
            .I(N__20469));
    SRMux I__4880 (
            .O(N__20697),
            .I(N__20469));
    SRMux I__4879 (
            .O(N__20696),
            .I(N__20469));
    SRMux I__4878 (
            .O(N__20695),
            .I(N__20469));
    SRMux I__4877 (
            .O(N__20694),
            .I(N__20469));
    SRMux I__4876 (
            .O(N__20693),
            .I(N__20469));
    SRMux I__4875 (
            .O(N__20692),
            .I(N__20469));
    SRMux I__4874 (
            .O(N__20691),
            .I(N__20469));
    SRMux I__4873 (
            .O(N__20690),
            .I(N__20469));
    SRMux I__4872 (
            .O(N__20689),
            .I(N__20469));
    SRMux I__4871 (
            .O(N__20688),
            .I(N__20469));
    SRMux I__4870 (
            .O(N__20687),
            .I(N__20469));
    SRMux I__4869 (
            .O(N__20686),
            .I(N__20469));
    SRMux I__4868 (
            .O(N__20685),
            .I(N__20469));
    SRMux I__4867 (
            .O(N__20684),
            .I(N__20469));
    SRMux I__4866 (
            .O(N__20683),
            .I(N__20469));
    SRMux I__4865 (
            .O(N__20682),
            .I(N__20469));
    SRMux I__4864 (
            .O(N__20681),
            .I(N__20469));
    SRMux I__4863 (
            .O(N__20680),
            .I(N__20469));
    SRMux I__4862 (
            .O(N__20679),
            .I(N__20469));
    SRMux I__4861 (
            .O(N__20678),
            .I(N__20469));
    SRMux I__4860 (
            .O(N__20677),
            .I(N__20469));
    SRMux I__4859 (
            .O(N__20676),
            .I(N__20469));
    SRMux I__4858 (
            .O(N__20675),
            .I(N__20469));
    SRMux I__4857 (
            .O(N__20674),
            .I(N__20469));
    SRMux I__4856 (
            .O(N__20673),
            .I(N__20469));
    SRMux I__4855 (
            .O(N__20672),
            .I(N__20469));
    SRMux I__4854 (
            .O(N__20671),
            .I(N__20469));
    SRMux I__4853 (
            .O(N__20670),
            .I(N__20469));
    SRMux I__4852 (
            .O(N__20669),
            .I(N__20469));
    SRMux I__4851 (
            .O(N__20668),
            .I(N__20469));
    SRMux I__4850 (
            .O(N__20667),
            .I(N__20469));
    SRMux I__4849 (
            .O(N__20666),
            .I(N__20469));
    SRMux I__4848 (
            .O(N__20665),
            .I(N__20469));
    SRMux I__4847 (
            .O(N__20664),
            .I(N__20469));
    SRMux I__4846 (
            .O(N__20663),
            .I(N__20469));
    SRMux I__4845 (
            .O(N__20662),
            .I(N__20469));
    SRMux I__4844 (
            .O(N__20661),
            .I(N__20469));
    SRMux I__4843 (
            .O(N__20660),
            .I(N__20469));
    SRMux I__4842 (
            .O(N__20659),
            .I(N__20469));
    SRMux I__4841 (
            .O(N__20658),
            .I(N__20469));
    Glb2LocalMux I__4840 (
            .O(N__20655),
            .I(N__20469));
    Glb2LocalMux I__4839 (
            .O(N__20652),
            .I(N__20469));
    Glb2LocalMux I__4838 (
            .O(N__20649),
            .I(N__20469));
    Glb2LocalMux I__4837 (
            .O(N__20646),
            .I(N__20469));
    Glb2LocalMux I__4836 (
            .O(N__20643),
            .I(N__20469));
    Glb2LocalMux I__4835 (
            .O(N__20640),
            .I(N__20469));
    Glb2LocalMux I__4834 (
            .O(N__20637),
            .I(N__20469));
    Glb2LocalMux I__4833 (
            .O(N__20634),
            .I(N__20469));
    Glb2LocalMux I__4832 (
            .O(N__20631),
            .I(N__20469));
    SRMux I__4831 (
            .O(N__20630),
            .I(N__20469));
    SRMux I__4830 (
            .O(N__20629),
            .I(N__20469));
    SRMux I__4829 (
            .O(N__20628),
            .I(N__20469));
    SRMux I__4828 (
            .O(N__20627),
            .I(N__20469));
    SRMux I__4827 (
            .O(N__20626),
            .I(N__20469));
    SRMux I__4826 (
            .O(N__20625),
            .I(N__20469));
    SRMux I__4825 (
            .O(N__20624),
            .I(N__20469));
    SRMux I__4824 (
            .O(N__20623),
            .I(N__20469));
    SRMux I__4823 (
            .O(N__20622),
            .I(N__20469));
    SRMux I__4822 (
            .O(N__20621),
            .I(N__20469));
    SRMux I__4821 (
            .O(N__20620),
            .I(N__20469));
    SRMux I__4820 (
            .O(N__20619),
            .I(N__20469));
    SRMux I__4819 (
            .O(N__20618),
            .I(N__20469));
    SRMux I__4818 (
            .O(N__20617),
            .I(N__20469));
    Glb2LocalMux I__4817 (
            .O(N__20614),
            .I(N__20469));
    Glb2LocalMux I__4816 (
            .O(N__20611),
            .I(N__20469));
    Glb2LocalMux I__4815 (
            .O(N__20608),
            .I(N__20469));
    GlobalMux I__4814 (
            .O(N__20469),
            .I(N__20466));
    gio2CtrlBuf I__4813 (
            .O(N__20466),
            .I(rst_g));
    CascadeMux I__4812 (
            .O(N__20463),
            .I(N__20458));
    CascadeMux I__4811 (
            .O(N__20462),
            .I(N__20454));
    InMux I__4810 (
            .O(N__20461),
            .I(N__20446));
    InMux I__4809 (
            .O(N__20458),
            .I(N__20446));
    InMux I__4808 (
            .O(N__20457),
            .I(N__20439));
    InMux I__4807 (
            .O(N__20454),
            .I(N__20439));
    InMux I__4806 (
            .O(N__20453),
            .I(N__20439));
    InMux I__4805 (
            .O(N__20452),
            .I(N__20433));
    InMux I__4804 (
            .O(N__20451),
            .I(N__20433));
    LocalMux I__4803 (
            .O(N__20446),
            .I(N__20428));
    LocalMux I__4802 (
            .O(N__20439),
            .I(N__20428));
    CascadeMux I__4801 (
            .O(N__20438),
            .I(N__20425));
    LocalMux I__4800 (
            .O(N__20433),
            .I(N__20414));
    Span4Mux_s2_v I__4799 (
            .O(N__20428),
            .I(N__20411));
    InMux I__4798 (
            .O(N__20425),
            .I(N__20408));
    InMux I__4797 (
            .O(N__20424),
            .I(N__20391));
    InMux I__4796 (
            .O(N__20423),
            .I(N__20391));
    InMux I__4795 (
            .O(N__20422),
            .I(N__20391));
    InMux I__4794 (
            .O(N__20421),
            .I(N__20391));
    InMux I__4793 (
            .O(N__20420),
            .I(N__20391));
    InMux I__4792 (
            .O(N__20419),
            .I(N__20391));
    InMux I__4791 (
            .O(N__20418),
            .I(N__20391));
    InMux I__4790 (
            .O(N__20417),
            .I(N__20391));
    Span4Mux_h I__4789 (
            .O(N__20414),
            .I(N__20388));
    Sp12to4 I__4788 (
            .O(N__20411),
            .I(N__20385));
    LocalMux I__4787 (
            .O(N__20408),
            .I(vbuf_tx_data_rdy));
    LocalMux I__4786 (
            .O(N__20391),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__4785 (
            .O(N__20388),
            .I(vbuf_tx_data_rdy));
    Odrv12 I__4784 (
            .O(N__20385),
            .I(vbuf_tx_data_rdy));
    CEMux I__4783 (
            .O(N__20376),
            .I(N__20373));
    LocalMux I__4782 (
            .O(N__20373),
            .I(N__20369));
    CEMux I__4781 (
            .O(N__20372),
            .I(N__20366));
    Span4Mux_s2_v I__4780 (
            .O(N__20369),
            .I(N__20363));
    LocalMux I__4779 (
            .O(N__20366),
            .I(N__20360));
    Span4Mux_h I__4778 (
            .O(N__20363),
            .I(N__20357));
    Span4Mux_h I__4777 (
            .O(N__20360),
            .I(N__20354));
    Span4Mux_h I__4776 (
            .O(N__20357),
            .I(N__20351));
    Span4Mux_s0_v I__4775 (
            .O(N__20354),
            .I(N__20348));
    Odrv4 I__4774 (
            .O(N__20351),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__4773 (
            .O(N__20348),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    InMux I__4772 (
            .O(N__20343),
            .I(N__20337));
    CascadeMux I__4771 (
            .O(N__20342),
            .I(N__20334));
    CascadeMux I__4770 (
            .O(N__20341),
            .I(N__20329));
    InMux I__4769 (
            .O(N__20340),
            .I(N__20326));
    LocalMux I__4768 (
            .O(N__20337),
            .I(N__20323));
    InMux I__4767 (
            .O(N__20334),
            .I(N__20318));
    InMux I__4766 (
            .O(N__20333),
            .I(N__20318));
    InMux I__4765 (
            .O(N__20332),
            .I(N__20313));
    InMux I__4764 (
            .O(N__20329),
            .I(N__20313));
    LocalMux I__4763 (
            .O(N__20326),
            .I(N__20306));
    Span4Mux_s2_h I__4762 (
            .O(N__20323),
            .I(N__20306));
    LocalMux I__4761 (
            .O(N__20318),
            .I(N__20306));
    LocalMux I__4760 (
            .O(N__20313),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__4759 (
            .O(N__20306),
            .I(\uu2.w_addr_userZ0Z_1 ));
    InMux I__4758 (
            .O(N__20301),
            .I(N__20298));
    LocalMux I__4757 (
            .O(N__20298),
            .I(N__20291));
    InMux I__4756 (
            .O(N__20297),
            .I(N__20282));
    InMux I__4755 (
            .O(N__20296),
            .I(N__20282));
    InMux I__4754 (
            .O(N__20295),
            .I(N__20282));
    InMux I__4753 (
            .O(N__20294),
            .I(N__20282));
    Span4Mux_s1_v I__4752 (
            .O(N__20291),
            .I(N__20279));
    LocalMux I__4751 (
            .O(N__20282),
            .I(N__20270));
    Span4Mux_h I__4750 (
            .O(N__20279),
            .I(N__20267));
    InMux I__4749 (
            .O(N__20278),
            .I(N__20256));
    InMux I__4748 (
            .O(N__20277),
            .I(N__20256));
    InMux I__4747 (
            .O(N__20276),
            .I(N__20256));
    InMux I__4746 (
            .O(N__20275),
            .I(N__20256));
    InMux I__4745 (
            .O(N__20274),
            .I(N__20256));
    InMux I__4744 (
            .O(N__20273),
            .I(N__20253));
    Span4Mux_h I__4743 (
            .O(N__20270),
            .I(N__20250));
    Odrv4 I__4742 (
            .O(N__20267),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__4741 (
            .O(N__20256),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__4740 (
            .O(N__20253),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__4739 (
            .O(N__20250),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__4738 (
            .O(N__20241),
            .I(N__20238));
    InMux I__4737 (
            .O(N__20238),
            .I(N__20235));
    LocalMux I__4736 (
            .O(N__20235),
            .I(N__20232));
    Odrv12 I__4735 (
            .O(N__20232),
            .I(\uu2.mem0.w_addr_1 ));
    InMux I__4734 (
            .O(N__20229),
            .I(N__20225));
    InMux I__4733 (
            .O(N__20228),
            .I(N__20222));
    LocalMux I__4732 (
            .O(N__20225),
            .I(N__20219));
    LocalMux I__4731 (
            .O(N__20222),
            .I(\Lab_UT.dictrl.N_8_0 ));
    Odrv4 I__4730 (
            .O(N__20219),
            .I(\Lab_UT.dictrl.N_8_0 ));
    InMux I__4729 (
            .O(N__20214),
            .I(N__20211));
    LocalMux I__4728 (
            .O(N__20211),
            .I(N__20208));
    Odrv4 I__4727 (
            .O(N__20208),
            .I(\Lab_UT.dictrl.i8_mux ));
    InMux I__4726 (
            .O(N__20205),
            .I(N__20200));
    CascadeMux I__4725 (
            .O(N__20204),
            .I(N__20197));
    InMux I__4724 (
            .O(N__20203),
            .I(N__20193));
    LocalMux I__4723 (
            .O(N__20200),
            .I(N__20189));
    InMux I__4722 (
            .O(N__20197),
            .I(N__20184));
    InMux I__4721 (
            .O(N__20196),
            .I(N__20184));
    LocalMux I__4720 (
            .O(N__20193),
            .I(N__20180));
    InMux I__4719 (
            .O(N__20192),
            .I(N__20177));
    Span4Mux_s3_v I__4718 (
            .O(N__20189),
            .I(N__20174));
    LocalMux I__4717 (
            .O(N__20184),
            .I(N__20171));
    InMux I__4716 (
            .O(N__20183),
            .I(N__20168));
    Odrv4 I__4715 (
            .O(N__20180),
            .I(bu_rx_data_fast_2));
    LocalMux I__4714 (
            .O(N__20177),
            .I(bu_rx_data_fast_2));
    Odrv4 I__4713 (
            .O(N__20174),
            .I(bu_rx_data_fast_2));
    Odrv12 I__4712 (
            .O(N__20171),
            .I(bu_rx_data_fast_2));
    LocalMux I__4711 (
            .O(N__20168),
            .I(bu_rx_data_fast_2));
    CascadeMux I__4710 (
            .O(N__20157),
            .I(N__20153));
    CascadeMux I__4709 (
            .O(N__20156),
            .I(N__20149));
    InMux I__4708 (
            .O(N__20153),
            .I(N__20144));
    InMux I__4707 (
            .O(N__20152),
            .I(N__20144));
    InMux I__4706 (
            .O(N__20149),
            .I(N__20141));
    LocalMux I__4705 (
            .O(N__20144),
            .I(N__20136));
    LocalMux I__4704 (
            .O(N__20141),
            .I(N__20132));
    CascadeMux I__4703 (
            .O(N__20140),
            .I(N__20129));
    InMux I__4702 (
            .O(N__20139),
            .I(N__20122));
    Span4Mux_v I__4701 (
            .O(N__20136),
            .I(N__20119));
    InMux I__4700 (
            .O(N__20135),
            .I(N__20116));
    Span4Mux_h I__4699 (
            .O(N__20132),
            .I(N__20113));
    InMux I__4698 (
            .O(N__20129),
            .I(N__20110));
    InMux I__4697 (
            .O(N__20128),
            .I(N__20107));
    InMux I__4696 (
            .O(N__20127),
            .I(N__20104));
    InMux I__4695 (
            .O(N__20126),
            .I(N__20099));
    InMux I__4694 (
            .O(N__20125),
            .I(N__20099));
    LocalMux I__4693 (
            .O(N__20122),
            .I(N__20096));
    Span4Mux_s3_v I__4692 (
            .O(N__20119),
            .I(N__20079));
    LocalMux I__4691 (
            .O(N__20116),
            .I(N__20079));
    Span4Mux_s3_v I__4690 (
            .O(N__20113),
            .I(N__20079));
    LocalMux I__4689 (
            .O(N__20110),
            .I(N__20079));
    LocalMux I__4688 (
            .O(N__20107),
            .I(N__20079));
    LocalMux I__4687 (
            .O(N__20104),
            .I(N__20079));
    LocalMux I__4686 (
            .O(N__20099),
            .I(N__20079));
    Span4Mux_h I__4685 (
            .O(N__20096),
            .I(N__20076));
    InMux I__4684 (
            .O(N__20095),
            .I(N__20071));
    InMux I__4683 (
            .O(N__20094),
            .I(N__20071));
    Span4Mux_v I__4682 (
            .O(N__20079),
            .I(N__20068));
    Odrv4 I__4681 (
            .O(N__20076),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    LocalMux I__4680 (
            .O(N__20071),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    Odrv4 I__4679 (
            .O(N__20068),
            .I(\Lab_UT.dictrl.state_0_rep1 ));
    CascadeMux I__4678 (
            .O(N__20061),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_ ));
    InMux I__4677 (
            .O(N__20058),
            .I(N__20055));
    LocalMux I__4676 (
            .O(N__20055),
            .I(\Lab_UT.dictrl.N_3 ));
    InMux I__4675 (
            .O(N__20052),
            .I(N__20047));
    InMux I__4674 (
            .O(N__20051),
            .I(N__20043));
    InMux I__4673 (
            .O(N__20050),
            .I(N__20040));
    LocalMux I__4672 (
            .O(N__20047),
            .I(N__20037));
    InMux I__4671 (
            .O(N__20046),
            .I(N__20034));
    LocalMux I__4670 (
            .O(N__20043),
            .I(N__20027));
    LocalMux I__4669 (
            .O(N__20040),
            .I(N__20020));
    Span4Mux_h I__4668 (
            .O(N__20037),
            .I(N__20020));
    LocalMux I__4667 (
            .O(N__20034),
            .I(N__20020));
    InMux I__4666 (
            .O(N__20033),
            .I(N__20017));
    InMux I__4665 (
            .O(N__20032),
            .I(N__20014));
    InMux I__4664 (
            .O(N__20031),
            .I(N__20011));
    InMux I__4663 (
            .O(N__20030),
            .I(N__20008));
    Span4Mux_v I__4662 (
            .O(N__20027),
            .I(N__20003));
    Span4Mux_v I__4661 (
            .O(N__20020),
            .I(N__20000));
    LocalMux I__4660 (
            .O(N__20017),
            .I(N__19991));
    LocalMux I__4659 (
            .O(N__20014),
            .I(N__19991));
    LocalMux I__4658 (
            .O(N__20011),
            .I(N__19991));
    LocalMux I__4657 (
            .O(N__20008),
            .I(N__19991));
    InMux I__4656 (
            .O(N__20007),
            .I(N__19986));
    InMux I__4655 (
            .O(N__20006),
            .I(N__19982));
    Span4Mux_v I__4654 (
            .O(N__20003),
            .I(N__19977));
    Span4Mux_v I__4653 (
            .O(N__20000),
            .I(N__19977));
    Span4Mux_v I__4652 (
            .O(N__19991),
            .I(N__19974));
    InMux I__4651 (
            .O(N__19990),
            .I(N__19971));
    InMux I__4650 (
            .O(N__19989),
            .I(N__19968));
    LocalMux I__4649 (
            .O(N__19986),
            .I(N__19965));
    InMux I__4648 (
            .O(N__19985),
            .I(N__19962));
    LocalMux I__4647 (
            .O(N__19982),
            .I(N__19959));
    Odrv4 I__4646 (
            .O(N__19977),
            .I(bu_rx_data_0));
    Odrv4 I__4645 (
            .O(N__19974),
            .I(bu_rx_data_0));
    LocalMux I__4644 (
            .O(N__19971),
            .I(bu_rx_data_0));
    LocalMux I__4643 (
            .O(N__19968),
            .I(bu_rx_data_0));
    Odrv12 I__4642 (
            .O(N__19965),
            .I(bu_rx_data_0));
    LocalMux I__4641 (
            .O(N__19962),
            .I(bu_rx_data_0));
    Odrv4 I__4640 (
            .O(N__19959),
            .I(bu_rx_data_0));
    CascadeMux I__4639 (
            .O(N__19944),
            .I(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_ ));
    InMux I__4638 (
            .O(N__19941),
            .I(N__19938));
    LocalMux I__4637 (
            .O(N__19938),
            .I(\Lab_UT.dictrl.next_state_RNO_5Z0Z_0 ));
    InMux I__4636 (
            .O(N__19935),
            .I(N__19932));
    LocalMux I__4635 (
            .O(N__19932),
            .I(\Lab_UT.dictrl.i9_mux ));
    CascadeMux I__4634 (
            .O(N__19929),
            .I(N__19924));
    InMux I__4633 (
            .O(N__19928),
            .I(N__19911));
    InMux I__4632 (
            .O(N__19927),
            .I(N__19911));
    InMux I__4631 (
            .O(N__19924),
            .I(N__19906));
    InMux I__4630 (
            .O(N__19923),
            .I(N__19903));
    InMux I__4629 (
            .O(N__19922),
            .I(N__19900));
    InMux I__4628 (
            .O(N__19921),
            .I(N__19897));
    InMux I__4627 (
            .O(N__19920),
            .I(N__19894));
    InMux I__4626 (
            .O(N__19919),
            .I(N__19889));
    InMux I__4625 (
            .O(N__19918),
            .I(N__19889));
    InMux I__4624 (
            .O(N__19917),
            .I(N__19877));
    InMux I__4623 (
            .O(N__19916),
            .I(N__19877));
    LocalMux I__4622 (
            .O(N__19911),
            .I(N__19874));
    InMux I__4621 (
            .O(N__19910),
            .I(N__19869));
    InMux I__4620 (
            .O(N__19909),
            .I(N__19869));
    LocalMux I__4619 (
            .O(N__19906),
            .I(N__19866));
    LocalMux I__4618 (
            .O(N__19903),
            .I(N__19860));
    LocalMux I__4617 (
            .O(N__19900),
            .I(N__19857));
    LocalMux I__4616 (
            .O(N__19897),
            .I(N__19850));
    LocalMux I__4615 (
            .O(N__19894),
            .I(N__19850));
    LocalMux I__4614 (
            .O(N__19889),
            .I(N__19850));
    InMux I__4613 (
            .O(N__19888),
            .I(N__19845));
    InMux I__4612 (
            .O(N__19887),
            .I(N__19845));
    InMux I__4611 (
            .O(N__19886),
            .I(N__19842));
    InMux I__4610 (
            .O(N__19885),
            .I(N__19837));
    InMux I__4609 (
            .O(N__19884),
            .I(N__19837));
    InMux I__4608 (
            .O(N__19883),
            .I(N__19832));
    InMux I__4607 (
            .O(N__19882),
            .I(N__19832));
    LocalMux I__4606 (
            .O(N__19877),
            .I(N__19822));
    Span4Mux_v I__4605 (
            .O(N__19874),
            .I(N__19822));
    LocalMux I__4604 (
            .O(N__19869),
            .I(N__19822));
    Span4Mux_h I__4603 (
            .O(N__19866),
            .I(N__19822));
    InMux I__4602 (
            .O(N__19865),
            .I(N__19819));
    InMux I__4601 (
            .O(N__19864),
            .I(N__19814));
    InMux I__4600 (
            .O(N__19863),
            .I(N__19814));
    Span4Mux_h I__4599 (
            .O(N__19860),
            .I(N__19803));
    Span4Mux_v I__4598 (
            .O(N__19857),
            .I(N__19803));
    Span4Mux_v I__4597 (
            .O(N__19850),
            .I(N__19803));
    LocalMux I__4596 (
            .O(N__19845),
            .I(N__19803));
    LocalMux I__4595 (
            .O(N__19842),
            .I(N__19803));
    LocalMux I__4594 (
            .O(N__19837),
            .I(N__19800));
    LocalMux I__4593 (
            .O(N__19832),
            .I(N__19797));
    InMux I__4592 (
            .O(N__19831),
            .I(N__19794));
    Odrv4 I__4591 (
            .O(N__19822),
            .I(Lab_UT_dictrl_state_1));
    LocalMux I__4590 (
            .O(N__19819),
            .I(Lab_UT_dictrl_state_1));
    LocalMux I__4589 (
            .O(N__19814),
            .I(Lab_UT_dictrl_state_1));
    Odrv4 I__4588 (
            .O(N__19803),
            .I(Lab_UT_dictrl_state_1));
    Odrv12 I__4587 (
            .O(N__19800),
            .I(Lab_UT_dictrl_state_1));
    Odrv4 I__4586 (
            .O(N__19797),
            .I(Lab_UT_dictrl_state_1));
    LocalMux I__4585 (
            .O(N__19794),
            .I(Lab_UT_dictrl_state_1));
    CascadeMux I__4584 (
            .O(N__19779),
            .I(N__19770));
    InMux I__4583 (
            .O(N__19778),
            .I(N__19763));
    InMux I__4582 (
            .O(N__19777),
            .I(N__19763));
    InMux I__4581 (
            .O(N__19776),
            .I(N__19763));
    CascadeMux I__4580 (
            .O(N__19775),
            .I(N__19760));
    CascadeMux I__4579 (
            .O(N__19774),
            .I(N__19757));
    InMux I__4578 (
            .O(N__19773),
            .I(N__19753));
    InMux I__4577 (
            .O(N__19770),
            .I(N__19750));
    LocalMux I__4576 (
            .O(N__19763),
            .I(N__19747));
    InMux I__4575 (
            .O(N__19760),
            .I(N__19744));
    InMux I__4574 (
            .O(N__19757),
            .I(N__19741));
    InMux I__4573 (
            .O(N__19756),
            .I(N__19736));
    LocalMux I__4572 (
            .O(N__19753),
            .I(N__19733));
    LocalMux I__4571 (
            .O(N__19750),
            .I(N__19726));
    Span4Mux_v I__4570 (
            .O(N__19747),
            .I(N__19726));
    LocalMux I__4569 (
            .O(N__19744),
            .I(N__19726));
    LocalMux I__4568 (
            .O(N__19741),
            .I(N__19723));
    InMux I__4567 (
            .O(N__19740),
            .I(N__19720));
    InMux I__4566 (
            .O(N__19739),
            .I(N__19717));
    LocalMux I__4565 (
            .O(N__19736),
            .I(N__19712));
    Span4Mux_s2_v I__4564 (
            .O(N__19733),
            .I(N__19712));
    Span4Mux_h I__4563 (
            .O(N__19726),
            .I(N__19709));
    Odrv4 I__4562 (
            .O(N__19723),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4561 (
            .O(N__19720),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4560 (
            .O(N__19717),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4559 (
            .O(N__19712),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4558 (
            .O(N__19709),
            .I(bu_rx_data_2_rep1));
    InMux I__4557 (
            .O(N__19698),
            .I(N__19692));
    InMux I__4556 (
            .O(N__19697),
            .I(N__19688));
    InMux I__4555 (
            .O(N__19696),
            .I(N__19684));
    InMux I__4554 (
            .O(N__19695),
            .I(N__19681));
    LocalMux I__4553 (
            .O(N__19692),
            .I(N__19678));
    InMux I__4552 (
            .O(N__19691),
            .I(N__19675));
    LocalMux I__4551 (
            .O(N__19688),
            .I(N__19672));
    InMux I__4550 (
            .O(N__19687),
            .I(N__19669));
    LocalMux I__4549 (
            .O(N__19684),
            .I(N__19663));
    LocalMux I__4548 (
            .O(N__19681),
            .I(N__19663));
    Span4Mux_h I__4547 (
            .O(N__19678),
            .I(N__19660));
    LocalMux I__4546 (
            .O(N__19675),
            .I(N__19653));
    Span4Mux_v I__4545 (
            .O(N__19672),
            .I(N__19653));
    LocalMux I__4544 (
            .O(N__19669),
            .I(N__19653));
    InMux I__4543 (
            .O(N__19668),
            .I(N__19650));
    Odrv4 I__4542 (
            .O(N__19663),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__4541 (
            .O(N__19660),
            .I(bu_rx_data_0_rep1));
    Odrv4 I__4540 (
            .O(N__19653),
            .I(bu_rx_data_0_rep1));
    LocalMux I__4539 (
            .O(N__19650),
            .I(bu_rx_data_0_rep1));
    InMux I__4538 (
            .O(N__19641),
            .I(N__19635));
    InMux I__4537 (
            .O(N__19640),
            .I(N__19635));
    LocalMux I__4536 (
            .O(N__19635),
            .I(N__19632));
    Odrv4 I__4535 (
            .O(N__19632),
            .I(\Lab_UT.dictrl.N_67_mux ));
    CascadeMux I__4534 (
            .O(N__19629),
            .I(N__19623));
    CascadeMux I__4533 (
            .O(N__19628),
            .I(N__19619));
    CascadeMux I__4532 (
            .O(N__19627),
            .I(N__19614));
    InMux I__4531 (
            .O(N__19626),
            .I(N__19611));
    InMux I__4530 (
            .O(N__19623),
            .I(N__19608));
    CascadeMux I__4529 (
            .O(N__19622),
            .I(N__19602));
    InMux I__4528 (
            .O(N__19619),
            .I(N__19597));
    InMux I__4527 (
            .O(N__19618),
            .I(N__19590));
    InMux I__4526 (
            .O(N__19617),
            .I(N__19585));
    InMux I__4525 (
            .O(N__19614),
            .I(N__19585));
    LocalMux I__4524 (
            .O(N__19611),
            .I(N__19582));
    LocalMux I__4523 (
            .O(N__19608),
            .I(N__19578));
    InMux I__4522 (
            .O(N__19607),
            .I(N__19575));
    InMux I__4521 (
            .O(N__19606),
            .I(N__19570));
    InMux I__4520 (
            .O(N__19605),
            .I(N__19570));
    InMux I__4519 (
            .O(N__19602),
            .I(N__19565));
    InMux I__4518 (
            .O(N__19601),
            .I(N__19565));
    InMux I__4517 (
            .O(N__19600),
            .I(N__19562));
    LocalMux I__4516 (
            .O(N__19597),
            .I(N__19559));
    InMux I__4515 (
            .O(N__19596),
            .I(N__19556));
    InMux I__4514 (
            .O(N__19595),
            .I(N__19549));
    InMux I__4513 (
            .O(N__19594),
            .I(N__19549));
    InMux I__4512 (
            .O(N__19593),
            .I(N__19549));
    LocalMux I__4511 (
            .O(N__19590),
            .I(N__19542));
    LocalMux I__4510 (
            .O(N__19585),
            .I(N__19542));
    Span4Mux_v I__4509 (
            .O(N__19582),
            .I(N__19542));
    InMux I__4508 (
            .O(N__19581),
            .I(N__19539));
    Span4Mux_h I__4507 (
            .O(N__19578),
            .I(N__19528));
    LocalMux I__4506 (
            .O(N__19575),
            .I(N__19528));
    LocalMux I__4505 (
            .O(N__19570),
            .I(N__19528));
    LocalMux I__4504 (
            .O(N__19565),
            .I(N__19528));
    LocalMux I__4503 (
            .O(N__19562),
            .I(N__19528));
    Odrv4 I__4502 (
            .O(N__19559),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4501 (
            .O(N__19556),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4500 (
            .O(N__19549),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4499 (
            .O(N__19542),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    LocalMux I__4498 (
            .O(N__19539),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    Odrv4 I__4497 (
            .O(N__19528),
            .I(\Lab_UT.dictrl.stateZ0Z_3 ));
    CascadeMux I__4496 (
            .O(N__19515),
            .I(G_6_0_a6_3_3_cascade_));
    InMux I__4495 (
            .O(N__19512),
            .I(N__19503));
    InMux I__4494 (
            .O(N__19511),
            .I(N__19497));
    InMux I__4493 (
            .O(N__19510),
            .I(N__19491));
    InMux I__4492 (
            .O(N__19509),
            .I(N__19491));
    CascadeMux I__4491 (
            .O(N__19508),
            .I(N__19488));
    InMux I__4490 (
            .O(N__19507),
            .I(N__19485));
    InMux I__4489 (
            .O(N__19506),
            .I(N__19482));
    LocalMux I__4488 (
            .O(N__19503),
            .I(N__19479));
    InMux I__4487 (
            .O(N__19502),
            .I(N__19472));
    InMux I__4486 (
            .O(N__19501),
            .I(N__19472));
    InMux I__4485 (
            .O(N__19500),
            .I(N__19472));
    LocalMux I__4484 (
            .O(N__19497),
            .I(N__19468));
    InMux I__4483 (
            .O(N__19496),
            .I(N__19465));
    LocalMux I__4482 (
            .O(N__19491),
            .I(N__19462));
    InMux I__4481 (
            .O(N__19488),
            .I(N__19455));
    LocalMux I__4480 (
            .O(N__19485),
            .I(N__19452));
    LocalMux I__4479 (
            .O(N__19482),
            .I(N__19445));
    Span4Mux_v I__4478 (
            .O(N__19479),
            .I(N__19445));
    LocalMux I__4477 (
            .O(N__19472),
            .I(N__19445));
    InMux I__4476 (
            .O(N__19471),
            .I(N__19442));
    Span4Mux_h I__4475 (
            .O(N__19468),
            .I(N__19435));
    LocalMux I__4474 (
            .O(N__19465),
            .I(N__19435));
    Span4Mux_h I__4473 (
            .O(N__19462),
            .I(N__19435));
    InMux I__4472 (
            .O(N__19461),
            .I(N__19430));
    InMux I__4471 (
            .O(N__19460),
            .I(N__19430));
    InMux I__4470 (
            .O(N__19459),
            .I(N__19427));
    InMux I__4469 (
            .O(N__19458),
            .I(N__19424));
    LocalMux I__4468 (
            .O(N__19455),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4467 (
            .O(N__19452),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4466 (
            .O(N__19445),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4465 (
            .O(N__19442),
            .I(\Lab_UT.stateZ0Z_0 ));
    Odrv4 I__4464 (
            .O(N__19435),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4463 (
            .O(N__19430),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4462 (
            .O(N__19427),
            .I(\Lab_UT.stateZ0Z_0 ));
    LocalMux I__4461 (
            .O(N__19424),
            .I(\Lab_UT.stateZ0Z_0 ));
    InMux I__4460 (
            .O(N__19407),
            .I(N__19404));
    LocalMux I__4459 (
            .O(N__19404),
            .I(\Lab_UT.dictrl.N_12 ));
    InMux I__4458 (
            .O(N__19401),
            .I(N__19397));
    InMux I__4457 (
            .O(N__19400),
            .I(N__19394));
    LocalMux I__4456 (
            .O(N__19397),
            .I(N__19388));
    LocalMux I__4455 (
            .O(N__19394),
            .I(N__19385));
    InMux I__4454 (
            .O(N__19393),
            .I(N__19382));
    InMux I__4453 (
            .O(N__19392),
            .I(N__19377));
    InMux I__4452 (
            .O(N__19391),
            .I(N__19377));
    Span4Mux_v I__4451 (
            .O(N__19388),
            .I(N__19374));
    Span4Mux_h I__4450 (
            .O(N__19385),
            .I(N__19371));
    LocalMux I__4449 (
            .O(N__19382),
            .I(bu_rx_data_fast_1));
    LocalMux I__4448 (
            .O(N__19377),
            .I(bu_rx_data_fast_1));
    Odrv4 I__4447 (
            .O(N__19374),
            .I(bu_rx_data_fast_1));
    Odrv4 I__4446 (
            .O(N__19371),
            .I(bu_rx_data_fast_1));
    InMux I__4445 (
            .O(N__19362),
            .I(N__19352));
    InMux I__4444 (
            .O(N__19361),
            .I(N__19352));
    InMux I__4443 (
            .O(N__19360),
            .I(N__19352));
    InMux I__4442 (
            .O(N__19359),
            .I(N__19349));
    LocalMux I__4441 (
            .O(N__19352),
            .I(N__19342));
    LocalMux I__4440 (
            .O(N__19349),
            .I(N__19339));
    InMux I__4439 (
            .O(N__19348),
            .I(N__19333));
    InMux I__4438 (
            .O(N__19347),
            .I(N__19333));
    InMux I__4437 (
            .O(N__19346),
            .I(N__19330));
    InMux I__4436 (
            .O(N__19345),
            .I(N__19327));
    Span4Mux_v I__4435 (
            .O(N__19342),
            .I(N__19322));
    Span4Mux_h I__4434 (
            .O(N__19339),
            .I(N__19322));
    InMux I__4433 (
            .O(N__19338),
            .I(N__19319));
    LocalMux I__4432 (
            .O(N__19333),
            .I(N__19316));
    LocalMux I__4431 (
            .O(N__19330),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4430 (
            .O(N__19327),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__4429 (
            .O(N__19322),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4428 (
            .O(N__19319),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__4427 (
            .O(N__19316),
            .I(bu_rx_data_1_rep1));
    InMux I__4426 (
            .O(N__19305),
            .I(N__19301));
    InMux I__4425 (
            .O(N__19304),
            .I(N__19298));
    LocalMux I__4424 (
            .O(N__19301),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    LocalMux I__4423 (
            .O(N__19298),
            .I(\Lab_UT.dictrl.next_state_0_0 ));
    CascadeMux I__4422 (
            .O(N__19293),
            .I(N__19283));
    InMux I__4421 (
            .O(N__19292),
            .I(N__19278));
    InMux I__4420 (
            .O(N__19291),
            .I(N__19275));
    InMux I__4419 (
            .O(N__19290),
            .I(N__19272));
    InMux I__4418 (
            .O(N__19289),
            .I(N__19265));
    InMux I__4417 (
            .O(N__19288),
            .I(N__19265));
    InMux I__4416 (
            .O(N__19287),
            .I(N__19265));
    InMux I__4415 (
            .O(N__19286),
            .I(N__19258));
    InMux I__4414 (
            .O(N__19283),
            .I(N__19258));
    InMux I__4413 (
            .O(N__19282),
            .I(N__19258));
    CascadeMux I__4412 (
            .O(N__19281),
            .I(N__19249));
    LocalMux I__4411 (
            .O(N__19278),
            .I(N__19242));
    LocalMux I__4410 (
            .O(N__19275),
            .I(N__19242));
    LocalMux I__4409 (
            .O(N__19272),
            .I(N__19235));
    LocalMux I__4408 (
            .O(N__19265),
            .I(N__19235));
    LocalMux I__4407 (
            .O(N__19258),
            .I(N__19235));
    InMux I__4406 (
            .O(N__19257),
            .I(N__19232));
    CascadeMux I__4405 (
            .O(N__19256),
            .I(N__19224));
    InMux I__4404 (
            .O(N__19255),
            .I(N__19217));
    InMux I__4403 (
            .O(N__19254),
            .I(N__19217));
    InMux I__4402 (
            .O(N__19253),
            .I(N__19217));
    InMux I__4401 (
            .O(N__19252),
            .I(N__19214));
    InMux I__4400 (
            .O(N__19249),
            .I(N__19211));
    InMux I__4399 (
            .O(N__19248),
            .I(N__19206));
    InMux I__4398 (
            .O(N__19247),
            .I(N__19206));
    Span4Mux_v I__4397 (
            .O(N__19242),
            .I(N__19201));
    Span4Mux_v I__4396 (
            .O(N__19235),
            .I(N__19201));
    LocalMux I__4395 (
            .O(N__19232),
            .I(N__19198));
    InMux I__4394 (
            .O(N__19231),
            .I(N__19191));
    InMux I__4393 (
            .O(N__19230),
            .I(N__19191));
    InMux I__4392 (
            .O(N__19229),
            .I(N__19191));
    InMux I__4391 (
            .O(N__19228),
            .I(N__19184));
    InMux I__4390 (
            .O(N__19227),
            .I(N__19184));
    InMux I__4389 (
            .O(N__19224),
            .I(N__19184));
    LocalMux I__4388 (
            .O(N__19217),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4387 (
            .O(N__19214),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4386 (
            .O(N__19211),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4385 (
            .O(N__19206),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv4 I__4384 (
            .O(N__19201),
            .I(\Lab_UT.un1_next_state66_0 ));
    Odrv4 I__4383 (
            .O(N__19198),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4382 (
            .O(N__19191),
            .I(\Lab_UT.un1_next_state66_0 ));
    LocalMux I__4381 (
            .O(N__19184),
            .I(\Lab_UT.un1_next_state66_0 ));
    CascadeMux I__4380 (
            .O(N__19167),
            .I(\Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ));
    CascadeMux I__4379 (
            .O(N__19164),
            .I(N__19160));
    InMux I__4378 (
            .O(N__19163),
            .I(N__19155));
    InMux I__4377 (
            .O(N__19160),
            .I(N__19155));
    LocalMux I__4376 (
            .O(N__19155),
            .I(\Lab_UT.dictrl.N_60 ));
    CascadeMux I__4375 (
            .O(N__19152),
            .I(N__19149));
    InMux I__4374 (
            .O(N__19149),
            .I(N__19143));
    InMux I__4373 (
            .O(N__19148),
            .I(N__19143));
    LocalMux I__4372 (
            .O(N__19143),
            .I(N__19140));
    Odrv12 I__4371 (
            .O(N__19140),
            .I(\Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ));
    InMux I__4370 (
            .O(N__19137),
            .I(N__19130));
    InMux I__4369 (
            .O(N__19136),
            .I(N__19127));
    InMux I__4368 (
            .O(N__19135),
            .I(N__19124));
    InMux I__4367 (
            .O(N__19134),
            .I(N__19121));
    CascadeMux I__4366 (
            .O(N__19133),
            .I(N__19117));
    LocalMux I__4365 (
            .O(N__19130),
            .I(N__19114));
    LocalMux I__4364 (
            .O(N__19127),
            .I(N__19107));
    LocalMux I__4363 (
            .O(N__19124),
            .I(N__19107));
    LocalMux I__4362 (
            .O(N__19121),
            .I(N__19107));
    InMux I__4361 (
            .O(N__19120),
            .I(N__19104));
    InMux I__4360 (
            .O(N__19117),
            .I(N__19100));
    Span4Mux_v I__4359 (
            .O(N__19114),
            .I(N__19097));
    Span4Mux_v I__4358 (
            .O(N__19107),
            .I(N__19094));
    LocalMux I__4357 (
            .O(N__19104),
            .I(N__19091));
    InMux I__4356 (
            .O(N__19103),
            .I(N__19088));
    LocalMux I__4355 (
            .O(N__19100),
            .I(\Lab_UT.dicLdSones_1 ));
    Odrv4 I__4354 (
            .O(N__19097),
            .I(\Lab_UT.dicLdSones_1 ));
    Odrv4 I__4353 (
            .O(N__19094),
            .I(\Lab_UT.dicLdSones_1 ));
    Odrv4 I__4352 (
            .O(N__19091),
            .I(\Lab_UT.dicLdSones_1 ));
    LocalMux I__4351 (
            .O(N__19088),
            .I(\Lab_UT.dicLdSones_1 ));
    CascadeMux I__4350 (
            .O(N__19077),
            .I(G_6_0_a6_2_cascade_));
    InMux I__4349 (
            .O(N__19074),
            .I(N__19071));
    LocalMux I__4348 (
            .O(N__19071),
            .I(\Lab_UT.dictrl.G_6_0_0_1 ));
    CascadeMux I__4347 (
            .O(N__19068),
            .I(\Lab_UT.dictrl.G_6_0_0_cascade_ ));
    InMux I__4346 (
            .O(N__19065),
            .I(N__19062));
    LocalMux I__4345 (
            .O(N__19062),
            .I(N__19059));
    Odrv4 I__4344 (
            .O(N__19059),
            .I(\Lab_UT.dictrl.G_6_0_1_0 ));
    InMux I__4343 (
            .O(N__19056),
            .I(N__19050));
    InMux I__4342 (
            .O(N__19055),
            .I(N__19050));
    LocalMux I__4341 (
            .O(N__19050),
            .I(N__19047));
    Span4Mux_h I__4340 (
            .O(N__19047),
            .I(N__19044));
    Odrv4 I__4339 (
            .O(N__19044),
            .I(\Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ));
    InMux I__4338 (
            .O(N__19041),
            .I(N__19037));
    InMux I__4337 (
            .O(N__19040),
            .I(N__19033));
    LocalMux I__4336 (
            .O(N__19037),
            .I(N__19030));
    CascadeMux I__4335 (
            .O(N__19036),
            .I(N__19024));
    LocalMux I__4334 (
            .O(N__19033),
            .I(N__19019));
    Span4Mux_v I__4333 (
            .O(N__19030),
            .I(N__19019));
    InMux I__4332 (
            .O(N__19029),
            .I(N__19016));
    InMux I__4331 (
            .O(N__19028),
            .I(N__19011));
    InMux I__4330 (
            .O(N__19027),
            .I(N__19011));
    InMux I__4329 (
            .O(N__19024),
            .I(N__19008));
    Odrv4 I__4328 (
            .O(N__19019),
            .I(\Lab_UT.dictrl.m13_out ));
    LocalMux I__4327 (
            .O(N__19016),
            .I(\Lab_UT.dictrl.m13_out ));
    LocalMux I__4326 (
            .O(N__19011),
            .I(\Lab_UT.dictrl.m13_out ));
    LocalMux I__4325 (
            .O(N__19008),
            .I(\Lab_UT.dictrl.m13_out ));
    InMux I__4324 (
            .O(N__18999),
            .I(N__18993));
    InMux I__4323 (
            .O(N__18998),
            .I(N__18993));
    LocalMux I__4322 (
            .O(N__18993),
            .I(N__18990));
    Odrv4 I__4321 (
            .O(N__18990),
            .I(\Lab_UT.dictrl.N_15_0 ));
    InMux I__4320 (
            .O(N__18987),
            .I(N__18983));
    InMux I__4319 (
            .O(N__18986),
            .I(N__18978));
    LocalMux I__4318 (
            .O(N__18983),
            .I(N__18975));
    InMux I__4317 (
            .O(N__18982),
            .I(N__18970));
    InMux I__4316 (
            .O(N__18981),
            .I(N__18970));
    LocalMux I__4315 (
            .O(N__18978),
            .I(\Lab_UT.dictrl.N_72_mux ));
    Odrv4 I__4314 (
            .O(N__18975),
            .I(\Lab_UT.dictrl.N_72_mux ));
    LocalMux I__4313 (
            .O(N__18970),
            .I(\Lab_UT.dictrl.N_72_mux ));
    InMux I__4312 (
            .O(N__18963),
            .I(N__18957));
    InMux I__4311 (
            .O(N__18962),
            .I(N__18957));
    LocalMux I__4310 (
            .O(N__18957),
            .I(\Lab_UT.dictrl.N_59 ));
    CascadeMux I__4309 (
            .O(N__18954),
            .I(shifter_1_rep1_RNI0FPF_cascade_));
    InMux I__4308 (
            .O(N__18951),
            .I(N__18945));
    InMux I__4307 (
            .O(N__18950),
            .I(N__18945));
    LocalMux I__4306 (
            .O(N__18945),
            .I(\Lab_UT.dictrl.N_33_0 ));
    CascadeMux I__4305 (
            .O(N__18942),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ));
    CascadeMux I__4304 (
            .O(N__18939),
            .I(N__18935));
    CascadeMux I__4303 (
            .O(N__18938),
            .I(N__18932));
    InMux I__4302 (
            .O(N__18935),
            .I(N__18925));
    InMux I__4301 (
            .O(N__18932),
            .I(N__18925));
    InMux I__4300 (
            .O(N__18931),
            .I(N__18920));
    InMux I__4299 (
            .O(N__18930),
            .I(N__18920));
    LocalMux I__4298 (
            .O(N__18925),
            .I(\Lab_UT.dictrl.G_14_0_1 ));
    LocalMux I__4297 (
            .O(N__18920),
            .I(\Lab_UT.dictrl.G_14_0_1 ));
    CascadeMux I__4296 (
            .O(N__18915),
            .I(N__18910));
    CascadeMux I__4295 (
            .O(N__18914),
            .I(N__18907));
    CascadeMux I__4294 (
            .O(N__18913),
            .I(N__18898));
    InMux I__4293 (
            .O(N__18910),
            .I(N__18891));
    InMux I__4292 (
            .O(N__18907),
            .I(N__18891));
    InMux I__4291 (
            .O(N__18906),
            .I(N__18891));
    CascadeMux I__4290 (
            .O(N__18905),
            .I(N__18888));
    CascadeMux I__4289 (
            .O(N__18904),
            .I(N__18883));
    CascadeMux I__4288 (
            .O(N__18903),
            .I(N__18880));
    InMux I__4287 (
            .O(N__18902),
            .I(N__18877));
    InMux I__4286 (
            .O(N__18901),
            .I(N__18872));
    InMux I__4285 (
            .O(N__18898),
            .I(N__18872));
    LocalMux I__4284 (
            .O(N__18891),
            .I(N__18869));
    InMux I__4283 (
            .O(N__18888),
            .I(N__18864));
    InMux I__4282 (
            .O(N__18887),
            .I(N__18864));
    InMux I__4281 (
            .O(N__18886),
            .I(N__18861));
    InMux I__4280 (
            .O(N__18883),
            .I(N__18858));
    InMux I__4279 (
            .O(N__18880),
            .I(N__18855));
    LocalMux I__4278 (
            .O(N__18877),
            .I(N__18846));
    LocalMux I__4277 (
            .O(N__18872),
            .I(N__18846));
    Span12Mux_s4_h I__4276 (
            .O(N__18869),
            .I(N__18846));
    LocalMux I__4275 (
            .O(N__18864),
            .I(N__18846));
    LocalMux I__4274 (
            .O(N__18861),
            .I(bu_rx_data_3_rep1));
    LocalMux I__4273 (
            .O(N__18858),
            .I(bu_rx_data_3_rep1));
    LocalMux I__4272 (
            .O(N__18855),
            .I(bu_rx_data_3_rep1));
    Odrv12 I__4271 (
            .O(N__18846),
            .I(bu_rx_data_3_rep1));
    InMux I__4270 (
            .O(N__18837),
            .I(N__18834));
    LocalMux I__4269 (
            .O(N__18834),
            .I(N__18831));
    Odrv12 I__4268 (
            .O(N__18831),
            .I(\Lab_UT.dictrl.G_14_0_a2_1 ));
    CascadeMux I__4267 (
            .O(N__18828),
            .I(N_15_cascade_));
    CascadeMux I__4266 (
            .O(N__18825),
            .I(N__18819));
    CascadeMux I__4265 (
            .O(N__18824),
            .I(N__18816));
    InMux I__4264 (
            .O(N__18823),
            .I(N__18807));
    InMux I__4263 (
            .O(N__18822),
            .I(N__18807));
    InMux I__4262 (
            .O(N__18819),
            .I(N__18807));
    InMux I__4261 (
            .O(N__18816),
            .I(N__18807));
    LocalMux I__4260 (
            .O(N__18807),
            .I(\Lab_UT.dictrl.N_20_0 ));
    CascadeMux I__4259 (
            .O(N__18804),
            .I(N__18800));
    InMux I__4258 (
            .O(N__18803),
            .I(N__18794));
    InMux I__4257 (
            .O(N__18800),
            .I(N__18794));
    InMux I__4256 (
            .O(N__18799),
            .I(N__18791));
    LocalMux I__4255 (
            .O(N__18794),
            .I(N__18788));
    LocalMux I__4254 (
            .O(N__18791),
            .I(N__18785));
    Span4Mux_h I__4253 (
            .O(N__18788),
            .I(N__18782));
    Span4Mux_h I__4252 (
            .O(N__18785),
            .I(N__18779));
    Odrv4 I__4251 (
            .O(N__18782),
            .I(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ));
    Odrv4 I__4250 (
            .O(N__18779),
            .I(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ));
    CascadeMux I__4249 (
            .O(N__18774),
            .I(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ));
    CEMux I__4248 (
            .O(N__18771),
            .I(N__18768));
    LocalMux I__4247 (
            .O(N__18768),
            .I(N__18765));
    Span4Mux_v I__4246 (
            .O(N__18765),
            .I(N__18760));
    CEMux I__4245 (
            .O(N__18764),
            .I(N__18757));
    CEMux I__4244 (
            .O(N__18763),
            .I(N__18754));
    Span4Mux_v I__4243 (
            .O(N__18760),
            .I(N__18749));
    LocalMux I__4242 (
            .O(N__18757),
            .I(N__18749));
    LocalMux I__4241 (
            .O(N__18754),
            .I(N__18745));
    Span4Mux_v I__4240 (
            .O(N__18749),
            .I(N__18742));
    CEMux I__4239 (
            .O(N__18748),
            .I(N__18739));
    Span4Mux_v I__4238 (
            .O(N__18745),
            .I(N__18736));
    Span4Mux_h I__4237 (
            .O(N__18742),
            .I(N__18731));
    LocalMux I__4236 (
            .O(N__18739),
            .I(N__18731));
    Span4Mux_s2_h I__4235 (
            .O(N__18736),
            .I(N__18728));
    Span4Mux_h I__4234 (
            .O(N__18731),
            .I(N__18725));
    Odrv4 I__4233 (
            .O(N__18728),
            .I(\Lab_UT.g0_0 ));
    Odrv4 I__4232 (
            .O(N__18725),
            .I(\Lab_UT.g0_0 ));
    CascadeMux I__4231 (
            .O(N__18720),
            .I(\Lab_UT.dictrl.N_15_0_cascade_ ));
    CascadeMux I__4230 (
            .O(N__18717),
            .I(\Lab_UT.dictrl.N_60_cascade_ ));
    InMux I__4229 (
            .O(N__18714),
            .I(N__18711));
    LocalMux I__4228 (
            .O(N__18711),
            .I(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ));
    InMux I__4227 (
            .O(N__18708),
            .I(N__18705));
    LocalMux I__4226 (
            .O(N__18705),
            .I(N__18701));
    InMux I__4225 (
            .O(N__18704),
            .I(N__18697));
    Span4Mux_v I__4224 (
            .O(N__18701),
            .I(N__18694));
    InMux I__4223 (
            .O(N__18700),
            .I(N__18691));
    LocalMux I__4222 (
            .O(N__18697),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    Odrv4 I__4221 (
            .O(N__18694),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    LocalMux I__4220 (
            .O(N__18691),
            .I(\Lab_UT.dictrl.state_i_4_1 ));
    InMux I__4219 (
            .O(N__18684),
            .I(N__18681));
    LocalMux I__4218 (
            .O(N__18681),
            .I(N__18678));
    Span4Mux_h I__4217 (
            .O(N__18678),
            .I(N__18675));
    Odrv4 I__4216 (
            .O(N__18675),
            .I(\Lab_UT.dictrl.m19_1_0 ));
    InMux I__4215 (
            .O(N__18672),
            .I(N__18667));
    InMux I__4214 (
            .O(N__18671),
            .I(N__18662));
    InMux I__4213 (
            .O(N__18670),
            .I(N__18662));
    LocalMux I__4212 (
            .O(N__18667),
            .I(N__18657));
    LocalMux I__4211 (
            .O(N__18662),
            .I(N__18657));
    Odrv4 I__4210 (
            .O(N__18657),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    CascadeMux I__4209 (
            .O(N__18654),
            .I(N__18651));
    InMux I__4208 (
            .O(N__18651),
            .I(N__18644));
    InMux I__4207 (
            .O(N__18650),
            .I(N__18644));
    CascadeMux I__4206 (
            .O(N__18649),
            .I(N__18641));
    LocalMux I__4205 (
            .O(N__18644),
            .I(N__18638));
    InMux I__4204 (
            .O(N__18641),
            .I(N__18635));
    Span4Mux_h I__4203 (
            .O(N__18638),
            .I(N__18630));
    LocalMux I__4202 (
            .O(N__18635),
            .I(N__18630));
    Span4Mux_v I__4201 (
            .O(N__18630),
            .I(N__18625));
    InMux I__4200 (
            .O(N__18629),
            .I(N__18622));
    InMux I__4199 (
            .O(N__18628),
            .I(N__18619));
    Odrv4 I__4198 (
            .O(N__18625),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    LocalMux I__4197 (
            .O(N__18622),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    LocalMux I__4196 (
            .O(N__18619),
            .I(\Lab_UT.dictrl.next_state_0_3 ));
    CascadeMux I__4195 (
            .O(N__18612),
            .I(N__18608));
    CascadeMux I__4194 (
            .O(N__18611),
            .I(N__18604));
    InMux I__4193 (
            .O(N__18608),
            .I(N__18593));
    InMux I__4192 (
            .O(N__18607),
            .I(N__18593));
    InMux I__4191 (
            .O(N__18604),
            .I(N__18593));
    InMux I__4190 (
            .O(N__18603),
            .I(N__18593));
    InMux I__4189 (
            .O(N__18602),
            .I(N__18587));
    LocalMux I__4188 (
            .O(N__18593),
            .I(N__18584));
    InMux I__4187 (
            .O(N__18592),
            .I(N__18579));
    InMux I__4186 (
            .O(N__18591),
            .I(N__18579));
    InMux I__4185 (
            .O(N__18590),
            .I(N__18576));
    LocalMux I__4184 (
            .O(N__18587),
            .I(N__18573));
    Sp12to4 I__4183 (
            .O(N__18584),
            .I(N__18568));
    LocalMux I__4182 (
            .O(N__18579),
            .I(N__18568));
    LocalMux I__4181 (
            .O(N__18576),
            .I(\Lab_UT.next_state_1 ));
    Odrv4 I__4180 (
            .O(N__18573),
            .I(\Lab_UT.next_state_1 ));
    Odrv12 I__4179 (
            .O(N__18568),
            .I(\Lab_UT.next_state_1 ));
    CascadeMux I__4178 (
            .O(N__18561),
            .I(N__18558));
    InMux I__4177 (
            .O(N__18558),
            .I(N__18554));
    InMux I__4176 (
            .O(N__18557),
            .I(N__18551));
    LocalMux I__4175 (
            .O(N__18554),
            .I(N__18546));
    LocalMux I__4174 (
            .O(N__18551),
            .I(N__18543));
    InMux I__4173 (
            .O(N__18550),
            .I(N__18538));
    InMux I__4172 (
            .O(N__18549),
            .I(N__18538));
    Span4Mux_h I__4171 (
            .O(N__18546),
            .I(N__18535));
    Span4Mux_v I__4170 (
            .O(N__18543),
            .I(N__18530));
    LocalMux I__4169 (
            .O(N__18538),
            .I(N__18530));
    Span4Mux_v I__4168 (
            .O(N__18535),
            .I(N__18527));
    Span4Mux_h I__4167 (
            .O(N__18530),
            .I(N__18524));
    Odrv4 I__4166 (
            .O(N__18527),
            .I(\Lab_UT.dictrl.next_state66_2 ));
    Odrv4 I__4165 (
            .O(N__18524),
            .I(\Lab_UT.dictrl.next_state66_2 ));
    CEMux I__4164 (
            .O(N__18519),
            .I(N__18516));
    LocalMux I__4163 (
            .O(N__18516),
            .I(N__18511));
    CEMux I__4162 (
            .O(N__18515),
            .I(N__18508));
    CEMux I__4161 (
            .O(N__18514),
            .I(N__18504));
    Span4Mux_s3_h I__4160 (
            .O(N__18511),
            .I(N__18499));
    LocalMux I__4159 (
            .O(N__18508),
            .I(N__18499));
    CEMux I__4158 (
            .O(N__18507),
            .I(N__18496));
    LocalMux I__4157 (
            .O(N__18504),
            .I(N__18493));
    Span4Mux_v I__4156 (
            .O(N__18499),
            .I(N__18488));
    LocalMux I__4155 (
            .O(N__18496),
            .I(N__18488));
    Span4Mux_h I__4154 (
            .O(N__18493),
            .I(N__18483));
    Span4Mux_h I__4153 (
            .O(N__18488),
            .I(N__18483));
    Odrv4 I__4152 (
            .O(N__18483),
            .I(\Lab_UT.bu_rx_data_rdy_0 ));
    InMux I__4151 (
            .O(N__18480),
            .I(N__18474));
    CascadeMux I__4150 (
            .O(N__18479),
            .I(N__18470));
    InMux I__4149 (
            .O(N__18478),
            .I(N__18465));
    InMux I__4148 (
            .O(N__18477),
            .I(N__18462));
    LocalMux I__4147 (
            .O(N__18474),
            .I(N__18459));
    InMux I__4146 (
            .O(N__18473),
            .I(N__18456));
    InMux I__4145 (
            .O(N__18470),
            .I(N__18452));
    CascadeMux I__4144 (
            .O(N__18469),
            .I(N__18449));
    CascadeMux I__4143 (
            .O(N__18468),
            .I(N__18446));
    LocalMux I__4142 (
            .O(N__18465),
            .I(N__18442));
    LocalMux I__4141 (
            .O(N__18462),
            .I(N__18438));
    Span4Mux_s3_v I__4140 (
            .O(N__18459),
            .I(N__18433));
    LocalMux I__4139 (
            .O(N__18456),
            .I(N__18433));
    InMux I__4138 (
            .O(N__18455),
            .I(N__18430));
    LocalMux I__4137 (
            .O(N__18452),
            .I(N__18427));
    InMux I__4136 (
            .O(N__18449),
            .I(N__18424));
    InMux I__4135 (
            .O(N__18446),
            .I(N__18413));
    InMux I__4134 (
            .O(N__18445),
            .I(N__18413));
    Span4Mux_v I__4133 (
            .O(N__18442),
            .I(N__18410));
    InMux I__4132 (
            .O(N__18441),
            .I(N__18407));
    Span4Mux_h I__4131 (
            .O(N__18438),
            .I(N__18396));
    Span4Mux_v I__4130 (
            .O(N__18433),
            .I(N__18396));
    LocalMux I__4129 (
            .O(N__18430),
            .I(N__18396));
    Span4Mux_h I__4128 (
            .O(N__18427),
            .I(N__18396));
    LocalMux I__4127 (
            .O(N__18424),
            .I(N__18396));
    InMux I__4126 (
            .O(N__18423),
            .I(N__18387));
    InMux I__4125 (
            .O(N__18422),
            .I(N__18387));
    InMux I__4124 (
            .O(N__18421),
            .I(N__18387));
    InMux I__4123 (
            .O(N__18420),
            .I(N__18387));
    InMux I__4122 (
            .O(N__18419),
            .I(N__18384));
    InMux I__4121 (
            .O(N__18418),
            .I(N__18381));
    LocalMux I__4120 (
            .O(N__18413),
            .I(N__18378));
    Odrv4 I__4119 (
            .O(N__18410),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__4118 (
            .O(N__18407),
            .I(\Lab_UT.state_i_4_3 ));
    Odrv4 I__4117 (
            .O(N__18396),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__4116 (
            .O(N__18387),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__4115 (
            .O(N__18384),
            .I(\Lab_UT.state_i_4_3 ));
    LocalMux I__4114 (
            .O(N__18381),
            .I(\Lab_UT.state_i_4_3 ));
    Odrv4 I__4113 (
            .O(N__18378),
            .I(\Lab_UT.state_i_4_3 ));
    CascadeMux I__4112 (
            .O(N__18363),
            .I(N__18360));
    InMux I__4111 (
            .O(N__18360),
            .I(N__18356));
    InMux I__4110 (
            .O(N__18359),
            .I(N__18353));
    LocalMux I__4109 (
            .O(N__18356),
            .I(\Lab_UT.dictrl.dicRun_1 ));
    LocalMux I__4108 (
            .O(N__18353),
            .I(\Lab_UT.dictrl.dicRun_1 ));
    InMux I__4107 (
            .O(N__18348),
            .I(N__18342));
    InMux I__4106 (
            .O(N__18347),
            .I(N__18331));
    InMux I__4105 (
            .O(N__18346),
            .I(N__18327));
    InMux I__4104 (
            .O(N__18345),
            .I(N__18324));
    LocalMux I__4103 (
            .O(N__18342),
            .I(N__18321));
    InMux I__4102 (
            .O(N__18341),
            .I(N__18318));
    InMux I__4101 (
            .O(N__18340),
            .I(N__18311));
    InMux I__4100 (
            .O(N__18339),
            .I(N__18311));
    InMux I__4099 (
            .O(N__18338),
            .I(N__18311));
    InMux I__4098 (
            .O(N__18337),
            .I(N__18302));
    InMux I__4097 (
            .O(N__18336),
            .I(N__18302));
    InMux I__4096 (
            .O(N__18335),
            .I(N__18302));
    InMux I__4095 (
            .O(N__18334),
            .I(N__18302));
    LocalMux I__4094 (
            .O(N__18331),
            .I(N__18294));
    InMux I__4093 (
            .O(N__18330),
            .I(N__18291));
    LocalMux I__4092 (
            .O(N__18327),
            .I(N__18288));
    LocalMux I__4091 (
            .O(N__18324),
            .I(N__18285));
    Span4Mux_v I__4090 (
            .O(N__18321),
            .I(N__18278));
    LocalMux I__4089 (
            .O(N__18318),
            .I(N__18278));
    LocalMux I__4088 (
            .O(N__18311),
            .I(N__18278));
    LocalMux I__4087 (
            .O(N__18302),
            .I(N__18275));
    InMux I__4086 (
            .O(N__18301),
            .I(N__18270));
    InMux I__4085 (
            .O(N__18300),
            .I(N__18270));
    InMux I__4084 (
            .O(N__18299),
            .I(N__18263));
    InMux I__4083 (
            .O(N__18298),
            .I(N__18263));
    InMux I__4082 (
            .O(N__18297),
            .I(N__18263));
    Odrv12 I__4081 (
            .O(N__18294),
            .I(\Lab_UT.state_2 ));
    LocalMux I__4080 (
            .O(N__18291),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4079 (
            .O(N__18288),
            .I(\Lab_UT.state_2 ));
    Odrv12 I__4078 (
            .O(N__18285),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4077 (
            .O(N__18278),
            .I(\Lab_UT.state_2 ));
    Odrv4 I__4076 (
            .O(N__18275),
            .I(\Lab_UT.state_2 ));
    LocalMux I__4075 (
            .O(N__18270),
            .I(\Lab_UT.state_2 ));
    LocalMux I__4074 (
            .O(N__18263),
            .I(\Lab_UT.state_2 ));
    InMux I__4073 (
            .O(N__18246),
            .I(N__18243));
    LocalMux I__4072 (
            .O(N__18243),
            .I(N__18240));
    Span4Mux_h I__4071 (
            .O(N__18240),
            .I(N__18236));
    InMux I__4070 (
            .O(N__18239),
            .I(N__18233));
    Odrv4 I__4069 (
            .O(N__18236),
            .I(\Lab_UT.LdASones ));
    LocalMux I__4068 (
            .O(N__18233),
            .I(\Lab_UT.LdASones ));
    InMux I__4067 (
            .O(N__18228),
            .I(N__18223));
    InMux I__4066 (
            .O(N__18227),
            .I(N__18217));
    InMux I__4065 (
            .O(N__18226),
            .I(N__18214));
    LocalMux I__4064 (
            .O(N__18223),
            .I(N__18211));
    InMux I__4063 (
            .O(N__18222),
            .I(N__18208));
    InMux I__4062 (
            .O(N__18221),
            .I(N__18203));
    CascadeMux I__4061 (
            .O(N__18220),
            .I(N__18198));
    LocalMux I__4060 (
            .O(N__18217),
            .I(N__18189));
    LocalMux I__4059 (
            .O(N__18214),
            .I(N__18189));
    Span4Mux_v I__4058 (
            .O(N__18211),
            .I(N__18184));
    LocalMux I__4057 (
            .O(N__18208),
            .I(N__18184));
    InMux I__4056 (
            .O(N__18207),
            .I(N__18181));
    InMux I__4055 (
            .O(N__18206),
            .I(N__18178));
    LocalMux I__4054 (
            .O(N__18203),
            .I(N__18175));
    InMux I__4053 (
            .O(N__18202),
            .I(N__18172));
    InMux I__4052 (
            .O(N__18201),
            .I(N__18167));
    InMux I__4051 (
            .O(N__18198),
            .I(N__18167));
    InMux I__4050 (
            .O(N__18197),
            .I(N__18162));
    InMux I__4049 (
            .O(N__18196),
            .I(N__18162));
    InMux I__4048 (
            .O(N__18195),
            .I(N__18159));
    InMux I__4047 (
            .O(N__18194),
            .I(N__18156));
    Span4Mux_v I__4046 (
            .O(N__18189),
            .I(N__18153));
    Span4Mux_h I__4045 (
            .O(N__18184),
            .I(N__18150));
    LocalMux I__4044 (
            .O(N__18181),
            .I(N__18145));
    LocalMux I__4043 (
            .O(N__18178),
            .I(N__18145));
    Span4Mux_v I__4042 (
            .O(N__18175),
            .I(N__18140));
    LocalMux I__4041 (
            .O(N__18172),
            .I(N__18140));
    LocalMux I__4040 (
            .O(N__18167),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4039 (
            .O(N__18162),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4038 (
            .O(N__18159),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__4037 (
            .O(N__18156),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__4036 (
            .O(N__18153),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__4035 (
            .O(N__18150),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv12 I__4034 (
            .O(N__18145),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__4033 (
            .O(N__18140),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    InMux I__4032 (
            .O(N__18123),
            .I(N__18107));
    InMux I__4031 (
            .O(N__18122),
            .I(N__18107));
    InMux I__4030 (
            .O(N__18121),
            .I(N__18100));
    InMux I__4029 (
            .O(N__18120),
            .I(N__18100));
    InMux I__4028 (
            .O(N__18119),
            .I(N__18100));
    InMux I__4027 (
            .O(N__18118),
            .I(N__18097));
    InMux I__4026 (
            .O(N__18117),
            .I(N__18094));
    InMux I__4025 (
            .O(N__18116),
            .I(N__18087));
    InMux I__4024 (
            .O(N__18115),
            .I(N__18087));
    InMux I__4023 (
            .O(N__18114),
            .I(N__18082));
    InMux I__4022 (
            .O(N__18113),
            .I(N__18082));
    InMux I__4021 (
            .O(N__18112),
            .I(N__18074));
    LocalMux I__4020 (
            .O(N__18107),
            .I(N__18069));
    LocalMux I__4019 (
            .O(N__18100),
            .I(N__18069));
    LocalMux I__4018 (
            .O(N__18097),
            .I(N__18064));
    LocalMux I__4017 (
            .O(N__18094),
            .I(N__18064));
    InMux I__4016 (
            .O(N__18093),
            .I(N__18061));
    InMux I__4015 (
            .O(N__18092),
            .I(N__18058));
    LocalMux I__4014 (
            .O(N__18087),
            .I(N__18053));
    LocalMux I__4013 (
            .O(N__18082),
            .I(N__18053));
    InMux I__4012 (
            .O(N__18081),
            .I(N__18048));
    InMux I__4011 (
            .O(N__18080),
            .I(N__18048));
    InMux I__4010 (
            .O(N__18079),
            .I(N__18043));
    InMux I__4009 (
            .O(N__18078),
            .I(N__18043));
    InMux I__4008 (
            .O(N__18077),
            .I(N__18040));
    LocalMux I__4007 (
            .O(N__18074),
            .I(N__18037));
    Span4Mux_v I__4006 (
            .O(N__18069),
            .I(N__18028));
    Span4Mux_v I__4005 (
            .O(N__18064),
            .I(N__18028));
    LocalMux I__4004 (
            .O(N__18061),
            .I(N__18028));
    LocalMux I__4003 (
            .O(N__18058),
            .I(N__18028));
    Span4Mux_v I__4002 (
            .O(N__18053),
            .I(N__18025));
    LocalMux I__4001 (
            .O(N__18048),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__4000 (
            .O(N__18043),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__3999 (
            .O(N__18040),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv12 I__3998 (
            .O(N__18037),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__3997 (
            .O(N__18028),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__3996 (
            .O(N__18025),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    InMux I__3995 (
            .O(N__18012),
            .I(N__18009));
    LocalMux I__3994 (
            .O(N__18009),
            .I(N__18004));
    CascadeMux I__3993 (
            .O(N__18008),
            .I(N__17999));
    InMux I__3992 (
            .O(N__18007),
            .I(N__17994));
    Span4Mux_v I__3991 (
            .O(N__18004),
            .I(N__17991));
    InMux I__3990 (
            .O(N__18003),
            .I(N__17986));
    InMux I__3989 (
            .O(N__18002),
            .I(N__17986));
    InMux I__3988 (
            .O(N__17999),
            .I(N__17983));
    CascadeMux I__3987 (
            .O(N__17998),
            .I(N__17977));
    InMux I__3986 (
            .O(N__17997),
            .I(N__17972));
    LocalMux I__3985 (
            .O(N__17994),
            .I(N__17963));
    Span4Mux_h I__3984 (
            .O(N__17991),
            .I(N__17963));
    LocalMux I__3983 (
            .O(N__17986),
            .I(N__17963));
    LocalMux I__3982 (
            .O(N__17983),
            .I(N__17963));
    InMux I__3981 (
            .O(N__17982),
            .I(N__17958));
    InMux I__3980 (
            .O(N__17981),
            .I(N__17958));
    InMux I__3979 (
            .O(N__17980),
            .I(N__17955));
    InMux I__3978 (
            .O(N__17977),
            .I(N__17950));
    InMux I__3977 (
            .O(N__17976),
            .I(N__17950));
    InMux I__3976 (
            .O(N__17975),
            .I(N__17947));
    LocalMux I__3975 (
            .O(N__17972),
            .I(N__17940));
    Span4Mux_v I__3974 (
            .O(N__17963),
            .I(N__17940));
    LocalMux I__3973 (
            .O(N__17958),
            .I(N__17940));
    LocalMux I__3972 (
            .O(N__17955),
            .I(N__17935));
    LocalMux I__3971 (
            .O(N__17950),
            .I(N__17935));
    LocalMux I__3970 (
            .O(N__17947),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__3969 (
            .O(N__17940),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__3968 (
            .O(N__17935),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    InMux I__3967 (
            .O(N__17928),
            .I(N__17925));
    LocalMux I__3966 (
            .O(N__17925),
            .I(N__17922));
    Span4Mux_h I__3965 (
            .O(N__17922),
            .I(N__17919));
    Odrv4 I__3964 (
            .O(N__17919),
            .I(\Lab_UT.dictrl.g1_4_0 ));
    CascadeMux I__3963 (
            .O(N__17916),
            .I(\Lab_UT.dictrl.g1_5_0_cascade_ ));
    CascadeMux I__3962 (
            .O(N__17913),
            .I(\Lab_UT.dictrl.G_14_0_a2_4_2_cascade_ ));
    InMux I__3961 (
            .O(N__17910),
            .I(N__17902));
    InMux I__3960 (
            .O(N__17909),
            .I(N__17902));
    InMux I__3959 (
            .O(N__17908),
            .I(N__17897));
    InMux I__3958 (
            .O(N__17907),
            .I(N__17897));
    LocalMux I__3957 (
            .O(N__17902),
            .I(\Lab_UT.dictrl.G_14_0_0 ));
    LocalMux I__3956 (
            .O(N__17897),
            .I(\Lab_UT.dictrl.G_14_0_0 ));
    InMux I__3955 (
            .O(N__17892),
            .I(N__17888));
    CascadeMux I__3954 (
            .O(N__17891),
            .I(N__17885));
    LocalMux I__3953 (
            .O(N__17888),
            .I(N__17878));
    InMux I__3952 (
            .O(N__17885),
            .I(N__17870));
    InMux I__3951 (
            .O(N__17884),
            .I(N__17870));
    InMux I__3950 (
            .O(N__17883),
            .I(N__17870));
    InMux I__3949 (
            .O(N__17882),
            .I(N__17867));
    InMux I__3948 (
            .O(N__17881),
            .I(N__17862));
    Span4Mux_h I__3947 (
            .O(N__17878),
            .I(N__17859));
    InMux I__3946 (
            .O(N__17877),
            .I(N__17856));
    LocalMux I__3945 (
            .O(N__17870),
            .I(N__17853));
    LocalMux I__3944 (
            .O(N__17867),
            .I(N__17850));
    InMux I__3943 (
            .O(N__17866),
            .I(N__17845));
    InMux I__3942 (
            .O(N__17865),
            .I(N__17845));
    LocalMux I__3941 (
            .O(N__17862),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3940 (
            .O(N__17859),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3939 (
            .O(N__17856),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3938 (
            .O(N__17853),
            .I(\Lab_UT.di_Sones_1 ));
    Odrv4 I__3937 (
            .O(N__17850),
            .I(\Lab_UT.di_Sones_1 ));
    LocalMux I__3936 (
            .O(N__17845),
            .I(\Lab_UT.di_Sones_1 ));
    InMux I__3935 (
            .O(N__17832),
            .I(N__17828));
    InMux I__3934 (
            .O(N__17831),
            .I(N__17824));
    LocalMux I__3933 (
            .O(N__17828),
            .I(N__17821));
    InMux I__3932 (
            .O(N__17827),
            .I(N__17818));
    LocalMux I__3931 (
            .O(N__17824),
            .I(N__17815));
    Span4Mux_h I__3930 (
            .O(N__17821),
            .I(N__17812));
    LocalMux I__3929 (
            .O(N__17818),
            .I(N__17809));
    Odrv4 I__3928 (
            .O(N__17815),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__3927 (
            .O(N__17812),
            .I(\Lab_UT.di_ASones_1 ));
    Odrv4 I__3926 (
            .O(N__17809),
            .I(\Lab_UT.di_ASones_1 ));
    CascadeMux I__3925 (
            .O(N__17802),
            .I(N__17787));
    InMux I__3924 (
            .O(N__17801),
            .I(N__17775));
    InMux I__3923 (
            .O(N__17800),
            .I(N__17775));
    InMux I__3922 (
            .O(N__17799),
            .I(N__17775));
    InMux I__3921 (
            .O(N__17798),
            .I(N__17775));
    InMux I__3920 (
            .O(N__17797),
            .I(N__17775));
    InMux I__3919 (
            .O(N__17796),
            .I(N__17766));
    InMux I__3918 (
            .O(N__17795),
            .I(N__17766));
    InMux I__3917 (
            .O(N__17794),
            .I(N__17766));
    InMux I__3916 (
            .O(N__17793),
            .I(N__17757));
    InMux I__3915 (
            .O(N__17792),
            .I(N__17757));
    InMux I__3914 (
            .O(N__17791),
            .I(N__17757));
    InMux I__3913 (
            .O(N__17790),
            .I(N__17757));
    InMux I__3912 (
            .O(N__17787),
            .I(N__17752));
    InMux I__3911 (
            .O(N__17786),
            .I(N__17752));
    LocalMux I__3910 (
            .O(N__17775),
            .I(N__17749));
    InMux I__3909 (
            .O(N__17774),
            .I(N__17746));
    InMux I__3908 (
            .O(N__17773),
            .I(N__17743));
    LocalMux I__3907 (
            .O(N__17766),
            .I(N__17740));
    LocalMux I__3906 (
            .O(N__17757),
            .I(N__17733));
    LocalMux I__3905 (
            .O(N__17752),
            .I(N__17733));
    Span4Mux_s3_v I__3904 (
            .O(N__17749),
            .I(N__17733));
    LocalMux I__3903 (
            .O(N__17746),
            .I(\Lab_UT.loadalarm_0 ));
    LocalMux I__3902 (
            .O(N__17743),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv12 I__3901 (
            .O(N__17740),
            .I(\Lab_UT.loadalarm_0 ));
    Odrv4 I__3900 (
            .O(N__17733),
            .I(\Lab_UT.loadalarm_0 ));
    CascadeMux I__3899 (
            .O(N__17724),
            .I(N__17721));
    InMux I__3898 (
            .O(N__17721),
            .I(N__17713));
    InMux I__3897 (
            .O(N__17720),
            .I(N__17713));
    CascadeMux I__3896 (
            .O(N__17719),
            .I(N__17709));
    CascadeMux I__3895 (
            .O(N__17718),
            .I(N__17705));
    LocalMux I__3894 (
            .O(N__17713),
            .I(N__17701));
    InMux I__3893 (
            .O(N__17712),
            .I(N__17690));
    InMux I__3892 (
            .O(N__17709),
            .I(N__17690));
    InMux I__3891 (
            .O(N__17708),
            .I(N__17690));
    InMux I__3890 (
            .O(N__17705),
            .I(N__17690));
    InMux I__3889 (
            .O(N__17704),
            .I(N__17690));
    Span4Mux_h I__3888 (
            .O(N__17701),
            .I(N__17687));
    LocalMux I__3887 (
            .O(N__17690),
            .I(N__17684));
    Odrv4 I__3886 (
            .O(N__17687),
            .I(\Lab_UT.sec2_1 ));
    Odrv12 I__3885 (
            .O(N__17684),
            .I(\Lab_UT.sec2_1 ));
    InMux I__3884 (
            .O(N__17679),
            .I(N__17671));
    InMux I__3883 (
            .O(N__17678),
            .I(N__17666));
    InMux I__3882 (
            .O(N__17677),
            .I(N__17666));
    CascadeMux I__3881 (
            .O(N__17676),
            .I(N__17663));
    InMux I__3880 (
            .O(N__17675),
            .I(N__17658));
    InMux I__3879 (
            .O(N__17674),
            .I(N__17658));
    LocalMux I__3878 (
            .O(N__17671),
            .I(N__17653));
    LocalMux I__3877 (
            .O(N__17666),
            .I(N__17653));
    InMux I__3876 (
            .O(N__17663),
            .I(N__17650));
    LocalMux I__3875 (
            .O(N__17658),
            .I(N__17647));
    Span4Mux_v I__3874 (
            .O(N__17653),
            .I(N__17644));
    LocalMux I__3873 (
            .O(N__17650),
            .I(N__17641));
    Span4Mux_v I__3872 (
            .O(N__17647),
            .I(N__17638));
    Odrv4 I__3871 (
            .O(N__17644),
            .I(\Lab_UT.LdMtens ));
    Odrv4 I__3870 (
            .O(N__17641),
            .I(\Lab_UT.LdMtens ));
    Odrv4 I__3869 (
            .O(N__17638),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__3868 (
            .O(N__17631),
            .I(N__17628));
    InMux I__3867 (
            .O(N__17628),
            .I(N__17625));
    LocalMux I__3866 (
            .O(N__17625),
            .I(N__17622));
    Odrv4 I__3865 (
            .O(N__17622),
            .I(\Lab_UT.didp.countrce4.un13_qPone ));
    InMux I__3864 (
            .O(N__17619),
            .I(N__17615));
    InMux I__3863 (
            .O(N__17618),
            .I(N__17612));
    LocalMux I__3862 (
            .O(N__17615),
            .I(N__17604));
    LocalMux I__3861 (
            .O(N__17612),
            .I(N__17604));
    CascadeMux I__3860 (
            .O(N__17611),
            .I(N__17600));
    InMux I__3859 (
            .O(N__17610),
            .I(N__17595));
    InMux I__3858 (
            .O(N__17609),
            .I(N__17595));
    Span4Mux_h I__3857 (
            .O(N__17604),
            .I(N__17592));
    InMux I__3856 (
            .O(N__17603),
            .I(N__17587));
    InMux I__3855 (
            .O(N__17600),
            .I(N__17587));
    LocalMux I__3854 (
            .O(N__17595),
            .I(\Lab_UT.di_Mtens_2 ));
    Odrv4 I__3853 (
            .O(N__17592),
            .I(\Lab_UT.di_Mtens_2 ));
    LocalMux I__3852 (
            .O(N__17587),
            .I(\Lab_UT.di_Mtens_2 ));
    CascadeMux I__3851 (
            .O(N__17580),
            .I(N__17577));
    InMux I__3850 (
            .O(N__17577),
            .I(N__17574));
    LocalMux I__3849 (
            .O(N__17574),
            .I(\Lab_UT.didp.countrce4.q_5_2 ));
    CascadeMux I__3848 (
            .O(N__17571),
            .I(N__17568));
    InMux I__3847 (
            .O(N__17568),
            .I(N__17565));
    LocalMux I__3846 (
            .O(N__17565),
            .I(N__17562));
    Span4Mux_v I__3845 (
            .O(N__17562),
            .I(N__17559));
    Span4Mux_h I__3844 (
            .O(N__17559),
            .I(N__17555));
    InMux I__3843 (
            .O(N__17558),
            .I(N__17552));
    Odrv4 I__3842 (
            .O(N__17555),
            .I(uu0_sec_clkD));
    LocalMux I__3841 (
            .O(N__17552),
            .I(uu0_sec_clkD));
    InMux I__3840 (
            .O(N__17547),
            .I(N__17543));
    InMux I__3839 (
            .O(N__17546),
            .I(N__17539));
    LocalMux I__3838 (
            .O(N__17543),
            .I(N__17536));
    InMux I__3837 (
            .O(N__17542),
            .I(N__17532));
    LocalMux I__3836 (
            .O(N__17539),
            .I(N__17529));
    Span4Mux_s2_v I__3835 (
            .O(N__17536),
            .I(N__17526));
    InMux I__3834 (
            .O(N__17535),
            .I(N__17523));
    LocalMux I__3833 (
            .O(N__17532),
            .I(N__17520));
    Span4Mux_v I__3832 (
            .O(N__17529),
            .I(N__17513));
    Span4Mux_v I__3831 (
            .O(N__17526),
            .I(N__17513));
    LocalMux I__3830 (
            .O(N__17523),
            .I(N__17513));
    Span4Mux_v I__3829 (
            .O(N__17520),
            .I(N__17507));
    Span4Mux_h I__3828 (
            .O(N__17513),
            .I(N__17507));
    InMux I__3827 (
            .O(N__17512),
            .I(N__17504));
    Span4Mux_h I__3826 (
            .O(N__17507),
            .I(N__17501));
    LocalMux I__3825 (
            .O(N__17504),
            .I(o_One_Sec_Pulse));
    Odrv4 I__3824 (
            .O(N__17501),
            .I(o_One_Sec_Pulse));
    CascadeMux I__3823 (
            .O(N__17496),
            .I(N__17488));
    CascadeMux I__3822 (
            .O(N__17495),
            .I(N__17484));
    CascadeMux I__3821 (
            .O(N__17494),
            .I(N__17481));
    CascadeMux I__3820 (
            .O(N__17493),
            .I(N__17477));
    InMux I__3819 (
            .O(N__17492),
            .I(N__17472));
    InMux I__3818 (
            .O(N__17491),
            .I(N__17472));
    InMux I__3817 (
            .O(N__17488),
            .I(N__17465));
    InMux I__3816 (
            .O(N__17487),
            .I(N__17465));
    InMux I__3815 (
            .O(N__17484),
            .I(N__17465));
    InMux I__3814 (
            .O(N__17481),
            .I(N__17462));
    CascadeMux I__3813 (
            .O(N__17480),
            .I(N__17459));
    InMux I__3812 (
            .O(N__17477),
            .I(N__17456));
    LocalMux I__3811 (
            .O(N__17472),
            .I(N__17449));
    LocalMux I__3810 (
            .O(N__17465),
            .I(N__17449));
    LocalMux I__3809 (
            .O(N__17462),
            .I(N__17449));
    InMux I__3808 (
            .O(N__17459),
            .I(N__17446));
    LocalMux I__3807 (
            .O(N__17456),
            .I(N__17443));
    Span4Mux_v I__3806 (
            .O(N__17449),
            .I(N__17438));
    LocalMux I__3805 (
            .O(N__17446),
            .I(N__17438));
    Odrv12 I__3804 (
            .O(N__17443),
            .I(oneSecStrb));
    Odrv4 I__3803 (
            .O(N__17438),
            .I(oneSecStrb));
    CascadeMux I__3802 (
            .O(N__17433),
            .I(oneSecStrb_cascade_));
    CascadeMux I__3801 (
            .O(N__17430),
            .I(N__17426));
    InMux I__3800 (
            .O(N__17429),
            .I(N__17423));
    InMux I__3799 (
            .O(N__17426),
            .I(N__17420));
    LocalMux I__3798 (
            .O(N__17423),
            .I(N__17417));
    LocalMux I__3797 (
            .O(N__17420),
            .I(N__17414));
    Span4Mux_h I__3796 (
            .O(N__17417),
            .I(N__17411));
    Span4Mux_h I__3795 (
            .O(N__17414),
            .I(N__17408));
    Odrv4 I__3794 (
            .O(N__17411),
            .I(\Lab_UT.dispString.N_102 ));
    Odrv4 I__3793 (
            .O(N__17408),
            .I(\Lab_UT.dispString.N_102 ));
    InMux I__3792 (
            .O(N__17403),
            .I(N__17400));
    LocalMux I__3791 (
            .O(N__17400),
            .I(N__17396));
    InMux I__3790 (
            .O(N__17399),
            .I(N__17393));
    Span4Mux_v I__3789 (
            .O(N__17396),
            .I(N__17390));
    LocalMux I__3788 (
            .O(N__17393),
            .I(N__17387));
    Span4Mux_h I__3787 (
            .O(N__17390),
            .I(N__17384));
    Span4Mux_h I__3786 (
            .O(N__17387),
            .I(N__17381));
    Odrv4 I__3785 (
            .O(N__17384),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    Odrv4 I__3784 (
            .O(N__17381),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__3783 (
            .O(N__17376),
            .I(N__17373));
    LocalMux I__3782 (
            .O(N__17373),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    CascadeMux I__3781 (
            .O(N__17370),
            .I(N__17366));
    CascadeMux I__3780 (
            .O(N__17369),
            .I(N__17363));
    InMux I__3779 (
            .O(N__17366),
            .I(N__17360));
    InMux I__3778 (
            .O(N__17363),
            .I(N__17355));
    LocalMux I__3777 (
            .O(N__17360),
            .I(N__17352));
    InMux I__3776 (
            .O(N__17359),
            .I(N__17349));
    InMux I__3775 (
            .O(N__17358),
            .I(N__17346));
    LocalMux I__3774 (
            .O(N__17355),
            .I(N__17343));
    Span4Mux_v I__3773 (
            .O(N__17352),
            .I(N__17334));
    LocalMux I__3772 (
            .O(N__17349),
            .I(N__17334));
    LocalMux I__3771 (
            .O(N__17346),
            .I(N__17334));
    Span4Mux_v I__3770 (
            .O(N__17343),
            .I(N__17334));
    Odrv4 I__3769 (
            .O(N__17334),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    InMux I__3768 (
            .O(N__17331),
            .I(N__17325));
    InMux I__3767 (
            .O(N__17330),
            .I(N__17318));
    InMux I__3766 (
            .O(N__17329),
            .I(N__17318));
    InMux I__3765 (
            .O(N__17328),
            .I(N__17318));
    LocalMux I__3764 (
            .O(N__17325),
            .I(N__17311));
    LocalMux I__3763 (
            .O(N__17318),
            .I(N__17311));
    InMux I__3762 (
            .O(N__17317),
            .I(N__17306));
    InMux I__3761 (
            .O(N__17316),
            .I(N__17306));
    Odrv4 I__3760 (
            .O(N__17311),
            .I(\Lab_UT.LdMones ));
    LocalMux I__3759 (
            .O(N__17306),
            .I(\Lab_UT.LdMones ));
    InMux I__3758 (
            .O(N__17301),
            .I(N__17295));
    InMux I__3757 (
            .O(N__17300),
            .I(N__17289));
    InMux I__3756 (
            .O(N__17299),
            .I(N__17284));
    InMux I__3755 (
            .O(N__17298),
            .I(N__17284));
    LocalMux I__3754 (
            .O(N__17295),
            .I(N__17281));
    InMux I__3753 (
            .O(N__17294),
            .I(N__17278));
    InMux I__3752 (
            .O(N__17293),
            .I(N__17273));
    InMux I__3751 (
            .O(N__17292),
            .I(N__17273));
    LocalMux I__3750 (
            .O(N__17289),
            .I(N__17268));
    LocalMux I__3749 (
            .O(N__17284),
            .I(N__17268));
    Span4Mux_h I__3748 (
            .O(N__17281),
            .I(N__17265));
    LocalMux I__3747 (
            .O(N__17278),
            .I(N__17262));
    LocalMux I__3746 (
            .O(N__17273),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__3745 (
            .O(N__17268),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv4 I__3744 (
            .O(N__17265),
            .I(\Lab_UT.di_Mones_0 ));
    Odrv12 I__3743 (
            .O(N__17262),
            .I(\Lab_UT.di_Mones_0 ));
    CascadeMux I__3742 (
            .O(N__17253),
            .I(N__17249));
    CascadeMux I__3741 (
            .O(N__17252),
            .I(N__17244));
    InMux I__3740 (
            .O(N__17249),
            .I(N__17240));
    CascadeMux I__3739 (
            .O(N__17248),
            .I(N__17235));
    CascadeMux I__3738 (
            .O(N__17247),
            .I(N__17232));
    InMux I__3737 (
            .O(N__17244),
            .I(N__17228));
    InMux I__3736 (
            .O(N__17243),
            .I(N__17225));
    LocalMux I__3735 (
            .O(N__17240),
            .I(N__17222));
    InMux I__3734 (
            .O(N__17239),
            .I(N__17219));
    InMux I__3733 (
            .O(N__17238),
            .I(N__17216));
    InMux I__3732 (
            .O(N__17235),
            .I(N__17213));
    InMux I__3731 (
            .O(N__17232),
            .I(N__17208));
    InMux I__3730 (
            .O(N__17231),
            .I(N__17208));
    LocalMux I__3729 (
            .O(N__17228),
            .I(N__17205));
    LocalMux I__3728 (
            .O(N__17225),
            .I(N__17192));
    Span4Mux_h I__3727 (
            .O(N__17222),
            .I(N__17192));
    LocalMux I__3726 (
            .O(N__17219),
            .I(N__17192));
    LocalMux I__3725 (
            .O(N__17216),
            .I(N__17192));
    LocalMux I__3724 (
            .O(N__17213),
            .I(N__17192));
    LocalMux I__3723 (
            .O(N__17208),
            .I(N__17192));
    Span4Mux_v I__3722 (
            .O(N__17205),
            .I(N__17187));
    Span4Mux_v I__3721 (
            .O(N__17192),
            .I(N__17187));
    Odrv4 I__3720 (
            .O(N__17187),
            .I(\Lab_UT.dictrl.state_i_3_0 ));
    InMux I__3719 (
            .O(N__17184),
            .I(N__17181));
    LocalMux I__3718 (
            .O(N__17181),
            .I(N__17178));
    Sp12to4 I__3717 (
            .O(N__17178),
            .I(N__17175));
    Odrv12 I__3716 (
            .O(N__17175),
            .I(\Lab_UT.dictrl.state_ret_2_fast ));
    InMux I__3715 (
            .O(N__17172),
            .I(N__17169));
    LocalMux I__3714 (
            .O(N__17169),
            .I(N__17165));
    CascadeMux I__3713 (
            .O(N__17168),
            .I(N__17161));
    Span4Mux_s3_h I__3712 (
            .O(N__17165),
            .I(N__17158));
    InMux I__3711 (
            .O(N__17164),
            .I(N__17155));
    InMux I__3710 (
            .O(N__17161),
            .I(N__17152));
    Odrv4 I__3709 (
            .O(N__17158),
            .I(\Lab_UT.dictrl.N_20 ));
    LocalMux I__3708 (
            .O(N__17155),
            .I(\Lab_UT.dictrl.N_20 ));
    LocalMux I__3707 (
            .O(N__17152),
            .I(\Lab_UT.dictrl.N_20 ));
    InMux I__3706 (
            .O(N__17145),
            .I(N__17142));
    LocalMux I__3705 (
            .O(N__17142),
            .I(N__17137));
    InMux I__3704 (
            .O(N__17141),
            .I(N__17134));
    InMux I__3703 (
            .O(N__17140),
            .I(N__17131));
    Odrv4 I__3702 (
            .O(N__17137),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    LocalMux I__3701 (
            .O(N__17134),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    LocalMux I__3700 (
            .O(N__17131),
            .I(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ));
    InMux I__3699 (
            .O(N__17124),
            .I(N__17119));
    InMux I__3698 (
            .O(N__17123),
            .I(N__17114));
    InMux I__3697 (
            .O(N__17122),
            .I(N__17114));
    LocalMux I__3696 (
            .O(N__17119),
            .I(N__17111));
    LocalMux I__3695 (
            .O(N__17114),
            .I(N__17108));
    Odrv4 I__3694 (
            .O(N__17111),
            .I(\Lab_UT.dispString.N_144 ));
    Odrv12 I__3693 (
            .O(N__17108),
            .I(\Lab_UT.dispString.N_144 ));
    InMux I__3692 (
            .O(N__17103),
            .I(N__17097));
    InMux I__3691 (
            .O(N__17102),
            .I(N__17094));
    InMux I__3690 (
            .O(N__17101),
            .I(N__17091));
    InMux I__3689 (
            .O(N__17100),
            .I(N__17088));
    LocalMux I__3688 (
            .O(N__17097),
            .I(N__17084));
    LocalMux I__3687 (
            .O(N__17094),
            .I(N__17078));
    LocalMux I__3686 (
            .O(N__17091),
            .I(N__17078));
    LocalMux I__3685 (
            .O(N__17088),
            .I(N__17074));
    CascadeMux I__3684 (
            .O(N__17087),
            .I(N__17071));
    Span4Mux_h I__3683 (
            .O(N__17084),
            .I(N__17068));
    InMux I__3682 (
            .O(N__17083),
            .I(N__17065));
    Span4Mux_h I__3681 (
            .O(N__17078),
            .I(N__17062));
    InMux I__3680 (
            .O(N__17077),
            .I(N__17059));
    Span12Mux_s6_h I__3679 (
            .O(N__17074),
            .I(N__17056));
    InMux I__3678 (
            .O(N__17071),
            .I(N__17053));
    Odrv4 I__3677 (
            .O(N__17068),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3676 (
            .O(N__17065),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv4 I__3675 (
            .O(N__17062),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3674 (
            .O(N__17059),
            .I(\Lab_UT.di_Mtens_0 ));
    Odrv12 I__3673 (
            .O(N__17056),
            .I(\Lab_UT.di_Mtens_0 ));
    LocalMux I__3672 (
            .O(N__17053),
            .I(\Lab_UT.di_Mtens_0 ));
    CascadeMux I__3671 (
            .O(N__17040),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__3670 (
            .O(N__17037),
            .I(N__17033));
    InMux I__3669 (
            .O(N__17036),
            .I(N__17030));
    LocalMux I__3668 (
            .O(N__17033),
            .I(N__17022));
    LocalMux I__3667 (
            .O(N__17030),
            .I(N__17019));
    InMux I__3666 (
            .O(N__17029),
            .I(N__17016));
    InMux I__3665 (
            .O(N__17028),
            .I(N__17013));
    InMux I__3664 (
            .O(N__17027),
            .I(N__17008));
    InMux I__3663 (
            .O(N__17026),
            .I(N__17008));
    InMux I__3662 (
            .O(N__17025),
            .I(N__17005));
    Span4Mux_v I__3661 (
            .O(N__17022),
            .I(N__16998));
    Span4Mux_v I__3660 (
            .O(N__17019),
            .I(N__16998));
    LocalMux I__3659 (
            .O(N__17016),
            .I(N__16998));
    LocalMux I__3658 (
            .O(N__17013),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__3657 (
            .O(N__17008),
            .I(\Lab_UT.di_Mtens_1 ));
    LocalMux I__3656 (
            .O(N__17005),
            .I(\Lab_UT.di_Mtens_1 ));
    Odrv4 I__3655 (
            .O(N__16998),
            .I(\Lab_UT.di_Mtens_1 ));
    InMux I__3654 (
            .O(N__16989),
            .I(N__16986));
    LocalMux I__3653 (
            .O(N__16986),
            .I(N__16980));
    CascadeMux I__3652 (
            .O(N__16985),
            .I(N__16975));
    InMux I__3651 (
            .O(N__16984),
            .I(N__16970));
    InMux I__3650 (
            .O(N__16983),
            .I(N__16970));
    Span4Mux_v I__3649 (
            .O(N__16980),
            .I(N__16967));
    InMux I__3648 (
            .O(N__16979),
            .I(N__16964));
    InMux I__3647 (
            .O(N__16978),
            .I(N__16961));
    InMux I__3646 (
            .O(N__16975),
            .I(N__16958));
    LocalMux I__3645 (
            .O(N__16970),
            .I(\Lab_UT.di_Sones_2 ));
    Odrv4 I__3644 (
            .O(N__16967),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3643 (
            .O(N__16964),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3642 (
            .O(N__16961),
            .I(\Lab_UT.di_Sones_2 ));
    LocalMux I__3641 (
            .O(N__16958),
            .I(\Lab_UT.di_Sones_2 ));
    InMux I__3640 (
            .O(N__16947),
            .I(N__16944));
    LocalMux I__3639 (
            .O(N__16944),
            .I(N__16939));
    InMux I__3638 (
            .O(N__16943),
            .I(N__16936));
    InMux I__3637 (
            .O(N__16942),
            .I(N__16933));
    Span4Mux_h I__3636 (
            .O(N__16939),
            .I(N__16930));
    LocalMux I__3635 (
            .O(N__16936),
            .I(N__16927));
    LocalMux I__3634 (
            .O(N__16933),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__3633 (
            .O(N__16930),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__3632 (
            .O(N__16927),
            .I(\Lab_UT.di_ASones_2 ));
    InMux I__3631 (
            .O(N__16920),
            .I(N__16914));
    InMux I__3630 (
            .O(N__16919),
            .I(N__16914));
    LocalMux I__3629 (
            .O(N__16914),
            .I(N__16906));
    InMux I__3628 (
            .O(N__16913),
            .I(N__16895));
    InMux I__3627 (
            .O(N__16912),
            .I(N__16895));
    InMux I__3626 (
            .O(N__16911),
            .I(N__16895));
    InMux I__3625 (
            .O(N__16910),
            .I(N__16895));
    InMux I__3624 (
            .O(N__16909),
            .I(N__16895));
    Span4Mux_h I__3623 (
            .O(N__16906),
            .I(N__16892));
    LocalMux I__3622 (
            .O(N__16895),
            .I(N__16889));
    Odrv4 I__3621 (
            .O(N__16892),
            .I(\Lab_UT.sec2_2 ));
    Odrv12 I__3620 (
            .O(N__16889),
            .I(\Lab_UT.sec2_2 ));
    InMux I__3619 (
            .O(N__16884),
            .I(N__16875));
    InMux I__3618 (
            .O(N__16883),
            .I(N__16868));
    InMux I__3617 (
            .O(N__16882),
            .I(N__16868));
    InMux I__3616 (
            .O(N__16881),
            .I(N__16868));
    InMux I__3615 (
            .O(N__16880),
            .I(N__16865));
    InMux I__3614 (
            .O(N__16879),
            .I(N__16860));
    InMux I__3613 (
            .O(N__16878),
            .I(N__16860));
    LocalMux I__3612 (
            .O(N__16875),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3611 (
            .O(N__16868),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3610 (
            .O(N__16865),
            .I(\Lab_UT.di_Mones_1 ));
    LocalMux I__3609 (
            .O(N__16860),
            .I(\Lab_UT.di_Mones_1 ));
    InMux I__3608 (
            .O(N__16851),
            .I(N__16848));
    LocalMux I__3607 (
            .O(N__16848),
            .I(N__16845));
    Odrv4 I__3606 (
            .O(N__16845),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    InMux I__3605 (
            .O(N__16842),
            .I(N__16839));
    LocalMux I__3604 (
            .O(N__16839),
            .I(N__16835));
    InMux I__3603 (
            .O(N__16838),
            .I(N__16832));
    Span4Mux_v I__3602 (
            .O(N__16835),
            .I(N__16825));
    LocalMux I__3601 (
            .O(N__16832),
            .I(N__16825));
    InMux I__3600 (
            .O(N__16831),
            .I(N__16820));
    InMux I__3599 (
            .O(N__16830),
            .I(N__16820));
    Span4Mux_h I__3598 (
            .O(N__16825),
            .I(N__16817));
    LocalMux I__3597 (
            .O(N__16820),
            .I(N__16814));
    Odrv4 I__3596 (
            .O(N__16817),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    Odrv12 I__3595 (
            .O(N__16814),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    InMux I__3594 (
            .O(N__16809),
            .I(N__16805));
    InMux I__3593 (
            .O(N__16808),
            .I(N__16802));
    LocalMux I__3592 (
            .O(N__16805),
            .I(N__16799));
    LocalMux I__3591 (
            .O(N__16802),
            .I(N__16796));
    Span4Mux_h I__3590 (
            .O(N__16799),
            .I(N__16793));
    Odrv12 I__3589 (
            .O(N__16796),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    Odrv4 I__3588 (
            .O(N__16793),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    InMux I__3587 (
            .O(N__16788),
            .I(N__16785));
    LocalMux I__3586 (
            .O(N__16785),
            .I(N__16782));
    Span4Mux_h I__3585 (
            .O(N__16782),
            .I(N__16777));
    InMux I__3584 (
            .O(N__16781),
            .I(N__16774));
    InMux I__3583 (
            .O(N__16780),
            .I(N__16771));
    Odrv4 I__3582 (
            .O(N__16777),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    LocalMux I__3581 (
            .O(N__16774),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    LocalMux I__3580 (
            .O(N__16771),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    CascadeMux I__3579 (
            .O(N__16764),
            .I(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ));
    CascadeMux I__3578 (
            .O(N__16761),
            .I(\Lab_UT.didp.countrce3.q_5_2_cascade_ ));
    InMux I__3577 (
            .O(N__16758),
            .I(N__16755));
    LocalMux I__3576 (
            .O(N__16755),
            .I(N__16752));
    Odrv4 I__3575 (
            .O(N__16752),
            .I(\Lab_UT.didp.reset_12_1_3 ));
    InMux I__3574 (
            .O(N__16749),
            .I(N__16744));
    InMux I__3573 (
            .O(N__16748),
            .I(N__16738));
    InMux I__3572 (
            .O(N__16747),
            .I(N__16735));
    LocalMux I__3571 (
            .O(N__16744),
            .I(N__16732));
    InMux I__3570 (
            .O(N__16743),
            .I(N__16725));
    InMux I__3569 (
            .O(N__16742),
            .I(N__16725));
    InMux I__3568 (
            .O(N__16741),
            .I(N__16725));
    LocalMux I__3567 (
            .O(N__16738),
            .I(N__16720));
    LocalMux I__3566 (
            .O(N__16735),
            .I(N__16720));
    Span4Mux_h I__3565 (
            .O(N__16732),
            .I(N__16717));
    LocalMux I__3564 (
            .O(N__16725),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3563 (
            .O(N__16720),
            .I(\Lab_UT.di_Mones_2 ));
    Odrv4 I__3562 (
            .O(N__16717),
            .I(\Lab_UT.di_Mones_2 ));
    CascadeMux I__3561 (
            .O(N__16710),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    InMux I__3560 (
            .O(N__16707),
            .I(N__16703));
    CascadeMux I__3559 (
            .O(N__16706),
            .I(N__16698));
    LocalMux I__3558 (
            .O(N__16703),
            .I(N__16694));
    InMux I__3557 (
            .O(N__16702),
            .I(N__16691));
    InMux I__3556 (
            .O(N__16701),
            .I(N__16688));
    InMux I__3555 (
            .O(N__16698),
            .I(N__16685));
    InMux I__3554 (
            .O(N__16697),
            .I(N__16682));
    Span12Mux_v I__3553 (
            .O(N__16694),
            .I(N__16679));
    LocalMux I__3552 (
            .O(N__16691),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3551 (
            .O(N__16688),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3550 (
            .O(N__16685),
            .I(\Lab_UT.di_Mones_3 ));
    LocalMux I__3549 (
            .O(N__16682),
            .I(\Lab_UT.di_Mones_3 ));
    Odrv12 I__3548 (
            .O(N__16679),
            .I(\Lab_UT.di_Mones_3 ));
    InMux I__3547 (
            .O(N__16668),
            .I(N__16665));
    LocalMux I__3546 (
            .O(N__16665),
            .I(\Lab_UT.didp.countrce3.q_5_3 ));
    InMux I__3545 (
            .O(N__16662),
            .I(N__16658));
    InMux I__3544 (
            .O(N__16661),
            .I(N__16655));
    LocalMux I__3543 (
            .O(N__16658),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    LocalMux I__3542 (
            .O(N__16655),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    CascadeMux I__3541 (
            .O(N__16650),
            .I(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ));
    InMux I__3540 (
            .O(N__16647),
            .I(N__16644));
    LocalMux I__3539 (
            .O(N__16644),
            .I(N__16641));
    Span4Mux_s1_v I__3538 (
            .O(N__16641),
            .I(N__16638));
    Odrv4 I__3537 (
            .O(N__16638),
            .I(\uu2.bitmapZ0Z_111 ));
    InMux I__3536 (
            .O(N__16635),
            .I(N__16624));
    InMux I__3535 (
            .O(N__16634),
            .I(N__16624));
    InMux I__3534 (
            .O(N__16633),
            .I(N__16624));
    InMux I__3533 (
            .O(N__16632),
            .I(N__16618));
    InMux I__3532 (
            .O(N__16631),
            .I(N__16618));
    LocalMux I__3531 (
            .O(N__16624),
            .I(N__16613));
    InMux I__3530 (
            .O(N__16623),
            .I(N__16610));
    LocalMux I__3529 (
            .O(N__16618),
            .I(N__16607));
    CascadeMux I__3528 (
            .O(N__16617),
            .I(N__16604));
    InMux I__3527 (
            .O(N__16616),
            .I(N__16598));
    Span4Mux_s1_v I__3526 (
            .O(N__16613),
            .I(N__16595));
    LocalMux I__3525 (
            .O(N__16610),
            .I(N__16592));
    Span4Mux_h I__3524 (
            .O(N__16607),
            .I(N__16589));
    InMux I__3523 (
            .O(N__16604),
            .I(N__16584));
    InMux I__3522 (
            .O(N__16603),
            .I(N__16584));
    InMux I__3521 (
            .O(N__16602),
            .I(N__16581));
    InMux I__3520 (
            .O(N__16601),
            .I(N__16578));
    LocalMux I__3519 (
            .O(N__16598),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3518 (
            .O(N__16595),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv12 I__3517 (
            .O(N__16592),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__3516 (
            .O(N__16589),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3515 (
            .O(N__16584),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3514 (
            .O(N__16581),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__3513 (
            .O(N__16578),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__3512 (
            .O(N__16563),
            .I(N__16560));
    LocalMux I__3511 (
            .O(N__16560),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__3510 (
            .O(N__16557),
            .I(N__16545));
    InMux I__3509 (
            .O(N__16556),
            .I(N__16545));
    InMux I__3508 (
            .O(N__16555),
            .I(N__16545));
    InMux I__3507 (
            .O(N__16554),
            .I(N__16545));
    LocalMux I__3506 (
            .O(N__16545),
            .I(N__16537));
    InMux I__3505 (
            .O(N__16544),
            .I(N__16530));
    InMux I__3504 (
            .O(N__16543),
            .I(N__16530));
    InMux I__3503 (
            .O(N__16542),
            .I(N__16530));
    CascadeMux I__3502 (
            .O(N__16541),
            .I(N__16526));
    CascadeMux I__3501 (
            .O(N__16540),
            .I(N__16523));
    Span4Mux_s2_v I__3500 (
            .O(N__16537),
            .I(N__16518));
    LocalMux I__3499 (
            .O(N__16530),
            .I(N__16518));
    InMux I__3498 (
            .O(N__16529),
            .I(N__16515));
    InMux I__3497 (
            .O(N__16526),
            .I(N__16512));
    InMux I__3496 (
            .O(N__16523),
            .I(N__16509));
    Span4Mux_h I__3495 (
            .O(N__16518),
            .I(N__16506));
    LocalMux I__3494 (
            .O(N__16515),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3493 (
            .O(N__16512),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    LocalMux I__3492 (
            .O(N__16509),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    Odrv4 I__3491 (
            .O(N__16506),
            .I(\uu2.w_addr_displaying_0_repZ0Z1 ));
    InMux I__3490 (
            .O(N__16497),
            .I(N__16494));
    LocalMux I__3489 (
            .O(N__16494),
            .I(\uu2.bitmapZ0Z_90 ));
    InMux I__3488 (
            .O(N__16491),
            .I(N__16488));
    LocalMux I__3487 (
            .O(N__16488),
            .I(N__16485));
    Odrv4 I__3486 (
            .O(N__16485),
            .I(\uu2.bitmap_pmux_19_ns_1 ));
    InMux I__3485 (
            .O(N__16482),
            .I(N__16476));
    InMux I__3484 (
            .O(N__16481),
            .I(N__16476));
    LocalMux I__3483 (
            .O(N__16476),
            .I(N__16468));
    InMux I__3482 (
            .O(N__16475),
            .I(N__16457));
    InMux I__3481 (
            .O(N__16474),
            .I(N__16457));
    InMux I__3480 (
            .O(N__16473),
            .I(N__16457));
    InMux I__3479 (
            .O(N__16472),
            .I(N__16457));
    InMux I__3478 (
            .O(N__16471),
            .I(N__16457));
    Odrv4 I__3477 (
            .O(N__16468),
            .I(\Lab_UT.sec2_0 ));
    LocalMux I__3476 (
            .O(N__16457),
            .I(\Lab_UT.sec2_0 ));
    CascadeMux I__3475 (
            .O(N__16452),
            .I(N__16448));
    InMux I__3474 (
            .O(N__16451),
            .I(N__16440));
    InMux I__3473 (
            .O(N__16448),
            .I(N__16440));
    CascadeMux I__3472 (
            .O(N__16447),
            .I(N__16437));
    CascadeMux I__3471 (
            .O(N__16446),
            .I(N__16433));
    CascadeMux I__3470 (
            .O(N__16445),
            .I(N__16429));
    LocalMux I__3469 (
            .O(N__16440),
            .I(N__16426));
    InMux I__3468 (
            .O(N__16437),
            .I(N__16415));
    InMux I__3467 (
            .O(N__16436),
            .I(N__16415));
    InMux I__3466 (
            .O(N__16433),
            .I(N__16415));
    InMux I__3465 (
            .O(N__16432),
            .I(N__16415));
    InMux I__3464 (
            .O(N__16429),
            .I(N__16415));
    Span4Mux_s2_v I__3463 (
            .O(N__16426),
            .I(N__16410));
    LocalMux I__3462 (
            .O(N__16415),
            .I(N__16410));
    Odrv4 I__3461 (
            .O(N__16410),
            .I(\Lab_UT.sec2_3 ));
    InMux I__3460 (
            .O(N__16407),
            .I(N__16400));
    InMux I__3459 (
            .O(N__16406),
            .I(N__16393));
    InMux I__3458 (
            .O(N__16405),
            .I(N__16393));
    InMux I__3457 (
            .O(N__16404),
            .I(N__16393));
    InMux I__3456 (
            .O(N__16403),
            .I(N__16390));
    LocalMux I__3455 (
            .O(N__16400),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3454 (
            .O(N__16393),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__3453 (
            .O(N__16390),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    InMux I__3452 (
            .O(N__16383),
            .I(N__16380));
    LocalMux I__3451 (
            .O(N__16380),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__3450 (
            .O(N__16377),
            .I(N__16374));
    LocalMux I__3449 (
            .O(N__16374),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__3448 (
            .O(N__16371),
            .I(N__16367));
    InMux I__3447 (
            .O(N__16370),
            .I(N__16364));
    LocalMux I__3446 (
            .O(N__16367),
            .I(N__16361));
    LocalMux I__3445 (
            .O(N__16364),
            .I(\uu2.bitmapZ0Z_314 ));
    Odrv12 I__3444 (
            .O(N__16361),
            .I(\uu2.bitmapZ0Z_314 ));
    CascadeMux I__3443 (
            .O(N__16356),
            .I(\uu2.N_152_cascade_ ));
    CascadeMux I__3442 (
            .O(N__16353),
            .I(N__16350));
    InMux I__3441 (
            .O(N__16350),
            .I(N__16344));
    InMux I__3440 (
            .O(N__16349),
            .I(N__16341));
    CascadeMux I__3439 (
            .O(N__16348),
            .I(N__16338));
    InMux I__3438 (
            .O(N__16347),
            .I(N__16335));
    LocalMux I__3437 (
            .O(N__16344),
            .I(N__16330));
    LocalMux I__3436 (
            .O(N__16341),
            .I(N__16330));
    InMux I__3435 (
            .O(N__16338),
            .I(N__16327));
    LocalMux I__3434 (
            .O(N__16335),
            .I(N__16324));
    Span4Mux_v I__3433 (
            .O(N__16330),
            .I(N__16321));
    LocalMux I__3432 (
            .O(N__16327),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__3431 (
            .O(N__16324),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    Odrv4 I__3430 (
            .O(N__16321),
            .I(\uu2.w_addr_displaying_fastZ0Z_8 ));
    InMux I__3429 (
            .O(N__16314),
            .I(N__16308));
    InMux I__3428 (
            .O(N__16313),
            .I(N__16308));
    LocalMux I__3427 (
            .O(N__16308),
            .I(N__16305));
    Span4Mux_h I__3426 (
            .O(N__16305),
            .I(N__16302));
    Odrv4 I__3425 (
            .O(N__16302),
            .I(\uu2.bitmap_RNIM5E21Z0Z_314 ));
    InMux I__3424 (
            .O(N__16299),
            .I(N__16296));
    LocalMux I__3423 (
            .O(N__16296),
            .I(N__16291));
    InMux I__3422 (
            .O(N__16295),
            .I(N__16284));
    InMux I__3421 (
            .O(N__16294),
            .I(N__16284));
    Span4Mux_s0_v I__3420 (
            .O(N__16291),
            .I(N__16281));
    InMux I__3419 (
            .O(N__16290),
            .I(N__16276));
    InMux I__3418 (
            .O(N__16289),
            .I(N__16276));
    LocalMux I__3417 (
            .O(N__16284),
            .I(\uu2.w_addr_userZ0Z_4 ));
    Odrv4 I__3416 (
            .O(N__16281),
            .I(\uu2.w_addr_userZ0Z_4 ));
    LocalMux I__3415 (
            .O(N__16276),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__3414 (
            .O(N__16269),
            .I(\uu2.un3_w_addr_user_4_cascade_ ));
    InMux I__3413 (
            .O(N__16266),
            .I(N__16263));
    LocalMux I__3412 (
            .O(N__16263),
            .I(\uu2.un3_w_addr_user_5 ));
    InMux I__3411 (
            .O(N__16260),
            .I(N__16254));
    InMux I__3410 (
            .O(N__16259),
            .I(N__16254));
    LocalMux I__3409 (
            .O(N__16254),
            .I(N__16251));
    Span4Mux_h I__3408 (
            .O(N__16251),
            .I(N__16248));
    Odrv4 I__3407 (
            .O(N__16248),
            .I(\uu2.un3_w_addr_user ));
    InMux I__3406 (
            .O(N__16245),
            .I(N__16242));
    LocalMux I__3405 (
            .O(N__16242),
            .I(N__16239));
    Span4Mux_h I__3404 (
            .O(N__16239),
            .I(N__16235));
    CascadeMux I__3403 (
            .O(N__16238),
            .I(N__16228));
    Span4Mux_v I__3402 (
            .O(N__16235),
            .I(N__16224));
    InMux I__3401 (
            .O(N__16234),
            .I(N__16217));
    InMux I__3400 (
            .O(N__16233),
            .I(N__16217));
    InMux I__3399 (
            .O(N__16232),
            .I(N__16217));
    InMux I__3398 (
            .O(N__16231),
            .I(N__16210));
    InMux I__3397 (
            .O(N__16228),
            .I(N__16210));
    InMux I__3396 (
            .O(N__16227),
            .I(N__16210));
    Span4Mux_v I__3395 (
            .O(N__16224),
            .I(N__16207));
    LocalMux I__3394 (
            .O(N__16217),
            .I(N__16204));
    LocalMux I__3393 (
            .O(N__16210),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__3392 (
            .O(N__16207),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__3391 (
            .O(N__16204),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__3390 (
            .O(N__16197),
            .I(\uu2.un404_ci_cascade_ ));
    InMux I__3389 (
            .O(N__16194),
            .I(N__16188));
    InMux I__3388 (
            .O(N__16193),
            .I(N__16185));
    InMux I__3387 (
            .O(N__16192),
            .I(N__16182));
    InMux I__3386 (
            .O(N__16191),
            .I(N__16178));
    LocalMux I__3385 (
            .O(N__16188),
            .I(N__16171));
    LocalMux I__3384 (
            .O(N__16185),
            .I(N__16171));
    LocalMux I__3383 (
            .O(N__16182),
            .I(N__16171));
    InMux I__3382 (
            .O(N__16181),
            .I(N__16168));
    LocalMux I__3381 (
            .O(N__16178),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv12 I__3380 (
            .O(N__16171),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__3379 (
            .O(N__16168),
            .I(\uu2.w_addr_userZ0Z_6 ));
    InMux I__3378 (
            .O(N__16161),
            .I(N__16155));
    InMux I__3377 (
            .O(N__16160),
            .I(N__16155));
    LocalMux I__3376 (
            .O(N__16155),
            .I(N__16150));
    InMux I__3375 (
            .O(N__16154),
            .I(N__16145));
    InMux I__3374 (
            .O(N__16153),
            .I(N__16145));
    Odrv4 I__3373 (
            .O(N__16150),
            .I(\uu2.w_addr_userZ0Z_7 ));
    LocalMux I__3372 (
            .O(N__16145),
            .I(\uu2.w_addr_userZ0Z_7 ));
    CascadeMux I__3371 (
            .O(N__16140),
            .I(N__16136));
    InMux I__3370 (
            .O(N__16139),
            .I(N__16125));
    InMux I__3369 (
            .O(N__16136),
            .I(N__16125));
    InMux I__3368 (
            .O(N__16135),
            .I(N__16125));
    InMux I__3367 (
            .O(N__16134),
            .I(N__16125));
    LocalMux I__3366 (
            .O(N__16125),
            .I(\uu2.w_addr_userZ0Z_3 ));
    InMux I__3365 (
            .O(N__16122),
            .I(N__16117));
    CascadeMux I__3364 (
            .O(N__16121),
            .I(N__16110));
    CascadeMux I__3363 (
            .O(N__16120),
            .I(N__16107));
    LocalMux I__3362 (
            .O(N__16117),
            .I(N__16103));
    InMux I__3361 (
            .O(N__16116),
            .I(N__16100));
    CascadeMux I__3360 (
            .O(N__16115),
            .I(N__16095));
    InMux I__3359 (
            .O(N__16114),
            .I(N__16090));
    InMux I__3358 (
            .O(N__16113),
            .I(N__16090));
    InMux I__3357 (
            .O(N__16110),
            .I(N__16085));
    InMux I__3356 (
            .O(N__16107),
            .I(N__16085));
    InMux I__3355 (
            .O(N__16106),
            .I(N__16082));
    Span4Mux_h I__3354 (
            .O(N__16103),
            .I(N__16077));
    LocalMux I__3353 (
            .O(N__16100),
            .I(N__16077));
    InMux I__3352 (
            .O(N__16099),
            .I(N__16072));
    InMux I__3351 (
            .O(N__16098),
            .I(N__16072));
    InMux I__3350 (
            .O(N__16095),
            .I(N__16069));
    LocalMux I__3349 (
            .O(N__16090),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3348 (
            .O(N__16085),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3347 (
            .O(N__16082),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__3346 (
            .O(N__16077),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3345 (
            .O(N__16072),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__3344 (
            .O(N__16069),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    CascadeMux I__3343 (
            .O(N__16056),
            .I(N__16053));
    InMux I__3342 (
            .O(N__16053),
            .I(N__16050));
    LocalMux I__3341 (
            .O(N__16050),
            .I(N__16047));
    Span4Mux_h I__3340 (
            .O(N__16047),
            .I(N__16044));
    Odrv4 I__3339 (
            .O(N__16044),
            .I(\uu2.mem0.w_addr_3 ));
    InMux I__3338 (
            .O(N__16041),
            .I(N__16036));
    InMux I__3337 (
            .O(N__16040),
            .I(N__16033));
    CascadeMux I__3336 (
            .O(N__16039),
            .I(N__16030));
    LocalMux I__3335 (
            .O(N__16036),
            .I(N__16025));
    LocalMux I__3334 (
            .O(N__16033),
            .I(N__16025));
    InMux I__3333 (
            .O(N__16030),
            .I(N__16022));
    Odrv4 I__3332 (
            .O(N__16025),
            .I(\uu2.un426_ci_3 ));
    LocalMux I__3331 (
            .O(N__16022),
            .I(\uu2.un426_ci_3 ));
    CascadeMux I__3330 (
            .O(N__16017),
            .I(N__16013));
    InMux I__3329 (
            .O(N__16016),
            .I(N__16005));
    InMux I__3328 (
            .O(N__16013),
            .I(N__16005));
    InMux I__3327 (
            .O(N__16012),
            .I(N__16005));
    LocalMux I__3326 (
            .O(N__16005),
            .I(N__16002));
    Span4Mux_h I__3325 (
            .O(N__16002),
            .I(N__15998));
    InMux I__3324 (
            .O(N__16001),
            .I(N__15995));
    Odrv4 I__3323 (
            .O(N__15998),
            .I(\uu2.un404_ci ));
    LocalMux I__3322 (
            .O(N__15995),
            .I(\uu2.un404_ci ));
    CascadeMux I__3321 (
            .O(N__15990),
            .I(N__15987));
    InMux I__3320 (
            .O(N__15987),
            .I(N__15984));
    LocalMux I__3319 (
            .O(N__15984),
            .I(N__15981));
    Odrv12 I__3318 (
            .O(N__15981),
            .I(\uu2.vbuf_w_addr_user.un448_ci_0 ));
    InMux I__3317 (
            .O(N__15978),
            .I(N__15975));
    LocalMux I__3316 (
            .O(N__15975),
            .I(N__15970));
    InMux I__3315 (
            .O(N__15974),
            .I(N__15965));
    InMux I__3314 (
            .O(N__15973),
            .I(N__15965));
    Odrv12 I__3313 (
            .O(N__15970),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__3312 (
            .O(N__15965),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CEMux I__3311 (
            .O(N__15960),
            .I(N__15957));
    LocalMux I__3310 (
            .O(N__15957),
            .I(N__15954));
    Sp12to4 I__3309 (
            .O(N__15954),
            .I(N__15951));
    Odrv12 I__3308 (
            .O(N__15951),
            .I(\uu2.un28_w_addr_user_i_0 ));
    SRMux I__3307 (
            .O(N__15948),
            .I(N__15945));
    LocalMux I__3306 (
            .O(N__15945),
            .I(N__15942));
    Span4Mux_s0_v I__3305 (
            .O(N__15942),
            .I(N__15938));
    SRMux I__3304 (
            .O(N__15941),
            .I(N__15935));
    Span4Mux_h I__3303 (
            .O(N__15938),
            .I(N__15930));
    LocalMux I__3302 (
            .O(N__15935),
            .I(N__15930));
    Span4Mux_s0_v I__3301 (
            .O(N__15930),
            .I(N__15926));
    InMux I__3300 (
            .O(N__15929),
            .I(N__15923));
    Odrv4 I__3299 (
            .O(N__15926),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_4 ));
    LocalMux I__3298 (
            .O(N__15923),
            .I(\uu2.w_addr_user_RNI43E87Z0Z_4 ));
    InMux I__3297 (
            .O(N__15918),
            .I(N__15914));
    InMux I__3296 (
            .O(N__15917),
            .I(N__15911));
    LocalMux I__3295 (
            .O(N__15914),
            .I(N__15908));
    LocalMux I__3294 (
            .O(N__15911),
            .I(N__15905));
    Span4Mux_h I__3293 (
            .O(N__15908),
            .I(N__15902));
    Span4Mux_h I__3292 (
            .O(N__15905),
            .I(N__15899));
    Span4Mux_h I__3291 (
            .O(N__15902),
            .I(N__15896));
    Odrv4 I__3290 (
            .O(N__15899),
            .I(\uu2.N_44 ));
    Odrv4 I__3289 (
            .O(N__15896),
            .I(\uu2.N_44 ));
    InMux I__3288 (
            .O(N__15891),
            .I(N__15882));
    InMux I__3287 (
            .O(N__15890),
            .I(N__15882));
    InMux I__3286 (
            .O(N__15889),
            .I(N__15882));
    LocalMux I__3285 (
            .O(N__15882),
            .I(N__15873));
    InMux I__3284 (
            .O(N__15881),
            .I(N__15868));
    InMux I__3283 (
            .O(N__15880),
            .I(N__15868));
    InMux I__3282 (
            .O(N__15879),
            .I(N__15863));
    InMux I__3281 (
            .O(N__15878),
            .I(N__15856));
    InMux I__3280 (
            .O(N__15877),
            .I(N__15856));
    InMux I__3279 (
            .O(N__15876),
            .I(N__15856));
    Span4Mux_v I__3278 (
            .O(N__15873),
            .I(N__15853));
    LocalMux I__3277 (
            .O(N__15868),
            .I(N__15850));
    InMux I__3276 (
            .O(N__15867),
            .I(N__15845));
    InMux I__3275 (
            .O(N__15866),
            .I(N__15845));
    LocalMux I__3274 (
            .O(N__15863),
            .I(N__15842));
    LocalMux I__3273 (
            .O(N__15856),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    Odrv4 I__3272 (
            .O(N__15853),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    Odrv4 I__3271 (
            .O(N__15850),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    LocalMux I__3270 (
            .O(N__15845),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    Odrv4 I__3269 (
            .O(N__15842),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ));
    InMux I__3268 (
            .O(N__15831),
            .I(N__15828));
    LocalMux I__3267 (
            .O(N__15828),
            .I(N__15824));
    InMux I__3266 (
            .O(N__15827),
            .I(N__15821));
    Odrv4 I__3265 (
            .O(N__15824),
            .I(bu_rx_data_fast_6));
    LocalMux I__3264 (
            .O(N__15821),
            .I(bu_rx_data_fast_6));
    CascadeMux I__3263 (
            .O(N__15816),
            .I(N__15812));
    InMux I__3262 (
            .O(N__15815),
            .I(N__15809));
    InMux I__3261 (
            .O(N__15812),
            .I(N__15806));
    LocalMux I__3260 (
            .O(N__15809),
            .I(N__15801));
    LocalMux I__3259 (
            .O(N__15806),
            .I(N__15801));
    Odrv4 I__3258 (
            .O(N__15801),
            .I(bu_rx_data_fast_5));
    CascadeMux I__3257 (
            .O(N__15798),
            .I(\Lab_UT.dictrl.g1_0_4_cascade_ ));
    InMux I__3256 (
            .O(N__15795),
            .I(N__15792));
    LocalMux I__3255 (
            .O(N__15792),
            .I(\Lab_UT.dictrl.g1_0_xZ0Z1 ));
    InMux I__3254 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__3253 (
            .O(N__15786),
            .I(\Lab_UT.dictrl.g0_5Z0Z_4 ));
    InMux I__3252 (
            .O(N__15783),
            .I(N__15780));
    LocalMux I__3251 (
            .O(N__15780),
            .I(\Lab_UT.dictrl.g0_5_3 ));
    CascadeMux I__3250 (
            .O(N__15777),
            .I(\Lab_UT.dictrl.g1_0_cascade_ ));
    InMux I__3249 (
            .O(N__15774),
            .I(N__15770));
    InMux I__3248 (
            .O(N__15773),
            .I(N__15767));
    LocalMux I__3247 (
            .O(N__15770),
            .I(N__15764));
    LocalMux I__3246 (
            .O(N__15767),
            .I(N__15761));
    Span4Mux_v I__3245 (
            .O(N__15764),
            .I(N__15758));
    Span4Mux_v I__3244 (
            .O(N__15761),
            .I(N__15755));
    Odrv4 I__3243 (
            .O(N__15758),
            .I(\Lab_UT.dictrl.N_55_0 ));
    Odrv4 I__3242 (
            .O(N__15755),
            .I(\Lab_UT.dictrl.N_55_0 ));
    CascadeMux I__3241 (
            .O(N__15750),
            .I(\Lab_UT.dictrl.g0_3_4_cascade_ ));
    InMux I__3240 (
            .O(N__15747),
            .I(N__15731));
    InMux I__3239 (
            .O(N__15746),
            .I(N__15731));
    InMux I__3238 (
            .O(N__15745),
            .I(N__15728));
    InMux I__3237 (
            .O(N__15744),
            .I(N__15719));
    InMux I__3236 (
            .O(N__15743),
            .I(N__15719));
    InMux I__3235 (
            .O(N__15742),
            .I(N__15719));
    InMux I__3234 (
            .O(N__15741),
            .I(N__15719));
    InMux I__3233 (
            .O(N__15740),
            .I(N__15716));
    InMux I__3232 (
            .O(N__15739),
            .I(N__15711));
    InMux I__3231 (
            .O(N__15738),
            .I(N__15711));
    InMux I__3230 (
            .O(N__15737),
            .I(N__15706));
    InMux I__3229 (
            .O(N__15736),
            .I(N__15706));
    LocalMux I__3228 (
            .O(N__15731),
            .I(N__15699));
    LocalMux I__3227 (
            .O(N__15728),
            .I(N__15699));
    LocalMux I__3226 (
            .O(N__15719),
            .I(N__15699));
    LocalMux I__3225 (
            .O(N__15716),
            .I(N__15696));
    LocalMux I__3224 (
            .O(N__15711),
            .I(N__15691));
    LocalMux I__3223 (
            .O(N__15706),
            .I(N__15691));
    Span4Mux_v I__3222 (
            .O(N__15699),
            .I(N__15688));
    Odrv4 I__3221 (
            .O(N__15696),
            .I(bu_rx_data_5));
    Odrv4 I__3220 (
            .O(N__15691),
            .I(bu_rx_data_5));
    Odrv4 I__3219 (
            .O(N__15688),
            .I(bu_rx_data_5));
    InMux I__3218 (
            .O(N__15681),
            .I(N__15678));
    LocalMux I__3217 (
            .O(N__15678),
            .I(N__15675));
    Span4Mux_v I__3216 (
            .O(N__15675),
            .I(N__15672));
    Odrv4 I__3215 (
            .O(N__15672),
            .I(\Lab_UT.dictrl.N_72_mux_0 ));
    InMux I__3214 (
            .O(N__15669),
            .I(N__15662));
    InMux I__3213 (
            .O(N__15668),
            .I(N__15657));
    InMux I__3212 (
            .O(N__15667),
            .I(N__15657));
    InMux I__3211 (
            .O(N__15666),
            .I(N__15652));
    InMux I__3210 (
            .O(N__15665),
            .I(N__15652));
    LocalMux I__3209 (
            .O(N__15662),
            .I(bu_rx_data_6_rep1));
    LocalMux I__3208 (
            .O(N__15657),
            .I(bu_rx_data_6_rep1));
    LocalMux I__3207 (
            .O(N__15652),
            .I(bu_rx_data_6_rep1));
    CascadeMux I__3206 (
            .O(N__15645),
            .I(N__15638));
    InMux I__3205 (
            .O(N__15644),
            .I(N__15635));
    InMux I__3204 (
            .O(N__15643),
            .I(N__15630));
    InMux I__3203 (
            .O(N__15642),
            .I(N__15630));
    InMux I__3202 (
            .O(N__15641),
            .I(N__15625));
    InMux I__3201 (
            .O(N__15638),
            .I(N__15625));
    LocalMux I__3200 (
            .O(N__15635),
            .I(bu_rx_data_7_rep1));
    LocalMux I__3199 (
            .O(N__15630),
            .I(bu_rx_data_7_rep1));
    LocalMux I__3198 (
            .O(N__15625),
            .I(bu_rx_data_7_rep1));
    InMux I__3197 (
            .O(N__15618),
            .I(N__15615));
    LocalMux I__3196 (
            .O(N__15615),
            .I(\Lab_UT.dictrl.g0_3_3 ));
    InMux I__3195 (
            .O(N__15612),
            .I(N__15604));
    InMux I__3194 (
            .O(N__15611),
            .I(N__15604));
    CascadeMux I__3193 (
            .O(N__15610),
            .I(N__15597));
    InMux I__3192 (
            .O(N__15609),
            .I(N__15593));
    LocalMux I__3191 (
            .O(N__15604),
            .I(N__15590));
    CascadeMux I__3190 (
            .O(N__15603),
            .I(N__15584));
    InMux I__3189 (
            .O(N__15602),
            .I(N__15580));
    InMux I__3188 (
            .O(N__15601),
            .I(N__15577));
    InMux I__3187 (
            .O(N__15600),
            .I(N__15574));
    InMux I__3186 (
            .O(N__15597),
            .I(N__15571));
    InMux I__3185 (
            .O(N__15596),
            .I(N__15568));
    LocalMux I__3184 (
            .O(N__15593),
            .I(N__15565));
    Span4Mux_h I__3183 (
            .O(N__15590),
            .I(N__15562));
    InMux I__3182 (
            .O(N__15589),
            .I(N__15559));
    InMux I__3181 (
            .O(N__15588),
            .I(N__15556));
    InMux I__3180 (
            .O(N__15587),
            .I(N__15549));
    InMux I__3179 (
            .O(N__15584),
            .I(N__15549));
    InMux I__3178 (
            .O(N__15583),
            .I(N__15549));
    LocalMux I__3177 (
            .O(N__15580),
            .I(bu_rx_data_4));
    LocalMux I__3176 (
            .O(N__15577),
            .I(bu_rx_data_4));
    LocalMux I__3175 (
            .O(N__15574),
            .I(bu_rx_data_4));
    LocalMux I__3174 (
            .O(N__15571),
            .I(bu_rx_data_4));
    LocalMux I__3173 (
            .O(N__15568),
            .I(bu_rx_data_4));
    Odrv4 I__3172 (
            .O(N__15565),
            .I(bu_rx_data_4));
    Odrv4 I__3171 (
            .O(N__15562),
            .I(bu_rx_data_4));
    LocalMux I__3170 (
            .O(N__15559),
            .I(bu_rx_data_4));
    LocalMux I__3169 (
            .O(N__15556),
            .I(bu_rx_data_4));
    LocalMux I__3168 (
            .O(N__15549),
            .I(bu_rx_data_4));
    CascadeMux I__3167 (
            .O(N__15528),
            .I(N__15525));
    InMux I__3166 (
            .O(N__15525),
            .I(N__15522));
    LocalMux I__3165 (
            .O(N__15522),
            .I(N__15516));
    InMux I__3164 (
            .O(N__15521),
            .I(N__15513));
    InMux I__3163 (
            .O(N__15520),
            .I(N__15508));
    InMux I__3162 (
            .O(N__15519),
            .I(N__15508));
    Span4Mux_h I__3161 (
            .O(N__15516),
            .I(N__15505));
    LocalMux I__3160 (
            .O(N__15513),
            .I(\uu2.w_addr_userZ0Z_5 ));
    LocalMux I__3159 (
            .O(N__15508),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__3158 (
            .O(N__15505),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CascadeMux I__3157 (
            .O(N__15498),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ));
    CascadeMux I__3156 (
            .O(N__15495),
            .I(N__15491));
    InMux I__3155 (
            .O(N__15494),
            .I(N__15487));
    InMux I__3154 (
            .O(N__15491),
            .I(N__15481));
    InMux I__3153 (
            .O(N__15490),
            .I(N__15481));
    LocalMux I__3152 (
            .O(N__15487),
            .I(N__15478));
    CascadeMux I__3151 (
            .O(N__15486),
            .I(N__15475));
    LocalMux I__3150 (
            .O(N__15481),
            .I(N__15472));
    Span4Mux_v I__3149 (
            .O(N__15478),
            .I(N__15469));
    InMux I__3148 (
            .O(N__15475),
            .I(N__15466));
    Odrv12 I__3147 (
            .O(N__15472),
            .I(\Lab_UT.dictrl.N_18 ));
    Odrv4 I__3146 (
            .O(N__15469),
            .I(\Lab_UT.dictrl.N_18 ));
    LocalMux I__3145 (
            .O(N__15466),
            .I(\Lab_UT.dictrl.N_18 ));
    InMux I__3144 (
            .O(N__15459),
            .I(N__15451));
    InMux I__3143 (
            .O(N__15458),
            .I(N__15451));
    InMux I__3142 (
            .O(N__15457),
            .I(N__15446));
    InMux I__3141 (
            .O(N__15456),
            .I(N__15446));
    LocalMux I__3140 (
            .O(N__15451),
            .I(m7_a0));
    LocalMux I__3139 (
            .O(N__15446),
            .I(m7_a0));
    CascadeMux I__3138 (
            .O(N__15441),
            .I(N__15436));
    CascadeMux I__3137 (
            .O(N__15440),
            .I(N__15433));
    CascadeMux I__3136 (
            .O(N__15439),
            .I(N__15430));
    InMux I__3135 (
            .O(N__15436),
            .I(N__15427));
    InMux I__3134 (
            .O(N__15433),
            .I(N__15422));
    InMux I__3133 (
            .O(N__15430),
            .I(N__15422));
    LocalMux I__3132 (
            .O(N__15427),
            .I(N__15419));
    LocalMux I__3131 (
            .O(N__15422),
            .I(N__15416));
    Sp12to4 I__3130 (
            .O(N__15419),
            .I(N__15411));
    Sp12to4 I__3129 (
            .O(N__15416),
            .I(N__15411));
    Odrv12 I__3128 (
            .O(N__15411),
            .I(\Lab_UT.dictrl.state_fast_0 ));
    InMux I__3127 (
            .O(N__15408),
            .I(N__15405));
    LocalMux I__3126 (
            .O(N__15405),
            .I(N__15402));
    Span4Mux_h I__3125 (
            .O(N__15402),
            .I(N__15395));
    InMux I__3124 (
            .O(N__15401),
            .I(N__15388));
    InMux I__3123 (
            .O(N__15400),
            .I(N__15388));
    InMux I__3122 (
            .O(N__15399),
            .I(N__15388));
    InMux I__3121 (
            .O(N__15398),
            .I(N__15385));
    Odrv4 I__3120 (
            .O(N__15395),
            .I(buart__rx_shifter_fast_4));
    LocalMux I__3119 (
            .O(N__15388),
            .I(buart__rx_shifter_fast_4));
    LocalMux I__3118 (
            .O(N__15385),
            .I(buart__rx_shifter_fast_4));
    InMux I__3117 (
            .O(N__15378),
            .I(N__15371));
    InMux I__3116 (
            .O(N__15377),
            .I(N__15371));
    CascadeMux I__3115 (
            .O(N__15376),
            .I(N__15368));
    LocalMux I__3114 (
            .O(N__15371),
            .I(N__15364));
    InMux I__3113 (
            .O(N__15368),
            .I(N__15359));
    InMux I__3112 (
            .O(N__15367),
            .I(N__15359));
    Odrv4 I__3111 (
            .O(N__15364),
            .I(bu_rx_data_5_rep1));
    LocalMux I__3110 (
            .O(N__15359),
            .I(bu_rx_data_5_rep1));
    CascadeMux I__3109 (
            .O(N__15354),
            .I(\Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_ ));
    InMux I__3108 (
            .O(N__15351),
            .I(N__15348));
    LocalMux I__3107 (
            .O(N__15348),
            .I(N__15345));
    Odrv4 I__3106 (
            .O(N__15345),
            .I(\Lab_UT.dictrl.g0_6_3 ));
    CascadeMux I__3105 (
            .O(N__15342),
            .I(N__15338));
    InMux I__3104 (
            .O(N__15341),
            .I(N__15335));
    InMux I__3103 (
            .O(N__15338),
            .I(N__15332));
    LocalMux I__3102 (
            .O(N__15335),
            .I(\Lab_UT.dictrl.gZ0Z2 ));
    LocalMux I__3101 (
            .O(N__15332),
            .I(\Lab_UT.dictrl.gZ0Z2 ));
    CascadeMux I__3100 (
            .O(N__15327),
            .I(\Lab_UT.dictrl.g0_6_3_cascade_ ));
    InMux I__3099 (
            .O(N__15324),
            .I(N__15321));
    LocalMux I__3098 (
            .O(N__15321),
            .I(N__15317));
    InMux I__3097 (
            .O(N__15320),
            .I(N__15314));
    Odrv4 I__3096 (
            .O(N__15317),
            .I(\Lab_UT.dictrl.g1_1 ));
    LocalMux I__3095 (
            .O(N__15314),
            .I(\Lab_UT.dictrl.g1_1 ));
    InMux I__3094 (
            .O(N__15309),
            .I(N__15303));
    InMux I__3093 (
            .O(N__15308),
            .I(N__15303));
    LocalMux I__3092 (
            .O(N__15303),
            .I(N__15300));
    Span4Mux_v I__3091 (
            .O(N__15300),
            .I(N__15297));
    Odrv4 I__3090 (
            .O(N__15297),
            .I(\Lab_UT.dictrl.N_57_0 ));
    CascadeMux I__3089 (
            .O(N__15294),
            .I(N_5_cascade_));
    CascadeMux I__3088 (
            .O(N__15291),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ));
    InMux I__3087 (
            .O(N__15288),
            .I(N__15285));
    LocalMux I__3086 (
            .O(N__15285),
            .I(\Lab_UT.dictrl.N_59_1_0 ));
    InMux I__3085 (
            .O(N__15282),
            .I(N__15276));
    InMux I__3084 (
            .O(N__15281),
            .I(N__15276));
    LocalMux I__3083 (
            .O(N__15276),
            .I(\Lab_UT.dictrl.i8_mux_0 ));
    InMux I__3082 (
            .O(N__15273),
            .I(N__15270));
    LocalMux I__3081 (
            .O(N__15270),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13 ));
    CascadeMux I__3080 (
            .O(N__15267),
            .I(\Lab_UT.dictrl.m22_xZ0Z1_cascade_ ));
    InMux I__3079 (
            .O(N__15264),
            .I(N__15259));
    InMux I__3078 (
            .O(N__15263),
            .I(N__15253));
    InMux I__3077 (
            .O(N__15262),
            .I(N__15253));
    LocalMux I__3076 (
            .O(N__15259),
            .I(N__15250));
    InMux I__3075 (
            .O(N__15258),
            .I(N__15247));
    LocalMux I__3074 (
            .O(N__15253),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    Odrv4 I__3073 (
            .O(N__15250),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    LocalMux I__3072 (
            .O(N__15247),
            .I(\Lab_UT.dictrl.m22Z0Z_4 ));
    CascadeMux I__3071 (
            .O(N__15240),
            .I(\Lab_UT.dictrl.N_72_mux_cascade_ ));
    InMux I__3070 (
            .O(N__15237),
            .I(N__15234));
    LocalMux I__3069 (
            .O(N__15234),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ));
    CascadeMux I__3068 (
            .O(N__15231),
            .I(\Lab_UT.dictrl.m34_0_cascade_ ));
    CascadeMux I__3067 (
            .O(N__15228),
            .I(\Lab_UT.dictrl.next_state_1_3_cascade_ ));
    CascadeMux I__3066 (
            .O(N__15225),
            .I(N__15221));
    CascadeMux I__3065 (
            .O(N__15224),
            .I(N__15217));
    InMux I__3064 (
            .O(N__15221),
            .I(N__15210));
    InMux I__3063 (
            .O(N__15220),
            .I(N__15210));
    InMux I__3062 (
            .O(N__15217),
            .I(N__15210));
    LocalMux I__3061 (
            .O(N__15210),
            .I(N__15207));
    Span4Mux_v I__3060 (
            .O(N__15207),
            .I(N__15204));
    Odrv4 I__3059 (
            .O(N__15204),
            .I(\Lab_UT.dictrl.next_stateZ0Z_3 ));
    CascadeMux I__3058 (
            .O(N__15201),
            .I(\Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ));
    InMux I__3057 (
            .O(N__15198),
            .I(N__15186));
    InMux I__3056 (
            .O(N__15197),
            .I(N__15186));
    InMux I__3055 (
            .O(N__15196),
            .I(N__15186));
    InMux I__3054 (
            .O(N__15195),
            .I(N__15186));
    LocalMux I__3053 (
            .O(N__15186),
            .I(N__15183));
    Odrv4 I__3052 (
            .O(N__15183),
            .I(\Lab_UT.dictrl.N_26_0 ));
    InMux I__3051 (
            .O(N__15180),
            .I(N__15177));
    LocalMux I__3050 (
            .O(N__15177),
            .I(\Lab_UT.dictrl.m34_0 ));
    CascadeMux I__3049 (
            .O(N__15174),
            .I(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_ ));
    InMux I__3048 (
            .O(N__15171),
            .I(N__15168));
    LocalMux I__3047 (
            .O(N__15168),
            .I(\Lab_UT.dictrl.N_60_0_0 ));
    InMux I__3046 (
            .O(N__15165),
            .I(N__15159));
    InMux I__3045 (
            .O(N__15164),
            .I(N__15159));
    LocalMux I__3044 (
            .O(N__15159),
            .I(N__15156));
    Odrv4 I__3043 (
            .O(N__15156),
            .I(\Lab_UT.dictrl.m19_1 ));
    InMux I__3042 (
            .O(N__15153),
            .I(N__15149));
    InMux I__3041 (
            .O(N__15152),
            .I(N__15146));
    LocalMux I__3040 (
            .O(N__15149),
            .I(N__15141));
    LocalMux I__3039 (
            .O(N__15146),
            .I(N__15141));
    Odrv4 I__3038 (
            .O(N__15141),
            .I(\Lab_UT.dictrl.N_22 ));
    CascadeMux I__3037 (
            .O(N__15138),
            .I(N__15135));
    InMux I__3036 (
            .O(N__15135),
            .I(N__15132));
    LocalMux I__3035 (
            .O(N__15132),
            .I(N__15129));
    Odrv4 I__3034 (
            .O(N__15129),
            .I(\Lab_UT.dictrl.next_state_0_1 ));
    CascadeMux I__3033 (
            .O(N__15126),
            .I(N__15123));
    InMux I__3032 (
            .O(N__15123),
            .I(N__15120));
    LocalMux I__3031 (
            .O(N__15120),
            .I(N__15117));
    Odrv4 I__3030 (
            .O(N__15117),
            .I(\Lab_UT.dictrl.g2_0_0 ));
    InMux I__3029 (
            .O(N__15114),
            .I(N__15104));
    InMux I__3028 (
            .O(N__15113),
            .I(N__15104));
    InMux I__3027 (
            .O(N__15112),
            .I(N__15104));
    CascadeMux I__3026 (
            .O(N__15111),
            .I(N__15101));
    LocalMux I__3025 (
            .O(N__15104),
            .I(N__15098));
    InMux I__3024 (
            .O(N__15101),
            .I(N__15095));
    Odrv4 I__3023 (
            .O(N__15098),
            .I(\Lab_UT.dictrl.state_i_4_2 ));
    LocalMux I__3022 (
            .O(N__15095),
            .I(\Lab_UT.dictrl.state_i_4_2 ));
    CascadeMux I__3021 (
            .O(N__15090),
            .I(\Lab_UT.dictrl.N_20_0_0_cascade_ ));
    InMux I__3020 (
            .O(N__15087),
            .I(N__15084));
    LocalMux I__3019 (
            .O(N__15084),
            .I(N__15081));
    Span4Mux_v I__3018 (
            .O(N__15081),
            .I(N__15078));
    Odrv4 I__3017 (
            .O(N__15078),
            .I(\Lab_UT.dictrl.N_22_0_0 ));
    InMux I__3016 (
            .O(N__15075),
            .I(N__15064));
    InMux I__3015 (
            .O(N__15074),
            .I(N__15064));
    InMux I__3014 (
            .O(N__15073),
            .I(N__15060));
    InMux I__3013 (
            .O(N__15072),
            .I(N__15051));
    InMux I__3012 (
            .O(N__15071),
            .I(N__15051));
    InMux I__3011 (
            .O(N__15070),
            .I(N__15051));
    InMux I__3010 (
            .O(N__15069),
            .I(N__15051));
    LocalMux I__3009 (
            .O(N__15064),
            .I(N__15048));
    InMux I__3008 (
            .O(N__15063),
            .I(N__15045));
    LocalMux I__3007 (
            .O(N__15060),
            .I(\Lab_UT.next_state_0 ));
    LocalMux I__3006 (
            .O(N__15051),
            .I(\Lab_UT.next_state_0 ));
    Odrv4 I__3005 (
            .O(N__15048),
            .I(\Lab_UT.next_state_0 ));
    LocalMux I__3004 (
            .O(N__15045),
            .I(\Lab_UT.next_state_0 ));
    CascadeMux I__3003 (
            .O(N__15036),
            .I(\Lab_UT.next_state_1_0_0_1_cascade_ ));
    InMux I__3002 (
            .O(N__15033),
            .I(N__15024));
    InMux I__3001 (
            .O(N__15032),
            .I(N__15015));
    InMux I__3000 (
            .O(N__15031),
            .I(N__15015));
    InMux I__2999 (
            .O(N__15030),
            .I(N__15015));
    InMux I__2998 (
            .O(N__15029),
            .I(N__15015));
    InMux I__2997 (
            .O(N__15028),
            .I(N__15010));
    InMux I__2996 (
            .O(N__15027),
            .I(N__15010));
    LocalMux I__2995 (
            .O(N__15024),
            .I(N__15007));
    LocalMux I__2994 (
            .O(N__15015),
            .I(\Lab_UT.next_state_2 ));
    LocalMux I__2993 (
            .O(N__15010),
            .I(\Lab_UT.next_state_2 ));
    Odrv4 I__2992 (
            .O(N__15007),
            .I(\Lab_UT.next_state_2 ));
    InMux I__2991 (
            .O(N__15000),
            .I(N__14987));
    InMux I__2990 (
            .O(N__14999),
            .I(N__14987));
    InMux I__2989 (
            .O(N__14998),
            .I(N__14987));
    InMux I__2988 (
            .O(N__14997),
            .I(N__14987));
    InMux I__2987 (
            .O(N__14996),
            .I(N__14984));
    LocalMux I__2986 (
            .O(N__14987),
            .I(N__14981));
    LocalMux I__2985 (
            .O(N__14984),
            .I(N__14975));
    Span4Mux_v I__2984 (
            .O(N__14981),
            .I(N__14971));
    InMux I__2983 (
            .O(N__14980),
            .I(N__14968));
    InMux I__2982 (
            .O(N__14979),
            .I(N__14963));
    InMux I__2981 (
            .O(N__14978),
            .I(N__14963));
    Sp12to4 I__2980 (
            .O(N__14975),
            .I(N__14958));
    InMux I__2979 (
            .O(N__14974),
            .I(N__14955));
    Sp12to4 I__2978 (
            .O(N__14971),
            .I(N__14948));
    LocalMux I__2977 (
            .O(N__14968),
            .I(N__14948));
    LocalMux I__2976 (
            .O(N__14963),
            .I(N__14948));
    InMux I__2975 (
            .O(N__14962),
            .I(N__14945));
    InMux I__2974 (
            .O(N__14961),
            .I(N__14942));
    Span12Mux_s4_v I__2973 (
            .O(N__14958),
            .I(N__14937));
    LocalMux I__2972 (
            .O(N__14955),
            .I(N__14937));
    Span12Mux_s11_h I__2971 (
            .O(N__14948),
            .I(N__14934));
    LocalMux I__2970 (
            .O(N__14945),
            .I(bu_rx_data_rdy));
    LocalMux I__2969 (
            .O(N__14942),
            .I(bu_rx_data_rdy));
    Odrv12 I__2968 (
            .O(N__14937),
            .I(bu_rx_data_rdy));
    Odrv12 I__2967 (
            .O(N__14934),
            .I(bu_rx_data_rdy));
    InMux I__2966 (
            .O(N__14925),
            .I(N__14922));
    LocalMux I__2965 (
            .O(N__14922),
            .I(\Lab_UT.didp.g0_0_2Z0Z_1 ));
    CascadeMux I__2964 (
            .O(N__14919),
            .I(N__14916));
    InMux I__2963 (
            .O(N__14916),
            .I(N__14911));
    CascadeMux I__2962 (
            .O(N__14915),
            .I(N__14907));
    IoInMux I__2961 (
            .O(N__14914),
            .I(N__14904));
    LocalMux I__2960 (
            .O(N__14911),
            .I(N__14901));
    InMux I__2959 (
            .O(N__14910),
            .I(N__14898));
    InMux I__2958 (
            .O(N__14907),
            .I(N__14895));
    LocalMux I__2957 (
            .O(N__14904),
            .I(N__14892));
    Sp12to4 I__2956 (
            .O(N__14901),
            .I(N__14885));
    LocalMux I__2955 (
            .O(N__14898),
            .I(N__14885));
    LocalMux I__2954 (
            .O(N__14895),
            .I(N__14885));
    Span4Mux_s0_h I__2953 (
            .O(N__14892),
            .I(N__14882));
    Odrv12 I__2952 (
            .O(N__14885),
            .I(rst));
    Odrv4 I__2951 (
            .O(N__14882),
            .I(rst));
    InMux I__2950 (
            .O(N__14877),
            .I(N__14874));
    LocalMux I__2949 (
            .O(N__14874),
            .I(\Lab_UT.didp.g0_0Z0Z_2 ));
    InMux I__2948 (
            .O(N__14871),
            .I(N__14865));
    InMux I__2947 (
            .O(N__14870),
            .I(N__14865));
    LocalMux I__2946 (
            .O(N__14865),
            .I(N__14862));
    Span4Mux_h I__2945 (
            .O(N__14862),
            .I(N__14859));
    Odrv4 I__2944 (
            .O(N__14859),
            .I(\Lab_UT.dictrl.next_state6 ));
    CascadeMux I__2943 (
            .O(N__14856),
            .I(\Lab_UT.dictrl.N_20_cascade_ ));
    CascadeMux I__2942 (
            .O(N__14853),
            .I(\Lab_UT.dictrl.un15_loadalarm_0_cascade_ ));
    InMux I__2941 (
            .O(N__14850),
            .I(N__14847));
    LocalMux I__2940 (
            .O(N__14847),
            .I(\Lab_UT.dictrl.loadalarm_0_0 ));
    InMux I__2939 (
            .O(N__14844),
            .I(N__14840));
    InMux I__2938 (
            .O(N__14843),
            .I(N__14837));
    LocalMux I__2937 (
            .O(N__14840),
            .I(N__14834));
    LocalMux I__2936 (
            .O(N__14837),
            .I(N__14831));
    Odrv4 I__2935 (
            .O(N__14834),
            .I(\Lab_UT.LdAStens ));
    Odrv4 I__2934 (
            .O(N__14831),
            .I(\Lab_UT.LdAStens ));
    CascadeMux I__2933 (
            .O(N__14826),
            .I(N__14823));
    InMux I__2932 (
            .O(N__14823),
            .I(N__14819));
    InMux I__2931 (
            .O(N__14822),
            .I(N__14816));
    LocalMux I__2930 (
            .O(N__14819),
            .I(\Lab_UT.dictrl.dicLdAMones_1 ));
    LocalMux I__2929 (
            .O(N__14816),
            .I(\Lab_UT.dictrl.dicLdAMones_1 ));
    InMux I__2928 (
            .O(N__14811),
            .I(N__14808));
    LocalMux I__2927 (
            .O(N__14808),
            .I(N__14805));
    Span4Mux_h I__2926 (
            .O(N__14805),
            .I(N__14802));
    Odrv4 I__2925 (
            .O(N__14802),
            .I(\Lab_UT.LdAMones ));
    CascadeMux I__2924 (
            .O(N__14799),
            .I(\Lab_UT.LdAMones_cascade_ ));
    InMux I__2923 (
            .O(N__14796),
            .I(N__14793));
    LocalMux I__2922 (
            .O(N__14793),
            .I(\Lab_UT.dictrl.g0_1_mb_rn_0 ));
    CascadeMux I__2921 (
            .O(N__14790),
            .I(\Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ));
    InMux I__2920 (
            .O(N__14787),
            .I(N__14784));
    LocalMux I__2919 (
            .O(N__14784),
            .I(N__14780));
    InMux I__2918 (
            .O(N__14783),
            .I(N__14777));
    Span4Mux_v I__2917 (
            .O(N__14780),
            .I(N__14774));
    LocalMux I__2916 (
            .O(N__14777),
            .I(N__14771));
    Span4Mux_v I__2915 (
            .O(N__14774),
            .I(N__14768));
    Span4Mux_h I__2914 (
            .O(N__14771),
            .I(N__14765));
    Odrv4 I__2913 (
            .O(N__14768),
            .I(\Lab_UT.dictrl.N_57_1 ));
    Odrv4 I__2912 (
            .O(N__14765),
            .I(\Lab_UT.dictrl.N_57_1 ));
    CascadeMux I__2911 (
            .O(N__14760),
            .I(N__14757));
    InMux I__2910 (
            .O(N__14757),
            .I(N__14754));
    LocalMux I__2909 (
            .O(N__14754),
            .I(N__14750));
    CascadeMux I__2908 (
            .O(N__14753),
            .I(N__14747));
    Span4Mux_s2_v I__2907 (
            .O(N__14750),
            .I(N__14744));
    InMux I__2906 (
            .O(N__14747),
            .I(N__14741));
    Span4Mux_v I__2905 (
            .O(N__14744),
            .I(N__14738));
    LocalMux I__2904 (
            .O(N__14741),
            .I(N__14735));
    Span4Mux_v I__2903 (
            .O(N__14738),
            .I(N__14732));
    Span4Mux_h I__2902 (
            .O(N__14735),
            .I(N__14729));
    Odrv4 I__2901 (
            .O(N__14732),
            .I(\Lab_UT.dictrl.N_55_1 ));
    Odrv4 I__2900 (
            .O(N__14729),
            .I(\Lab_UT.dictrl.N_55_1 ));
    InMux I__2899 (
            .O(N__14724),
            .I(N__14721));
    LocalMux I__2898 (
            .O(N__14721),
            .I(N__14717));
    CascadeMux I__2897 (
            .O(N__14720),
            .I(N__14713));
    Span4Mux_v I__2896 (
            .O(N__14717),
            .I(N__14710));
    InMux I__2895 (
            .O(N__14716),
            .I(N__14705));
    InMux I__2894 (
            .O(N__14713),
            .I(N__14705));
    Span4Mux_v I__2893 (
            .O(N__14710),
            .I(N__14702));
    LocalMux I__2892 (
            .O(N__14705),
            .I(N__14699));
    Odrv4 I__2891 (
            .O(N__14702),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    Odrv12 I__2890 (
            .O(N__14699),
            .I(\Lab_UT.dictrl.next_state_0_2 ));
    CascadeMux I__2889 (
            .O(N__14694),
            .I(\Lab_UT.dictrl.next_state_1_2_cascade_ ));
    InMux I__2888 (
            .O(N__14691),
            .I(N__14685));
    InMux I__2887 (
            .O(N__14690),
            .I(N__14685));
    LocalMux I__2886 (
            .O(N__14685),
            .I(\Lab_UT.dictrl.g0_1_mb_sn ));
    InMux I__2885 (
            .O(N__14682),
            .I(N__14675));
    InMux I__2884 (
            .O(N__14681),
            .I(N__14675));
    InMux I__2883 (
            .O(N__14680),
            .I(N__14672));
    LocalMux I__2882 (
            .O(N__14675),
            .I(N__14669));
    LocalMux I__2881 (
            .O(N__14672),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv12 I__2880 (
            .O(N__14669),
            .I(\Lab_UT.di_AMtens_2 ));
    InMux I__2879 (
            .O(N__14664),
            .I(N__14661));
    LocalMux I__2878 (
            .O(N__14661),
            .I(N__14652));
    InMux I__2877 (
            .O(N__14660),
            .I(N__14639));
    InMux I__2876 (
            .O(N__14659),
            .I(N__14639));
    InMux I__2875 (
            .O(N__14658),
            .I(N__14639));
    InMux I__2874 (
            .O(N__14657),
            .I(N__14639));
    InMux I__2873 (
            .O(N__14656),
            .I(N__14639));
    InMux I__2872 (
            .O(N__14655),
            .I(N__14639));
    Span4Mux_s2_v I__2871 (
            .O(N__14652),
            .I(N__14636));
    LocalMux I__2870 (
            .O(N__14639),
            .I(N__14633));
    Odrv4 I__2869 (
            .O(N__14636),
            .I(\Lab_UT.min1_2 ));
    Odrv12 I__2868 (
            .O(N__14633),
            .I(\Lab_UT.min1_2 ));
    CEMux I__2867 (
            .O(N__14628),
            .I(N__14625));
    LocalMux I__2866 (
            .O(N__14625),
            .I(N__14622));
    Span4Mux_v I__2865 (
            .O(N__14622),
            .I(N__14618));
    CEMux I__2864 (
            .O(N__14621),
            .I(N__14615));
    Span4Mux_h I__2863 (
            .O(N__14618),
            .I(N__14612));
    LocalMux I__2862 (
            .O(N__14615),
            .I(N__14609));
    Odrv4 I__2861 (
            .O(N__14612),
            .I(\Lab_UT.didp.regrce3.LdAMones_0 ));
    Odrv12 I__2860 (
            .O(N__14609),
            .I(\Lab_UT.didp.regrce3.LdAMones_0 ));
    InMux I__2859 (
            .O(N__14604),
            .I(N__14595));
    InMux I__2858 (
            .O(N__14603),
            .I(N__14595));
    InMux I__2857 (
            .O(N__14602),
            .I(N__14595));
    LocalMux I__2856 (
            .O(N__14595),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__2855 (
            .O(N__14592),
            .I(N__14588));
    InMux I__2854 (
            .O(N__14591),
            .I(N__14585));
    LocalMux I__2853 (
            .O(N__14588),
            .I(N__14580));
    LocalMux I__2852 (
            .O(N__14585),
            .I(N__14580));
    Span4Mux_v I__2851 (
            .O(N__14580),
            .I(N__14576));
    InMux I__2850 (
            .O(N__14579),
            .I(N__14573));
    Span4Mux_v I__2849 (
            .O(N__14576),
            .I(N__14570));
    LocalMux I__2848 (
            .O(N__14573),
            .I(N__14567));
    Odrv4 I__2847 (
            .O(N__14570),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv12 I__2846 (
            .O(N__14567),
            .I(\Lab_UT.di_AStens_1 ));
    CascadeMux I__2845 (
            .O(N__14562),
            .I(\Lab_UT.dispString.N_118_cascade_ ));
    InMux I__2844 (
            .O(N__14559),
            .I(N__14556));
    LocalMux I__2843 (
            .O(N__14556),
            .I(N__14553));
    Span4Mux_h I__2842 (
            .O(N__14553),
            .I(N__14550));
    Odrv4 I__2841 (
            .O(N__14550),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_1 ));
    InMux I__2840 (
            .O(N__14547),
            .I(N__14543));
    CascadeMux I__2839 (
            .O(N__14546),
            .I(N__14540));
    LocalMux I__2838 (
            .O(N__14543),
            .I(N__14537));
    InMux I__2837 (
            .O(N__14540),
            .I(N__14534));
    Span4Mux_v I__2836 (
            .O(N__14537),
            .I(N__14528));
    LocalMux I__2835 (
            .O(N__14534),
            .I(N__14528));
    InMux I__2834 (
            .O(N__14533),
            .I(N__14525));
    Odrv4 I__2833 (
            .O(N__14528),
            .I(\Lab_UT.dispString.N_145 ));
    LocalMux I__2832 (
            .O(N__14525),
            .I(\Lab_UT.dispString.N_145 ));
    InMux I__2831 (
            .O(N__14520),
            .I(N__14516));
    InMux I__2830 (
            .O(N__14519),
            .I(N__14512));
    LocalMux I__2829 (
            .O(N__14516),
            .I(N__14509));
    InMux I__2828 (
            .O(N__14515),
            .I(N__14506));
    LocalMux I__2827 (
            .O(N__14512),
            .I(N__14501));
    Span4Mux_v I__2826 (
            .O(N__14509),
            .I(N__14501));
    LocalMux I__2825 (
            .O(N__14506),
            .I(N__14498));
    Odrv4 I__2824 (
            .O(N__14501),
            .I(\Lab_UT.di_AMtens_1 ));
    Odrv12 I__2823 (
            .O(N__14498),
            .I(\Lab_UT.di_AMtens_1 ));
    CascadeMux I__2822 (
            .O(N__14493),
            .I(N__14487));
    CascadeMux I__2821 (
            .O(N__14492),
            .I(N__14483));
    CascadeMux I__2820 (
            .O(N__14491),
            .I(N__14479));
    InMux I__2819 (
            .O(N__14490),
            .I(N__14475));
    InMux I__2818 (
            .O(N__14487),
            .I(N__14462));
    InMux I__2817 (
            .O(N__14486),
            .I(N__14462));
    InMux I__2816 (
            .O(N__14483),
            .I(N__14462));
    InMux I__2815 (
            .O(N__14482),
            .I(N__14462));
    InMux I__2814 (
            .O(N__14479),
            .I(N__14462));
    InMux I__2813 (
            .O(N__14478),
            .I(N__14462));
    LocalMux I__2812 (
            .O(N__14475),
            .I(N__14457));
    LocalMux I__2811 (
            .O(N__14462),
            .I(N__14457));
    Odrv4 I__2810 (
            .O(N__14457),
            .I(\Lab_UT.min1_1 ));
    InMux I__2809 (
            .O(N__14454),
            .I(N__14443));
    InMux I__2808 (
            .O(N__14453),
            .I(N__14443));
    InMux I__2807 (
            .O(N__14452),
            .I(N__14443));
    InMux I__2806 (
            .O(N__14451),
            .I(N__14440));
    CascadeMux I__2805 (
            .O(N__14450),
            .I(N__14436));
    LocalMux I__2804 (
            .O(N__14443),
            .I(N__14431));
    LocalMux I__2803 (
            .O(N__14440),
            .I(N__14431));
    InMux I__2802 (
            .O(N__14439),
            .I(N__14426));
    InMux I__2801 (
            .O(N__14436),
            .I(N__14426));
    Odrv4 I__2800 (
            .O(N__14431),
            .I(\Lab_UT.di_Stens_2 ));
    LocalMux I__2799 (
            .O(N__14426),
            .I(\Lab_UT.di_Stens_2 ));
    InMux I__2798 (
            .O(N__14421),
            .I(N__14417));
    InMux I__2797 (
            .O(N__14420),
            .I(N__14414));
    LocalMux I__2796 (
            .O(N__14417),
            .I(N__14411));
    LocalMux I__2795 (
            .O(N__14414),
            .I(N__14405));
    Span4Mux_h I__2794 (
            .O(N__14411),
            .I(N__14405));
    InMux I__2793 (
            .O(N__14410),
            .I(N__14402));
    Span4Mux_v I__2792 (
            .O(N__14405),
            .I(N__14399));
    LocalMux I__2791 (
            .O(N__14402),
            .I(N__14396));
    Odrv4 I__2790 (
            .O(N__14399),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__2789 (
            .O(N__14396),
            .I(\Lab_UT.di_AStens_2 ));
    InMux I__2788 (
            .O(N__14391),
            .I(N__14373));
    InMux I__2787 (
            .O(N__14390),
            .I(N__14373));
    InMux I__2786 (
            .O(N__14389),
            .I(N__14373));
    InMux I__2785 (
            .O(N__14388),
            .I(N__14373));
    InMux I__2784 (
            .O(N__14387),
            .I(N__14373));
    InMux I__2783 (
            .O(N__14386),
            .I(N__14373));
    LocalMux I__2782 (
            .O(N__14373),
            .I(N__14369));
    InMux I__2781 (
            .O(N__14372),
            .I(N__14366));
    Odrv4 I__2780 (
            .O(N__14369),
            .I(\Lab_UT.sec1_2 ));
    LocalMux I__2779 (
            .O(N__14366),
            .I(\Lab_UT.sec1_2 ));
    InMux I__2778 (
            .O(N__14361),
            .I(N__14357));
    InMux I__2777 (
            .O(N__14360),
            .I(N__14352));
    LocalMux I__2776 (
            .O(N__14357),
            .I(N__14348));
    InMux I__2775 (
            .O(N__14356),
            .I(N__14343));
    InMux I__2774 (
            .O(N__14355),
            .I(N__14340));
    LocalMux I__2773 (
            .O(N__14352),
            .I(N__14337));
    InMux I__2772 (
            .O(N__14351),
            .I(N__14333));
    Span4Mux_h I__2771 (
            .O(N__14348),
            .I(N__14330));
    InMux I__2770 (
            .O(N__14347),
            .I(N__14327));
    InMux I__2769 (
            .O(N__14346),
            .I(N__14324));
    LocalMux I__2768 (
            .O(N__14343),
            .I(N__14317));
    LocalMux I__2767 (
            .O(N__14340),
            .I(N__14317));
    Span4Mux_s2_v I__2766 (
            .O(N__14337),
            .I(N__14317));
    InMux I__2765 (
            .O(N__14336),
            .I(N__14314));
    LocalMux I__2764 (
            .O(N__14333),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__2763 (
            .O(N__14330),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__2762 (
            .O(N__14327),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__2761 (
            .O(N__14324),
            .I(\Lab_UT.di_Sones_0 ));
    Odrv4 I__2760 (
            .O(N__14317),
            .I(\Lab_UT.di_Sones_0 ));
    LocalMux I__2759 (
            .O(N__14314),
            .I(\Lab_UT.di_Sones_0 ));
    InMux I__2758 (
            .O(N__14301),
            .I(N__14298));
    LocalMux I__2757 (
            .O(N__14298),
            .I(N__14295));
    Span4Mux_h I__2756 (
            .O(N__14295),
            .I(N__14289));
    CascadeMux I__2755 (
            .O(N__14294),
            .I(N__14286));
    InMux I__2754 (
            .O(N__14293),
            .I(N__14283));
    InMux I__2753 (
            .O(N__14292),
            .I(N__14280));
    Span4Mux_h I__2752 (
            .O(N__14289),
            .I(N__14277));
    InMux I__2751 (
            .O(N__14286),
            .I(N__14274));
    LocalMux I__2750 (
            .O(N__14283),
            .I(N__14271));
    LocalMux I__2749 (
            .O(N__14280),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__2748 (
            .O(N__14277),
            .I(\Lab_UT.LdSones ));
    LocalMux I__2747 (
            .O(N__14274),
            .I(\Lab_UT.LdSones ));
    Odrv12 I__2746 (
            .O(N__14271),
            .I(\Lab_UT.LdSones ));
    CascadeMux I__2745 (
            .O(N__14262),
            .I(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ));
    CascadeMux I__2744 (
            .O(N__14259),
            .I(N__14255));
    CascadeMux I__2743 (
            .O(N__14258),
            .I(N__14252));
    InMux I__2742 (
            .O(N__14255),
            .I(N__14246));
    InMux I__2741 (
            .O(N__14252),
            .I(N__14246));
    InMux I__2740 (
            .O(N__14251),
            .I(N__14243));
    LocalMux I__2739 (
            .O(N__14246),
            .I(N__14239));
    LocalMux I__2738 (
            .O(N__14243),
            .I(N__14236));
    InMux I__2737 (
            .O(N__14242),
            .I(N__14233));
    Span4Mux_v I__2736 (
            .O(N__14239),
            .I(N__14230));
    Span4Mux_v I__2735 (
            .O(N__14236),
            .I(N__14227));
    LocalMux I__2734 (
            .O(N__14233),
            .I(N__14224));
    Odrv4 I__2733 (
            .O(N__14230),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    Odrv4 I__2732 (
            .O(N__14227),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    Odrv12 I__2731 (
            .O(N__14224),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    CascadeMux I__2730 (
            .O(N__14217),
            .I(\Lab_UT.didp.countrce1.q_5_2_cascade_ ));
    InMux I__2729 (
            .O(N__14214),
            .I(N__14211));
    LocalMux I__2728 (
            .O(N__14211),
            .I(N__14205));
    InMux I__2727 (
            .O(N__14210),
            .I(N__14202));
    InMux I__2726 (
            .O(N__14209),
            .I(N__14199));
    InMux I__2725 (
            .O(N__14208),
            .I(N__14196));
    Odrv4 I__2724 (
            .O(N__14205),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    LocalMux I__2723 (
            .O(N__14202),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    LocalMux I__2722 (
            .O(N__14199),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    LocalMux I__2721 (
            .O(N__14196),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    InMux I__2720 (
            .O(N__14187),
            .I(N__14178));
    InMux I__2719 (
            .O(N__14186),
            .I(N__14178));
    InMux I__2718 (
            .O(N__14185),
            .I(N__14178));
    LocalMux I__2717 (
            .O(N__14178),
            .I(N__14175));
    Odrv4 I__2716 (
            .O(N__14175),
            .I(\Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ));
    InMux I__2715 (
            .O(N__14172),
            .I(N__14169));
    LocalMux I__2714 (
            .O(N__14169),
            .I(N__14166));
    Span4Mux_h I__2713 (
            .O(N__14166),
            .I(N__14163));
    Odrv4 I__2712 (
            .O(N__14163),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ));
    CascadeMux I__2711 (
            .O(N__14160),
            .I(N__14155));
    CascadeMux I__2710 (
            .O(N__14159),
            .I(N__14152));
    InMux I__2709 (
            .O(N__14158),
            .I(N__14140));
    InMux I__2708 (
            .O(N__14155),
            .I(N__14140));
    InMux I__2707 (
            .O(N__14152),
            .I(N__14140));
    InMux I__2706 (
            .O(N__14151),
            .I(N__14140));
    CascadeMux I__2705 (
            .O(N__14150),
            .I(N__14137));
    CascadeMux I__2704 (
            .O(N__14149),
            .I(N__14134));
    LocalMux I__2703 (
            .O(N__14140),
            .I(N__14130));
    InMux I__2702 (
            .O(N__14137),
            .I(N__14123));
    InMux I__2701 (
            .O(N__14134),
            .I(N__14123));
    InMux I__2700 (
            .O(N__14133),
            .I(N__14123));
    Span4Mux_h I__2699 (
            .O(N__14130),
            .I(N__14118));
    LocalMux I__2698 (
            .O(N__14123),
            .I(N__14118));
    Odrv4 I__2697 (
            .O(N__14118),
            .I(\Lab_UT.min2_1 ));
    CascadeMux I__2696 (
            .O(N__14115),
            .I(N__14106));
    CascadeMux I__2695 (
            .O(N__14114),
            .I(N__14103));
    CascadeMux I__2694 (
            .O(N__14113),
            .I(N__14100));
    CascadeMux I__2693 (
            .O(N__14112),
            .I(N__14097));
    CascadeMux I__2692 (
            .O(N__14111),
            .I(N__14094));
    CascadeMux I__2691 (
            .O(N__14110),
            .I(N__14091));
    CascadeMux I__2690 (
            .O(N__14109),
            .I(N__14088));
    InMux I__2689 (
            .O(N__14106),
            .I(N__14085));
    InMux I__2688 (
            .O(N__14103),
            .I(N__14076));
    InMux I__2687 (
            .O(N__14100),
            .I(N__14076));
    InMux I__2686 (
            .O(N__14097),
            .I(N__14076));
    InMux I__2685 (
            .O(N__14094),
            .I(N__14076));
    InMux I__2684 (
            .O(N__14091),
            .I(N__14071));
    InMux I__2683 (
            .O(N__14088),
            .I(N__14071));
    LocalMux I__2682 (
            .O(N__14085),
            .I(\Lab_UT.sec1_3 ));
    LocalMux I__2681 (
            .O(N__14076),
            .I(\Lab_UT.sec1_3 ));
    LocalMux I__2680 (
            .O(N__14071),
            .I(\Lab_UT.sec1_3 ));
    InMux I__2679 (
            .O(N__14064),
            .I(N__14055));
    InMux I__2678 (
            .O(N__14063),
            .I(N__14042));
    InMux I__2677 (
            .O(N__14062),
            .I(N__14042));
    InMux I__2676 (
            .O(N__14061),
            .I(N__14042));
    InMux I__2675 (
            .O(N__14060),
            .I(N__14042));
    InMux I__2674 (
            .O(N__14059),
            .I(N__14042));
    InMux I__2673 (
            .O(N__14058),
            .I(N__14042));
    LocalMux I__2672 (
            .O(N__14055),
            .I(\Lab_UT.sec1_0 ));
    LocalMux I__2671 (
            .O(N__14042),
            .I(\Lab_UT.sec1_0 ));
    InMux I__2670 (
            .O(N__14037),
            .I(N__14034));
    LocalMux I__2669 (
            .O(N__14034),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__2668 (
            .O(N__14031),
            .I(N__14028));
    LocalMux I__2667 (
            .O(N__14028),
            .I(\uu2.bitmapZ0Z_212 ));
    InMux I__2666 (
            .O(N__14025),
            .I(N__14022));
    LocalMux I__2665 (
            .O(N__14022),
            .I(\uu2.bitmap_pmux_17_ns_1 ));
    CascadeMux I__2664 (
            .O(N__14019),
            .I(N__14014));
    CascadeMux I__2663 (
            .O(N__14018),
            .I(N__14011));
    InMux I__2662 (
            .O(N__14017),
            .I(N__14004));
    InMux I__2661 (
            .O(N__14014),
            .I(N__14004));
    InMux I__2660 (
            .O(N__14011),
            .I(N__14004));
    LocalMux I__2659 (
            .O(N__14004),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__2658 (
            .O(N__14001),
            .I(N__13998));
    LocalMux I__2657 (
            .O(N__13998),
            .I(N__13995));
    Span4Mux_h I__2656 (
            .O(N__13995),
            .I(N__13992));
    Odrv4 I__2655 (
            .O(N__13992),
            .I(\uu2.bitmap_pmux_16_ns_1 ));
    InMux I__2654 (
            .O(N__13989),
            .I(N__13986));
    LocalMux I__2653 (
            .O(N__13986),
            .I(\uu2.bitmapZ0Z_72 ));
    InMux I__2652 (
            .O(N__13983),
            .I(N__13980));
    LocalMux I__2651 (
            .O(N__13980),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__2650 (
            .O(N__13977),
            .I(N__13965));
    InMux I__2649 (
            .O(N__13976),
            .I(N__13965));
    InMux I__2648 (
            .O(N__13975),
            .I(N__13965));
    InMux I__2647 (
            .O(N__13974),
            .I(N__13965));
    LocalMux I__2646 (
            .O(N__13965),
            .I(N__13959));
    InMux I__2645 (
            .O(N__13964),
            .I(N__13952));
    InMux I__2644 (
            .O(N__13963),
            .I(N__13952));
    InMux I__2643 (
            .O(N__13962),
            .I(N__13952));
    Odrv12 I__2642 (
            .O(N__13959),
            .I(\Lab_UT.min2_0 ));
    LocalMux I__2641 (
            .O(N__13952),
            .I(\Lab_UT.min2_0 ));
    CascadeMux I__2640 (
            .O(N__13947),
            .I(N__13942));
    CascadeMux I__2639 (
            .O(N__13946),
            .I(N__13937));
    CascadeMux I__2638 (
            .O(N__13945),
            .I(N__13932));
    InMux I__2637 (
            .O(N__13942),
            .I(N__13923));
    InMux I__2636 (
            .O(N__13941),
            .I(N__13923));
    InMux I__2635 (
            .O(N__13940),
            .I(N__13923));
    InMux I__2634 (
            .O(N__13937),
            .I(N__13923));
    InMux I__2633 (
            .O(N__13936),
            .I(N__13916));
    InMux I__2632 (
            .O(N__13935),
            .I(N__13916));
    InMux I__2631 (
            .O(N__13932),
            .I(N__13916));
    LocalMux I__2630 (
            .O(N__13923),
            .I(\Lab_UT.min2_3 ));
    LocalMux I__2629 (
            .O(N__13916),
            .I(\Lab_UT.min2_3 ));
    InMux I__2628 (
            .O(N__13911),
            .I(N__13899));
    InMux I__2627 (
            .O(N__13910),
            .I(N__13899));
    InMux I__2626 (
            .O(N__13909),
            .I(N__13899));
    InMux I__2625 (
            .O(N__13908),
            .I(N__13899));
    LocalMux I__2624 (
            .O(N__13899),
            .I(N__13893));
    InMux I__2623 (
            .O(N__13898),
            .I(N__13886));
    InMux I__2622 (
            .O(N__13897),
            .I(N__13886));
    InMux I__2621 (
            .O(N__13896),
            .I(N__13886));
    Odrv4 I__2620 (
            .O(N__13893),
            .I(\Lab_UT.min2_2 ));
    LocalMux I__2619 (
            .O(N__13886),
            .I(\Lab_UT.min2_2 ));
    InMux I__2618 (
            .O(N__13881),
            .I(N__13878));
    LocalMux I__2617 (
            .O(N__13878),
            .I(N__13875));
    Odrv4 I__2616 (
            .O(N__13875),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__2615 (
            .O(N__13872),
            .I(N__13866));
    InMux I__2614 (
            .O(N__13871),
            .I(N__13858));
    InMux I__2613 (
            .O(N__13870),
            .I(N__13858));
    InMux I__2612 (
            .O(N__13869),
            .I(N__13858));
    LocalMux I__2611 (
            .O(N__13866),
            .I(N__13855));
    InMux I__2610 (
            .O(N__13865),
            .I(N__13850));
    LocalMux I__2609 (
            .O(N__13858),
            .I(N__13845));
    Span4Mux_v I__2608 (
            .O(N__13855),
            .I(N__13845));
    InMux I__2607 (
            .O(N__13854),
            .I(N__13840));
    InMux I__2606 (
            .O(N__13853),
            .I(N__13840));
    LocalMux I__2605 (
            .O(N__13850),
            .I(\Lab_UT.di_Stens_1 ));
    Odrv4 I__2604 (
            .O(N__13845),
            .I(\Lab_UT.di_Stens_1 ));
    LocalMux I__2603 (
            .O(N__13840),
            .I(\Lab_UT.di_Stens_1 ));
    InMux I__2602 (
            .O(N__13833),
            .I(N__13818));
    InMux I__2601 (
            .O(N__13832),
            .I(N__13818));
    InMux I__2600 (
            .O(N__13831),
            .I(N__13818));
    InMux I__2599 (
            .O(N__13830),
            .I(N__13818));
    InMux I__2598 (
            .O(N__13829),
            .I(N__13813));
    InMux I__2597 (
            .O(N__13828),
            .I(N__13813));
    InMux I__2596 (
            .O(N__13827),
            .I(N__13810));
    LocalMux I__2595 (
            .O(N__13818),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__2594 (
            .O(N__13813),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__2593 (
            .O(N__13810),
            .I(\Lab_UT.sec1_1 ));
    InMux I__2592 (
            .O(N__13803),
            .I(N__13800));
    LocalMux I__2591 (
            .O(N__13800),
            .I(\uu2.bitmapZ0Z_290 ));
    InMux I__2590 (
            .O(N__13797),
            .I(N__13794));
    LocalMux I__2589 (
            .O(N__13794),
            .I(\uu2.bitmapZ0Z_34 ));
    CascadeMux I__2588 (
            .O(N__13791),
            .I(N__13786));
    CascadeMux I__2587 (
            .O(N__13790),
            .I(N__13783));
    CascadeMux I__2586 (
            .O(N__13789),
            .I(N__13779));
    InMux I__2585 (
            .O(N__13786),
            .I(N__13774));
    InMux I__2584 (
            .O(N__13783),
            .I(N__13771));
    InMux I__2583 (
            .O(N__13782),
            .I(N__13766));
    InMux I__2582 (
            .O(N__13779),
            .I(N__13766));
    InMux I__2581 (
            .O(N__13778),
            .I(N__13761));
    InMux I__2580 (
            .O(N__13777),
            .I(N__13761));
    LocalMux I__2579 (
            .O(N__13774),
            .I(N__13758));
    LocalMux I__2578 (
            .O(N__13771),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2577 (
            .O(N__13766),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2576 (
            .O(N__13761),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__2575 (
            .O(N__13758),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    InMux I__2574 (
            .O(N__13749),
            .I(N__13746));
    LocalMux I__2573 (
            .O(N__13746),
            .I(\uu2.bitmap_pmux_26_bm_1 ));
    InMux I__2572 (
            .O(N__13743),
            .I(N__13740));
    LocalMux I__2571 (
            .O(N__13740),
            .I(N__13737));
    Odrv4 I__2570 (
            .O(N__13737),
            .I(\uu2.bitmap_RNIP2JO1Z0Z_34 ));
    InMux I__2569 (
            .O(N__13734),
            .I(N__13731));
    LocalMux I__2568 (
            .O(N__13731),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__2567 (
            .O(N__13728),
            .I(N__13722));
    InMux I__2566 (
            .O(N__13727),
            .I(N__13714));
    InMux I__2565 (
            .O(N__13726),
            .I(N__13714));
    InMux I__2564 (
            .O(N__13725),
            .I(N__13714));
    LocalMux I__2563 (
            .O(N__13722),
            .I(N__13711));
    CascadeMux I__2562 (
            .O(N__13721),
            .I(N__13706));
    LocalMux I__2561 (
            .O(N__13714),
            .I(N__13703));
    Span12Mux_s6_v I__2560 (
            .O(N__13711),
            .I(N__13700));
    InMux I__2559 (
            .O(N__13710),
            .I(N__13693));
    InMux I__2558 (
            .O(N__13709),
            .I(N__13693));
    InMux I__2557 (
            .O(N__13706),
            .I(N__13693));
    Odrv4 I__2556 (
            .O(N__13703),
            .I(\Lab_UT.di_Sones_3 ));
    Odrv12 I__2555 (
            .O(N__13700),
            .I(\Lab_UT.di_Sones_3 ));
    LocalMux I__2554 (
            .O(N__13693),
            .I(\Lab_UT.di_Sones_3 ));
    CascadeMux I__2553 (
            .O(N__13686),
            .I(N__13683));
    InMux I__2552 (
            .O(N__13683),
            .I(N__13679));
    InMux I__2551 (
            .O(N__13682),
            .I(N__13676));
    LocalMux I__2550 (
            .O(N__13679),
            .I(N__13672));
    LocalMux I__2549 (
            .O(N__13676),
            .I(N__13669));
    InMux I__2548 (
            .O(N__13675),
            .I(N__13666));
    Span4Mux_h I__2547 (
            .O(N__13672),
            .I(N__13663));
    Span4Mux_v I__2546 (
            .O(N__13669),
            .I(N__13660));
    LocalMux I__2545 (
            .O(N__13666),
            .I(N__13657));
    Odrv4 I__2544 (
            .O(N__13663),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__2543 (
            .O(N__13660),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__2542 (
            .O(N__13657),
            .I(\Lab_UT.di_ASones_3 ));
    InMux I__2541 (
            .O(N__13650),
            .I(N__13646));
    InMux I__2540 (
            .O(N__13649),
            .I(N__13643));
    LocalMux I__2539 (
            .O(N__13646),
            .I(N__13640));
    LocalMux I__2538 (
            .O(N__13643),
            .I(N__13637));
    Span4Mux_h I__2537 (
            .O(N__13640),
            .I(N__13632));
    Span4Mux_s2_v I__2536 (
            .O(N__13637),
            .I(N__13632));
    Span4Mux_v I__2535 (
            .O(N__13632),
            .I(N__13628));
    InMux I__2534 (
            .O(N__13631),
            .I(N__13625));
    Odrv4 I__2533 (
            .O(N__13628),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__2532 (
            .O(N__13625),
            .I(\Lab_UT.di_ASones_0 ));
    InMux I__2531 (
            .O(N__13620),
            .I(N__13616));
    InMux I__2530 (
            .O(N__13619),
            .I(N__13613));
    LocalMux I__2529 (
            .O(N__13616),
            .I(N__13609));
    LocalMux I__2528 (
            .O(N__13613),
            .I(N__13606));
    InMux I__2527 (
            .O(N__13612),
            .I(N__13603));
    Span4Mux_v I__2526 (
            .O(N__13609),
            .I(N__13600));
    Span4Mux_v I__2525 (
            .O(N__13606),
            .I(N__13597));
    LocalMux I__2524 (
            .O(N__13603),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__2523 (
            .O(N__13600),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__2522 (
            .O(N__13597),
            .I(\Lab_UT.di_AMones_3 ));
    InMux I__2521 (
            .O(N__13590),
            .I(N__13586));
    InMux I__2520 (
            .O(N__13589),
            .I(N__13583));
    LocalMux I__2519 (
            .O(N__13586),
            .I(N__13580));
    LocalMux I__2518 (
            .O(N__13583),
            .I(N__13576));
    Span4Mux_h I__2517 (
            .O(N__13580),
            .I(N__13573));
    InMux I__2516 (
            .O(N__13579),
            .I(N__13570));
    Odrv4 I__2515 (
            .O(N__13576),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__2514 (
            .O(N__13573),
            .I(\Lab_UT.di_AMtens_0 ));
    LocalMux I__2513 (
            .O(N__13570),
            .I(\Lab_UT.di_AMtens_0 ));
    InMux I__2512 (
            .O(N__13563),
            .I(N__13554));
    InMux I__2511 (
            .O(N__13562),
            .I(N__13541));
    InMux I__2510 (
            .O(N__13561),
            .I(N__13541));
    InMux I__2509 (
            .O(N__13560),
            .I(N__13541));
    InMux I__2508 (
            .O(N__13559),
            .I(N__13541));
    InMux I__2507 (
            .O(N__13558),
            .I(N__13541));
    InMux I__2506 (
            .O(N__13557),
            .I(N__13541));
    LocalMux I__2505 (
            .O(N__13554),
            .I(\Lab_UT.min1_0 ));
    LocalMux I__2504 (
            .O(N__13541),
            .I(\Lab_UT.min1_0 ));
    InMux I__2503 (
            .O(N__13536),
            .I(N__13531));
    InMux I__2502 (
            .O(N__13535),
            .I(N__13526));
    InMux I__2501 (
            .O(N__13534),
            .I(N__13526));
    LocalMux I__2500 (
            .O(N__13531),
            .I(N__13523));
    LocalMux I__2499 (
            .O(N__13526),
            .I(N__13520));
    Span4Mux_h I__2498 (
            .O(N__13523),
            .I(N__13517));
    Span4Mux_h I__2497 (
            .O(N__13520),
            .I(N__13514));
    Odrv4 I__2496 (
            .O(N__13517),
            .I(\Lab_UT.di_AMtens_3 ));
    Odrv4 I__2495 (
            .O(N__13514),
            .I(\Lab_UT.di_AMtens_3 ));
    InMux I__2494 (
            .O(N__13509),
            .I(N__13505));
    InMux I__2493 (
            .O(N__13508),
            .I(N__13502));
    LocalMux I__2492 (
            .O(N__13505),
            .I(N__13499));
    LocalMux I__2491 (
            .O(N__13502),
            .I(N__13492));
    Span4Mux_h I__2490 (
            .O(N__13499),
            .I(N__13492));
    InMux I__2489 (
            .O(N__13498),
            .I(N__13486));
    InMux I__2488 (
            .O(N__13497),
            .I(N__13486));
    Span4Mux_v I__2487 (
            .O(N__13492),
            .I(N__13483));
    InMux I__2486 (
            .O(N__13491),
            .I(N__13480));
    LocalMux I__2485 (
            .O(N__13486),
            .I(\Lab_UT.di_Mtens_3 ));
    Odrv4 I__2484 (
            .O(N__13483),
            .I(\Lab_UT.di_Mtens_3 ));
    LocalMux I__2483 (
            .O(N__13480),
            .I(\Lab_UT.di_Mtens_3 ));
    CascadeMux I__2482 (
            .O(N__13473),
            .I(N__13470));
    InMux I__2481 (
            .O(N__13470),
            .I(N__13464));
    CascadeMux I__2480 (
            .O(N__13469),
            .I(N__13460));
    CascadeMux I__2479 (
            .O(N__13468),
            .I(N__13456));
    CascadeMux I__2478 (
            .O(N__13467),
            .I(N__13452));
    LocalMux I__2477 (
            .O(N__13464),
            .I(N__13449));
    InMux I__2476 (
            .O(N__13463),
            .I(N__13436));
    InMux I__2475 (
            .O(N__13460),
            .I(N__13436));
    InMux I__2474 (
            .O(N__13459),
            .I(N__13436));
    InMux I__2473 (
            .O(N__13456),
            .I(N__13436));
    InMux I__2472 (
            .O(N__13455),
            .I(N__13436));
    InMux I__2471 (
            .O(N__13452),
            .I(N__13436));
    Odrv4 I__2470 (
            .O(N__13449),
            .I(\Lab_UT.min1_3 ));
    LocalMux I__2469 (
            .O(N__13436),
            .I(\Lab_UT.min1_3 ));
    CascadeMux I__2468 (
            .O(N__13431),
            .I(N__13428));
    InMux I__2467 (
            .O(N__13428),
            .I(N__13423));
    CascadeMux I__2466 (
            .O(N__13427),
            .I(N__13419));
    CascadeMux I__2465 (
            .O(N__13426),
            .I(N__13414));
    LocalMux I__2464 (
            .O(N__13423),
            .I(N__13410));
    InMux I__2463 (
            .O(N__13422),
            .I(N__13397));
    InMux I__2462 (
            .O(N__13419),
            .I(N__13397));
    InMux I__2461 (
            .O(N__13418),
            .I(N__13397));
    InMux I__2460 (
            .O(N__13417),
            .I(N__13397));
    InMux I__2459 (
            .O(N__13414),
            .I(N__13397));
    InMux I__2458 (
            .O(N__13413),
            .I(N__13397));
    Span4Mux_s2_v I__2457 (
            .O(N__13410),
            .I(N__13394));
    LocalMux I__2456 (
            .O(N__13397),
            .I(N__13391));
    Odrv4 I__2455 (
            .O(N__13394),
            .I(\uu2.N_37 ));
    Odrv4 I__2454 (
            .O(N__13391),
            .I(\uu2.N_37 ));
    InMux I__2453 (
            .O(N__13386),
            .I(N__13377));
    InMux I__2452 (
            .O(N__13385),
            .I(N__13377));
    InMux I__2451 (
            .O(N__13384),
            .I(N__13374));
    InMux I__2450 (
            .O(N__13383),
            .I(N__13366));
    InMux I__2449 (
            .O(N__13382),
            .I(N__13363));
    LocalMux I__2448 (
            .O(N__13377),
            .I(N__13360));
    LocalMux I__2447 (
            .O(N__13374),
            .I(N__13357));
    InMux I__2446 (
            .O(N__13373),
            .I(N__13350));
    InMux I__2445 (
            .O(N__13372),
            .I(N__13350));
    InMux I__2444 (
            .O(N__13371),
            .I(N__13350));
    InMux I__2443 (
            .O(N__13370),
            .I(N__13345));
    InMux I__2442 (
            .O(N__13369),
            .I(N__13345));
    LocalMux I__2441 (
            .O(N__13366),
            .I(N__13342));
    LocalMux I__2440 (
            .O(N__13363),
            .I(N__13339));
    Span4Mux_h I__2439 (
            .O(N__13360),
            .I(N__13336));
    Odrv12 I__2438 (
            .O(N__13357),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2437 (
            .O(N__13350),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__2436 (
            .O(N__13345),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2435 (
            .O(N__13342),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2434 (
            .O(N__13339),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__2433 (
            .O(N__13336),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__2432 (
            .O(N__13323),
            .I(N__13320));
    InMux I__2431 (
            .O(N__13320),
            .I(N__13317));
    LocalMux I__2430 (
            .O(N__13317),
            .I(\uu2.N_45 ));
    InMux I__2429 (
            .O(N__13314),
            .I(N__13311));
    LocalMux I__2428 (
            .O(N__13311),
            .I(N__13308));
    Odrv4 I__2427 (
            .O(N__13308),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    CascadeMux I__2426 (
            .O(N__13305),
            .I(N__13301));
    InMux I__2425 (
            .O(N__13304),
            .I(N__13298));
    InMux I__2424 (
            .O(N__13301),
            .I(N__13290));
    LocalMux I__2423 (
            .O(N__13298),
            .I(N__13287));
    InMux I__2422 (
            .O(N__13297),
            .I(N__13282));
    InMux I__2421 (
            .O(N__13296),
            .I(N__13282));
    InMux I__2420 (
            .O(N__13295),
            .I(N__13275));
    InMux I__2419 (
            .O(N__13294),
            .I(N__13275));
    InMux I__2418 (
            .O(N__13293),
            .I(N__13275));
    LocalMux I__2417 (
            .O(N__13290),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv12 I__2416 (
            .O(N__13287),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2415 (
            .O(N__13282),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__2414 (
            .O(N__13275),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    InMux I__2413 (
            .O(N__13266),
            .I(N__13257));
    InMux I__2412 (
            .O(N__13265),
            .I(N__13257));
    InMux I__2411 (
            .O(N__13264),
            .I(N__13253));
    InMux I__2410 (
            .O(N__13263),
            .I(N__13250));
    InMux I__2409 (
            .O(N__13262),
            .I(N__13246));
    LocalMux I__2408 (
            .O(N__13257),
            .I(N__13243));
    CascadeMux I__2407 (
            .O(N__13256),
            .I(N__13237));
    LocalMux I__2406 (
            .O(N__13253),
            .I(N__13234));
    LocalMux I__2405 (
            .O(N__13250),
            .I(N__13231));
    InMux I__2404 (
            .O(N__13249),
            .I(N__13228));
    LocalMux I__2403 (
            .O(N__13246),
            .I(N__13225));
    Span4Mux_h I__2402 (
            .O(N__13243),
            .I(N__13222));
    InMux I__2401 (
            .O(N__13242),
            .I(N__13213));
    InMux I__2400 (
            .O(N__13241),
            .I(N__13213));
    InMux I__2399 (
            .O(N__13240),
            .I(N__13213));
    InMux I__2398 (
            .O(N__13237),
            .I(N__13213));
    Span4Mux_h I__2397 (
            .O(N__13234),
            .I(N__13208));
    Span4Mux_h I__2396 (
            .O(N__13231),
            .I(N__13208));
    LocalMux I__2395 (
            .O(N__13228),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv12 I__2394 (
            .O(N__13225),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2393 (
            .O(N__13222),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2392 (
            .O(N__13213),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2391 (
            .O(N__13208),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    InMux I__2390 (
            .O(N__13197),
            .I(N__13194));
    LocalMux I__2389 (
            .O(N__13194),
            .I(N__13190));
    CascadeMux I__2388 (
            .O(N__13193),
            .I(N__13185));
    Span4Mux_h I__2387 (
            .O(N__13190),
            .I(N__13180));
    InMux I__2386 (
            .O(N__13189),
            .I(N__13173));
    InMux I__2385 (
            .O(N__13188),
            .I(N__13173));
    InMux I__2384 (
            .O(N__13185),
            .I(N__13173));
    InMux I__2383 (
            .O(N__13184),
            .I(N__13168));
    InMux I__2382 (
            .O(N__13183),
            .I(N__13168));
    Odrv4 I__2381 (
            .O(N__13180),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2380 (
            .O(N__13173),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__2379 (
            .O(N__13168),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__2378 (
            .O(N__13161),
            .I(N__13158));
    LocalMux I__2377 (
            .O(N__13158),
            .I(N__13155));
    Span4Mux_h I__2376 (
            .O(N__13155),
            .I(N__13152));
    Odrv4 I__2375 (
            .O(N__13152),
            .I(\uu2.bitmap_pmux_sn_N_36 ));
    InMux I__2374 (
            .O(N__13149),
            .I(N__13146));
    LocalMux I__2373 (
            .O(N__13146),
            .I(\uu2.bitmapZ0Z_194 ));
    InMux I__2372 (
            .O(N__13143),
            .I(N__13140));
    LocalMux I__2371 (
            .O(N__13140),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__2370 (
            .O(N__13137),
            .I(N__13134));
    LocalMux I__2369 (
            .O(N__13134),
            .I(\uu2.bitmap_pmux_20_ns_1 ));
    InMux I__2368 (
            .O(N__13131),
            .I(N__13128));
    LocalMux I__2367 (
            .O(N__13128),
            .I(\uu2.bitmapZ0Z_162 ));
    CascadeMux I__2366 (
            .O(N__13125),
            .I(\Lab_UT.dictrl.g1_1_4_cascade_ ));
    InMux I__2365 (
            .O(N__13122),
            .I(N__13119));
    LocalMux I__2364 (
            .O(N__13119),
            .I(N__13116));
    Odrv4 I__2363 (
            .O(N__13116),
            .I(\Lab_UT.dictrl.g1_1Z0Z_5 ));
    CascadeMux I__2362 (
            .O(N__13113),
            .I(N__13108));
    CascadeMux I__2361 (
            .O(N__13112),
            .I(N__13105));
    InMux I__2360 (
            .O(N__13111),
            .I(N__13094));
    InMux I__2359 (
            .O(N__13108),
            .I(N__13094));
    InMux I__2358 (
            .O(N__13105),
            .I(N__13084));
    InMux I__2357 (
            .O(N__13104),
            .I(N__13084));
    InMux I__2356 (
            .O(N__13103),
            .I(N__13084));
    InMux I__2355 (
            .O(N__13102),
            .I(N__13081));
    InMux I__2354 (
            .O(N__13101),
            .I(N__13078));
    InMux I__2353 (
            .O(N__13100),
            .I(N__13073));
    InMux I__2352 (
            .O(N__13099),
            .I(N__13073));
    LocalMux I__2351 (
            .O(N__13094),
            .I(N__13070));
    InMux I__2350 (
            .O(N__13093),
            .I(N__13065));
    InMux I__2349 (
            .O(N__13092),
            .I(N__13065));
    InMux I__2348 (
            .O(N__13091),
            .I(N__13062));
    LocalMux I__2347 (
            .O(N__13084),
            .I(N__13059));
    LocalMux I__2346 (
            .O(N__13081),
            .I(N__13054));
    LocalMux I__2345 (
            .O(N__13078),
            .I(N__13054));
    LocalMux I__2344 (
            .O(N__13073),
            .I(N__13049));
    Span4Mux_v I__2343 (
            .O(N__13070),
            .I(N__13049));
    LocalMux I__2342 (
            .O(N__13065),
            .I(N__13042));
    LocalMux I__2341 (
            .O(N__13062),
            .I(N__13042));
    Span4Mux_h I__2340 (
            .O(N__13059),
            .I(N__13042));
    Odrv4 I__2339 (
            .O(N__13054),
            .I(bu_rx_data_7));
    Odrv4 I__2338 (
            .O(N__13049),
            .I(bu_rx_data_7));
    Odrv4 I__2337 (
            .O(N__13042),
            .I(bu_rx_data_7));
    InMux I__2336 (
            .O(N__13035),
            .I(N__13029));
    InMux I__2335 (
            .O(N__13034),
            .I(N__13029));
    LocalMux I__2334 (
            .O(N__13029),
            .I(N__13025));
    InMux I__2333 (
            .O(N__13028),
            .I(N__13022));
    Span4Mux_h I__2332 (
            .O(N__13025),
            .I(N__13017));
    LocalMux I__2331 (
            .O(N__13022),
            .I(N__13017));
    Span4Mux_h I__2330 (
            .O(N__13017),
            .I(N__13013));
    InMux I__2329 (
            .O(N__13016),
            .I(N__13010));
    Span4Mux_v I__2328 (
            .O(N__13013),
            .I(N__13005));
    LocalMux I__2327 (
            .O(N__13010),
            .I(N__13005));
    Odrv4 I__2326 (
            .O(N__13005),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__2325 (
            .O(N__13002),
            .I(N__12996));
    InMux I__2324 (
            .O(N__13001),
            .I(N__12996));
    LocalMux I__2323 (
            .O(N__12996),
            .I(bu_rx_data_fast_7));
    InMux I__2322 (
            .O(N__12993),
            .I(N__12983));
    InMux I__2321 (
            .O(N__12992),
            .I(N__12983));
    InMux I__2320 (
            .O(N__12991),
            .I(N__12983));
    CascadeMux I__2319 (
            .O(N__12990),
            .I(N__12978));
    LocalMux I__2318 (
            .O(N__12983),
            .I(N__12975));
    InMux I__2317 (
            .O(N__12982),
            .I(N__12968));
    InMux I__2316 (
            .O(N__12981),
            .I(N__12968));
    InMux I__2315 (
            .O(N__12978),
            .I(N__12968));
    Span4Mux_h I__2314 (
            .O(N__12975),
            .I(N__12965));
    LocalMux I__2313 (
            .O(N__12968),
            .I(\uu2.N_40 ));
    Odrv4 I__2312 (
            .O(N__12965),
            .I(\uu2.N_40 ));
    CascadeMux I__2311 (
            .O(N__12960),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ));
    CascadeMux I__2310 (
            .O(N__12957),
            .I(\Lab_UT.dictrl.m22Z0Z_1_cascade_ ));
    InMux I__2309 (
            .O(N__12954),
            .I(N__12951));
    LocalMux I__2308 (
            .O(N__12951),
            .I(\Lab_UT.dictrl.N_72_mux_1 ));
    CascadeMux I__2307 (
            .O(N__12948),
            .I(N__12945));
    InMux I__2306 (
            .O(N__12945),
            .I(N__12942));
    LocalMux I__2305 (
            .O(N__12942),
            .I(\Lab_UT.dictrl.g1_1_0_0 ));
    InMux I__2304 (
            .O(N__12939),
            .I(N__12935));
    InMux I__2303 (
            .O(N__12938),
            .I(N__12932));
    LocalMux I__2302 (
            .O(N__12935),
            .I(N__12929));
    LocalMux I__2301 (
            .O(N__12932),
            .I(\Lab_UT.dictrl.m22Z0Z_1 ));
    Odrv4 I__2300 (
            .O(N__12929),
            .I(\Lab_UT.dictrl.m22Z0Z_1 ));
    InMux I__2299 (
            .O(N__12924),
            .I(N__12921));
    LocalMux I__2298 (
            .O(N__12921),
            .I(\Lab_UT.dictrl.g1_1_0 ));
    CascadeMux I__2297 (
            .O(N__12918),
            .I(N__12915));
    InMux I__2296 (
            .O(N__12915),
            .I(N__12912));
    LocalMux I__2295 (
            .O(N__12912),
            .I(N__12909));
    Odrv12 I__2294 (
            .O(N__12909),
            .I(\Lab_UT.dictrl.g1_rn_0 ));
    InMux I__2293 (
            .O(N__12906),
            .I(N__12903));
    LocalMux I__2292 (
            .O(N__12903),
            .I(N__12900));
    Span4Mux_v I__2291 (
            .O(N__12900),
            .I(N__12896));
    InMux I__2290 (
            .O(N__12899),
            .I(N__12893));
    Odrv4 I__2289 (
            .O(N__12896),
            .I(\Lab_UT.dictrl.m34Z0Z_1 ));
    LocalMux I__2288 (
            .O(N__12893),
            .I(\Lab_UT.dictrl.m34Z0Z_1 ));
    CascadeMux I__2287 (
            .O(N__12888),
            .I(N__12884));
    CascadeMux I__2286 (
            .O(N__12887),
            .I(N__12881));
    InMux I__2285 (
            .O(N__12884),
            .I(N__12878));
    InMux I__2284 (
            .O(N__12881),
            .I(N__12875));
    LocalMux I__2283 (
            .O(N__12878),
            .I(bu_rx_data_fast_3));
    LocalMux I__2282 (
            .O(N__12875),
            .I(bu_rx_data_fast_3));
    InMux I__2281 (
            .O(N__12870),
            .I(N__12864));
    InMux I__2280 (
            .O(N__12869),
            .I(N__12864));
    LocalMux I__2279 (
            .O(N__12864),
            .I(N__12861));
    Odrv4 I__2278 (
            .O(N__12861),
            .I(bu_rx_data_fast_0));
    CascadeMux I__2277 (
            .O(N__12858),
            .I(\Lab_UT.dictrl.m13_out_cascade_ ));
    CascadeMux I__2276 (
            .O(N__12855),
            .I(\Lab_UT.dictrl.N_18_0_0_cascade_ ));
    InMux I__2275 (
            .O(N__12852),
            .I(N__12849));
    LocalMux I__2274 (
            .O(N__12849),
            .I(\Lab_UT.dictrl.G_25_i_o3_5 ));
    InMux I__2273 (
            .O(N__12846),
            .I(N__12843));
    LocalMux I__2272 (
            .O(N__12843),
            .I(N__12840));
    Odrv4 I__2271 (
            .O(N__12840),
            .I(\Lab_UT.dictrl.G_25_i_o3_4 ));
    CascadeMux I__2270 (
            .O(N__12837),
            .I(\Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ));
    InMux I__2269 (
            .O(N__12834),
            .I(N__12831));
    LocalMux I__2268 (
            .O(N__12831),
            .I(\Lab_UT.dictrl.N_11 ));
    CascadeMux I__2267 (
            .O(N__12828),
            .I(\Lab_UT.dictrl.m34Z0Z_1_cascade_ ));
    InMux I__2266 (
            .O(N__12825),
            .I(N__12818));
    InMux I__2265 (
            .O(N__12824),
            .I(N__12813));
    InMux I__2264 (
            .O(N__12823),
            .I(N__12813));
    InMux I__2263 (
            .O(N__12822),
            .I(N__12801));
    InMux I__2262 (
            .O(N__12821),
            .I(N__12801));
    LocalMux I__2261 (
            .O(N__12818),
            .I(N__12798));
    LocalMux I__2260 (
            .O(N__12813),
            .I(N__12795));
    InMux I__2259 (
            .O(N__12812),
            .I(N__12790));
    InMux I__2258 (
            .O(N__12811),
            .I(N__12790));
    InMux I__2257 (
            .O(N__12810),
            .I(N__12785));
    InMux I__2256 (
            .O(N__12809),
            .I(N__12785));
    InMux I__2255 (
            .O(N__12808),
            .I(N__12778));
    InMux I__2254 (
            .O(N__12807),
            .I(N__12778));
    InMux I__2253 (
            .O(N__12806),
            .I(N__12778));
    LocalMux I__2252 (
            .O(N__12801),
            .I(bu_rx_data_6));
    Odrv4 I__2251 (
            .O(N__12798),
            .I(bu_rx_data_6));
    Odrv4 I__2250 (
            .O(N__12795),
            .I(bu_rx_data_6));
    LocalMux I__2249 (
            .O(N__12790),
            .I(bu_rx_data_6));
    LocalMux I__2248 (
            .O(N__12785),
            .I(bu_rx_data_6));
    LocalMux I__2247 (
            .O(N__12778),
            .I(bu_rx_data_6));
    CascadeMux I__2246 (
            .O(N__12765),
            .I(\Lab_UT.i8_mux_0_cascade_ ));
    CascadeMux I__2245 (
            .O(N__12762),
            .I(N__12759));
    InMux I__2244 (
            .O(N__12759),
            .I(N__12756));
    LocalMux I__2243 (
            .O(N__12756),
            .I(\Lab_UT.dictrl.g0_0_sn ));
    CascadeMux I__2242 (
            .O(N__12753),
            .I(\Lab_UT.dictrl.g1_1_0_1_cascade_ ));
    InMux I__2241 (
            .O(N__12750),
            .I(N__12747));
    LocalMux I__2240 (
            .O(N__12747),
            .I(\Lab_UT.g1 ));
    InMux I__2239 (
            .O(N__12744),
            .I(N__12741));
    LocalMux I__2238 (
            .O(N__12741),
            .I(\Lab_UT.dictrl.g0_0_rn_0 ));
    InMux I__2237 (
            .O(N__12738),
            .I(N__12735));
    LocalMux I__2236 (
            .O(N__12735),
            .I(N__12732));
    Odrv4 I__2235 (
            .O(N__12732),
            .I(\Lab_UT.dictrl.G_25_i_0 ));
    InMux I__2234 (
            .O(N__12729),
            .I(N__12726));
    LocalMux I__2233 (
            .O(N__12726),
            .I(\Lab_UT.dictrl.G_25_i_1 ));
    InMux I__2232 (
            .O(N__12723),
            .I(N__12720));
    LocalMux I__2231 (
            .O(N__12720),
            .I(N__12717));
    Odrv4 I__2230 (
            .O(N__12717),
            .I(\Lab_UT.dictrl.g2Z0Z_0 ));
    CascadeMux I__2229 (
            .O(N__12714),
            .I(N__12711));
    InMux I__2228 (
            .O(N__12711),
            .I(N__12708));
    LocalMux I__2227 (
            .O(N__12708),
            .I(\Lab_UT.dictrl.g0_6_3_0 ));
    CEMux I__2226 (
            .O(N__12705),
            .I(N__12702));
    LocalMux I__2225 (
            .O(N__12702),
            .I(N__12699));
    Span4Mux_v I__2224 (
            .O(N__12699),
            .I(N__12696));
    Odrv4 I__2223 (
            .O(N__12696),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    CascadeMux I__2222 (
            .O(N__12693),
            .I(\Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_ ));
    CascadeMux I__2221 (
            .O(N__12690),
            .I(\Lab_UT.dictrl.G_25_i_a5_1_0_cascade_ ));
    InMux I__2220 (
            .O(N__12687),
            .I(N__12684));
    LocalMux I__2219 (
            .O(N__12684),
            .I(N__12681));
    Span4Mux_v I__2218 (
            .O(N__12681),
            .I(N__12678));
    Odrv4 I__2217 (
            .O(N__12678),
            .I(\Lab_UT.didp.N_90 ));
    InMux I__2216 (
            .O(N__12675),
            .I(N__12672));
    LocalMux I__2215 (
            .O(N__12672),
            .I(\Lab_UT.LdSones_i_4 ));
    InMux I__2214 (
            .O(N__12669),
            .I(N__12666));
    LocalMux I__2213 (
            .O(N__12666),
            .I(N__12663));
    Span4Mux_h I__2212 (
            .O(N__12663),
            .I(N__12660));
    Odrv4 I__2211 (
            .O(N__12660),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__2210 (
            .O(N__12657),
            .I(N__12648));
    InMux I__2209 (
            .O(N__12656),
            .I(N__12648));
    InMux I__2208 (
            .O(N__12655),
            .I(N__12648));
    LocalMux I__2207 (
            .O(N__12648),
            .I(N__12642));
    InMux I__2206 (
            .O(N__12647),
            .I(N__12637));
    InMux I__2205 (
            .O(N__12646),
            .I(N__12637));
    InMux I__2204 (
            .O(N__12645),
            .I(N__12634));
    Odrv4 I__2203 (
            .O(N__12642),
            .I(\Lab_UT.state_ret_8_ess ));
    LocalMux I__2202 (
            .O(N__12637),
            .I(\Lab_UT.state_ret_8_ess ));
    LocalMux I__2201 (
            .O(N__12634),
            .I(\Lab_UT.state_ret_8_ess ));
    CascadeMux I__2200 (
            .O(N__12627),
            .I(N__12621));
    CascadeMux I__2199 (
            .O(N__12626),
            .I(N__12617));
    CascadeMux I__2198 (
            .O(N__12625),
            .I(N__12612));
    CascadeMux I__2197 (
            .O(N__12624),
            .I(N__12609));
    InMux I__2196 (
            .O(N__12621),
            .I(N__12604));
    InMux I__2195 (
            .O(N__12620),
            .I(N__12604));
    InMux I__2194 (
            .O(N__12617),
            .I(N__12601));
    InMux I__2193 (
            .O(N__12616),
            .I(N__12598));
    InMux I__2192 (
            .O(N__12615),
            .I(N__12591));
    InMux I__2191 (
            .O(N__12612),
            .I(N__12591));
    InMux I__2190 (
            .O(N__12609),
            .I(N__12591));
    LocalMux I__2189 (
            .O(N__12604),
            .I(N__12586));
    LocalMux I__2188 (
            .O(N__12601),
            .I(N__12586));
    LocalMux I__2187 (
            .O(N__12598),
            .I(\Lab_UT.di_Stens_0 ));
    LocalMux I__2186 (
            .O(N__12591),
            .I(\Lab_UT.di_Stens_0 ));
    Odrv4 I__2185 (
            .O(N__12586),
            .I(\Lab_UT.di_Stens_0 ));
    CascadeMux I__2184 (
            .O(N__12579),
            .I(N__12576));
    InMux I__2183 (
            .O(N__12576),
            .I(N__12573));
    LocalMux I__2182 (
            .O(N__12573),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ));
    InMux I__2181 (
            .O(N__12570),
            .I(N__12567));
    LocalMux I__2180 (
            .O(N__12567),
            .I(\Lab_UT.didp.countrce1.q_5_1 ));
    InMux I__2179 (
            .O(N__12564),
            .I(N__12560));
    CascadeMux I__2178 (
            .O(N__12563),
            .I(N__12555));
    LocalMux I__2177 (
            .O(N__12560),
            .I(N__12552));
    InMux I__2176 (
            .O(N__12559),
            .I(N__12549));
    InMux I__2175 (
            .O(N__12558),
            .I(N__12546));
    InMux I__2174 (
            .O(N__12555),
            .I(N__12543));
    Span4Mux_v I__2173 (
            .O(N__12552),
            .I(N__12539));
    LocalMux I__2172 (
            .O(N__12549),
            .I(N__12532));
    LocalMux I__2171 (
            .O(N__12546),
            .I(N__12532));
    LocalMux I__2170 (
            .O(N__12543),
            .I(N__12532));
    InMux I__2169 (
            .O(N__12542),
            .I(N__12529));
    Odrv4 I__2168 (
            .O(N__12539),
            .I(\Lab_UT.dispString.N_143 ));
    Odrv4 I__2167 (
            .O(N__12532),
            .I(\Lab_UT.dispString.N_143 ));
    LocalMux I__2166 (
            .O(N__12529),
            .I(\Lab_UT.dispString.N_143 ));
    InMux I__2165 (
            .O(N__12522),
            .I(N__12519));
    LocalMux I__2164 (
            .O(N__12519),
            .I(N__12514));
    InMux I__2163 (
            .O(N__12518),
            .I(N__12511));
    InMux I__2162 (
            .O(N__12517),
            .I(N__12508));
    Span4Mux_v I__2161 (
            .O(N__12514),
            .I(N__12503));
    LocalMux I__2160 (
            .O(N__12511),
            .I(N__12503));
    LocalMux I__2159 (
            .O(N__12508),
            .I(N__12500));
    Odrv4 I__2158 (
            .O(N__12503),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__2157 (
            .O(N__12500),
            .I(\Lab_UT.di_AMones_0 ));
    InMux I__2156 (
            .O(N__12495),
            .I(N__12492));
    LocalMux I__2155 (
            .O(N__12492),
            .I(N__12489));
    Span4Mux_h I__2154 (
            .O(N__12489),
            .I(N__12486));
    Odrv4 I__2153 (
            .O(N__12486),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_0 ));
    InMux I__2152 (
            .O(N__12483),
            .I(N__12477));
    InMux I__2151 (
            .O(N__12482),
            .I(N__12477));
    LocalMux I__2150 (
            .O(N__12477),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    InMux I__2149 (
            .O(N__12474),
            .I(N__12471));
    LocalMux I__2148 (
            .O(N__12471),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_2 ));
    CascadeMux I__2147 (
            .O(N__12468),
            .I(\Lab_UT.didp.un1_dicLdStens_0_cascade_ ));
    CascadeMux I__2146 (
            .O(N__12465),
            .I(N__12460));
    InMux I__2145 (
            .O(N__12464),
            .I(N__12454));
    InMux I__2144 (
            .O(N__12463),
            .I(N__12454));
    InMux I__2143 (
            .O(N__12460),
            .I(N__12449));
    InMux I__2142 (
            .O(N__12459),
            .I(N__12449));
    LocalMux I__2141 (
            .O(N__12454),
            .I(N__12446));
    LocalMux I__2140 (
            .O(N__12449),
            .I(N__12443));
    Span4Mux_v I__2139 (
            .O(N__12446),
            .I(N__12440));
    Span4Mux_h I__2138 (
            .O(N__12443),
            .I(N__12437));
    Odrv4 I__2137 (
            .O(N__12440),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    Odrv4 I__2136 (
            .O(N__12437),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    InMux I__2135 (
            .O(N__12432),
            .I(N__12426));
    InMux I__2134 (
            .O(N__12431),
            .I(N__12426));
    LocalMux I__2133 (
            .O(N__12426),
            .I(N__12423));
    Odrv4 I__2132 (
            .O(N__12423),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__2131 (
            .O(N__12420),
            .I(N__12417));
    LocalMux I__2130 (
            .O(N__12417),
            .I(N__12414));
    Span4Mux_h I__2129 (
            .O(N__12414),
            .I(N__12411));
    Odrv4 I__2128 (
            .O(N__12411),
            .I(\Lab_UT.didp.countrce1.q_5_0 ));
    InMux I__2127 (
            .O(N__12408),
            .I(N__12405));
    LocalMux I__2126 (
            .O(N__12405),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ));
    InMux I__2125 (
            .O(N__12402),
            .I(N__12398));
    InMux I__2124 (
            .O(N__12401),
            .I(N__12394));
    LocalMux I__2123 (
            .O(N__12398),
            .I(N__12391));
    InMux I__2122 (
            .O(N__12397),
            .I(N__12388));
    LocalMux I__2121 (
            .O(N__12394),
            .I(N__12385));
    Span4Mux_v I__2120 (
            .O(N__12391),
            .I(N__12382));
    LocalMux I__2119 (
            .O(N__12388),
            .I(N__12379));
    Odrv4 I__2118 (
            .O(N__12385),
            .I(\Lab_UT.di_AStens_0 ));
    Odrv4 I__2117 (
            .O(N__12382),
            .I(\Lab_UT.di_AStens_0 ));
    Odrv12 I__2116 (
            .O(N__12379),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__2115 (
            .O(N__12372),
            .I(N__12369));
    LocalMux I__2114 (
            .O(N__12369),
            .I(N__12366));
    Span4Mux_h I__2113 (
            .O(N__12366),
            .I(N__12361));
    InMux I__2112 (
            .O(N__12365),
            .I(N__12356));
    InMux I__2111 (
            .O(N__12364),
            .I(N__12356));
    Span4Mux_v I__2110 (
            .O(N__12361),
            .I(N__12353));
    LocalMux I__2109 (
            .O(N__12356),
            .I(N__12350));
    Odrv4 I__2108 (
            .O(N__12353),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv12 I__2107 (
            .O(N__12350),
            .I(\Lab_UT.di_AStens_3 ));
    CascadeMux I__2106 (
            .O(N__12345),
            .I(N__12342));
    InMux I__2105 (
            .O(N__12342),
            .I(N__12339));
    LocalMux I__2104 (
            .O(N__12339),
            .I(\Lab_UT.didp.countrce2.N_93 ));
    InMux I__2103 (
            .O(N__12336),
            .I(N__12333));
    LocalMux I__2102 (
            .O(N__12333),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ));
    CascadeMux I__2101 (
            .O(N__12330),
            .I(\Lab_UT.didp.countrce2.N_96_cascade_ ));
    InMux I__2100 (
            .O(N__12327),
            .I(N__12324));
    LocalMux I__2099 (
            .O(N__12324),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_3 ));
    CascadeMux I__2098 (
            .O(N__12321),
            .I(N__12318));
    InMux I__2097 (
            .O(N__12318),
            .I(N__12315));
    LocalMux I__2096 (
            .O(N__12315),
            .I(N__12312));
    Odrv4 I__2095 (
            .O(N__12312),
            .I(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_1 ));
    CascadeMux I__2094 (
            .O(N__12309),
            .I(N__12302));
    InMux I__2093 (
            .O(N__12308),
            .I(N__12299));
    InMux I__2092 (
            .O(N__12307),
            .I(N__12296));
    InMux I__2091 (
            .O(N__12306),
            .I(N__12293));
    InMux I__2090 (
            .O(N__12305),
            .I(N__12288));
    InMux I__2089 (
            .O(N__12302),
            .I(N__12288));
    LocalMux I__2088 (
            .O(N__12299),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2087 (
            .O(N__12296),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2086 (
            .O(N__12293),
            .I(\Lab_UT.di_Stens_3 ));
    LocalMux I__2085 (
            .O(N__12288),
            .I(\Lab_UT.di_Stens_3 ));
    CascadeMux I__2084 (
            .O(N__12279),
            .I(N__12276));
    InMux I__2083 (
            .O(N__12276),
            .I(N__12268));
    InMux I__2082 (
            .O(N__12275),
            .I(N__12268));
    InMux I__2081 (
            .O(N__12274),
            .I(N__12263));
    InMux I__2080 (
            .O(N__12273),
            .I(N__12263));
    LocalMux I__2079 (
            .O(N__12268),
            .I(N__12259));
    LocalMux I__2078 (
            .O(N__12263),
            .I(N__12256));
    InMux I__2077 (
            .O(N__12262),
            .I(N__12253));
    Span4Mux_h I__2076 (
            .O(N__12259),
            .I(N__12250));
    Odrv4 I__2075 (
            .O(N__12256),
            .I(\Lab_UT.didp.un24_ce_3 ));
    LocalMux I__2074 (
            .O(N__12253),
            .I(\Lab_UT.didp.un24_ce_3 ));
    Odrv4 I__2073 (
            .O(N__12250),
            .I(\Lab_UT.didp.un24_ce_3 ));
    InMux I__2072 (
            .O(N__12243),
            .I(N__12240));
    LocalMux I__2071 (
            .O(N__12240),
            .I(N__12237));
    Span4Mux_h I__2070 (
            .O(N__12237),
            .I(N__12234));
    Odrv4 I__2069 (
            .O(N__12234),
            .I(\uu2.bitmapZ0Z_180 ));
    InMux I__2068 (
            .O(N__12231),
            .I(N__12228));
    LocalMux I__2067 (
            .O(N__12228),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__2066 (
            .O(N__12225),
            .I(N__12222));
    LocalMux I__2065 (
            .O(N__12222),
            .I(\uu2.bitmapZ0Z_52 ));
    InMux I__2064 (
            .O(N__12219),
            .I(N__12216));
    LocalMux I__2063 (
            .O(N__12216),
            .I(N__12213));
    Span4Mux_h I__2062 (
            .O(N__12213),
            .I(N__12210));
    Odrv4 I__2061 (
            .O(N__12210),
            .I(\uu2.N_149 ));
    InMux I__2060 (
            .O(N__12207),
            .I(N__12204));
    LocalMux I__2059 (
            .O(N__12204),
            .I(\uu2.bitmapZ0Z_84 ));
    CascadeMux I__2058 (
            .O(N__12201),
            .I(N__12198));
    InMux I__2057 (
            .O(N__12198),
            .I(N__12195));
    LocalMux I__2056 (
            .O(N__12195),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__2055 (
            .O(N__12192),
            .I(N__12189));
    LocalMux I__2054 (
            .O(N__12189),
            .I(\uu2.N_25 ));
    InMux I__2053 (
            .O(N__12186),
            .I(N__12177));
    InMux I__2052 (
            .O(N__12185),
            .I(N__12177));
    InMux I__2051 (
            .O(N__12184),
            .I(N__12177));
    LocalMux I__2050 (
            .O(N__12177),
            .I(\Lab_UT.didp.countrce1.ce_12_1_1 ));
    InMux I__2049 (
            .O(N__12174),
            .I(N__12170));
    InMux I__2048 (
            .O(N__12173),
            .I(N__12166));
    LocalMux I__2047 (
            .O(N__12170),
            .I(N__12163));
    InMux I__2046 (
            .O(N__12169),
            .I(N__12160));
    LocalMux I__2045 (
            .O(N__12166),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__2044 (
            .O(N__12163),
            .I(\Lab_UT.di_AMones_2 ));
    LocalMux I__2043 (
            .O(N__12160),
            .I(\Lab_UT.di_AMones_2 ));
    CascadeMux I__2042 (
            .O(N__12153),
            .I(N__12150));
    InMux I__2041 (
            .O(N__12150),
            .I(N__12147));
    LocalMux I__2040 (
            .O(N__12147),
            .I(N__12144));
    Span4Mux_v I__2039 (
            .O(N__12144),
            .I(N__12141));
    Odrv4 I__2038 (
            .O(N__12141),
            .I(\Lab_UT.didp.countrce4.un20_qPone ));
    InMux I__2037 (
            .O(N__12138),
            .I(N__12132));
    InMux I__2036 (
            .O(N__12137),
            .I(N__12132));
    LocalMux I__2035 (
            .O(N__12132),
            .I(N__12128));
    InMux I__2034 (
            .O(N__12131),
            .I(N__12124));
    Span4Mux_s2_v I__2033 (
            .O(N__12128),
            .I(N__12121));
    InMux I__2032 (
            .O(N__12127),
            .I(N__12118));
    LocalMux I__2031 (
            .O(N__12124),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    Odrv4 I__2030 (
            .O(N__12121),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    LocalMux I__2029 (
            .O(N__12118),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__2028 (
            .O(N__12111),
            .I(N__12108));
    LocalMux I__2027 (
            .O(N__12108),
            .I(N__12103));
    InMux I__2026 (
            .O(N__12107),
            .I(N__12100));
    InMux I__2025 (
            .O(N__12106),
            .I(N__12096));
    Span4Mux_v I__2024 (
            .O(N__12103),
            .I(N__12088));
    LocalMux I__2023 (
            .O(N__12100),
            .I(N__12085));
    CascadeMux I__2022 (
            .O(N__12099),
            .I(N__12081));
    LocalMux I__2021 (
            .O(N__12096),
            .I(N__12076));
    CascadeMux I__2020 (
            .O(N__12095),
            .I(N__12073));
    CascadeMux I__2019 (
            .O(N__12094),
            .I(N__12069));
    CascadeMux I__2018 (
            .O(N__12093),
            .I(N__12066));
    CascadeMux I__2017 (
            .O(N__12092),
            .I(N__12063));
    CascadeMux I__2016 (
            .O(N__12091),
            .I(N__12060));
    Span4Mux_h I__2015 (
            .O(N__12088),
            .I(N__12057));
    Span4Mux_s2_v I__2014 (
            .O(N__12085),
            .I(N__12054));
    InMux I__2013 (
            .O(N__12084),
            .I(N__12045));
    InMux I__2012 (
            .O(N__12081),
            .I(N__12045));
    InMux I__2011 (
            .O(N__12080),
            .I(N__12045));
    InMux I__2010 (
            .O(N__12079),
            .I(N__12045));
    Span4Mux_s2_v I__2009 (
            .O(N__12076),
            .I(N__12042));
    InMux I__2008 (
            .O(N__12073),
            .I(N__12033));
    InMux I__2007 (
            .O(N__12072),
            .I(N__12033));
    InMux I__2006 (
            .O(N__12069),
            .I(N__12033));
    InMux I__2005 (
            .O(N__12066),
            .I(N__12033));
    InMux I__2004 (
            .O(N__12063),
            .I(N__12028));
    InMux I__2003 (
            .O(N__12060),
            .I(N__12028));
    Odrv4 I__2002 (
            .O(N__12057),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2001 (
            .O(N__12054),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2000 (
            .O(N__12045),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__1999 (
            .O(N__12042),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__1998 (
            .O(N__12033),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__1997 (
            .O(N__12028),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__1996 (
            .O(N__12015),
            .I(N__12012));
    LocalMux I__1995 (
            .O(N__12012),
            .I(\uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ));
    CascadeMux I__1994 (
            .O(N__12009),
            .I(N__12006));
    InMux I__1993 (
            .O(N__12006),
            .I(N__12000));
    InMux I__1992 (
            .O(N__12005),
            .I(N__12000));
    LocalMux I__1991 (
            .O(N__12000),
            .I(N__11997));
    Span4Mux_s2_v I__1990 (
            .O(N__11997),
            .I(N__11994));
    Odrv4 I__1989 (
            .O(N__11994),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    InMux I__1988 (
            .O(N__11991),
            .I(N__11988));
    LocalMux I__1987 (
            .O(N__11988),
            .I(\uu2.bitmapZ0Z_75 ));
    CascadeMux I__1986 (
            .O(N__11985),
            .I(N__11982));
    InMux I__1985 (
            .O(N__11982),
            .I(N__11979));
    LocalMux I__1984 (
            .O(N__11979),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__1983 (
            .O(N__11976),
            .I(N__11973));
    LocalMux I__1982 (
            .O(N__11973),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__1981 (
            .O(N__11970),
            .I(N__11967));
    LocalMux I__1980 (
            .O(N__11967),
            .I(N__11964));
    Odrv4 I__1979 (
            .O(N__11964),
            .I(\uu2.w_addr_displaying_fastZ0Z_1 ));
    CascadeMux I__1978 (
            .O(N__11961),
            .I(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ));
    InMux I__1977 (
            .O(N__11958),
            .I(N__11955));
    LocalMux I__1976 (
            .O(N__11955),
            .I(\uu2.N_14 ));
    InMux I__1975 (
            .O(N__11952),
            .I(N__11949));
    LocalMux I__1974 (
            .O(N__11949),
            .I(N__11946));
    Odrv4 I__1973 (
            .O(N__11946),
            .I(\uu2.bitmap_RNI2Q8F1Z0Z_111 ));
    InMux I__1972 (
            .O(N__11943),
            .I(N__11940));
    LocalMux I__1971 (
            .O(N__11940),
            .I(\uu2.bitmapZ0Z_40 ));
    InMux I__1970 (
            .O(N__11937),
            .I(N__11930));
    InMux I__1969 (
            .O(N__11936),
            .I(N__11927));
    InMux I__1968 (
            .O(N__11935),
            .I(N__11920));
    InMux I__1967 (
            .O(N__11934),
            .I(N__11920));
    InMux I__1966 (
            .O(N__11933),
            .I(N__11920));
    LocalMux I__1965 (
            .O(N__11930),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__1964 (
            .O(N__11927),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__1963 (
            .O(N__11920),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__1962 (
            .O(N__11913),
            .I(N__11910));
    LocalMux I__1961 (
            .O(N__11910),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__1960 (
            .O(N__11907),
            .I(N__11904));
    LocalMux I__1959 (
            .O(N__11904),
            .I(\uu2.N_166 ));
    CEMux I__1958 (
            .O(N__11901),
            .I(N__11898));
    LocalMux I__1957 (
            .O(N__11898),
            .I(N__11894));
    CEMux I__1956 (
            .O(N__11897),
            .I(N__11891));
    Span4Mux_h I__1955 (
            .O(N__11894),
            .I(N__11887));
    LocalMux I__1954 (
            .O(N__11891),
            .I(N__11884));
    CEMux I__1953 (
            .O(N__11890),
            .I(N__11881));
    Span4Mux_h I__1952 (
            .O(N__11887),
            .I(N__11878));
    Span4Mux_s0_v I__1951 (
            .O(N__11884),
            .I(N__11875));
    LocalMux I__1950 (
            .O(N__11881),
            .I(N__11872));
    Odrv4 I__1949 (
            .O(N__11878),
            .I(\uu2.N_33_1 ));
    Odrv4 I__1948 (
            .O(N__11875),
            .I(\uu2.N_33_1 ));
    Odrv12 I__1947 (
            .O(N__11872),
            .I(\uu2.N_33_1 ));
    CascadeMux I__1946 (
            .O(N__11865),
            .I(N__11862));
    InMux I__1945 (
            .O(N__11862),
            .I(N__11859));
    LocalMux I__1944 (
            .O(N__11859),
            .I(N__11856));
    Span4Mux_s0_v I__1943 (
            .O(N__11856),
            .I(N__11853));
    Odrv4 I__1942 (
            .O(N__11853),
            .I(\uu2.mem0.w_addr_6 ));
    CascadeMux I__1941 (
            .O(N__11850),
            .I(N__11847));
    InMux I__1940 (
            .O(N__11847),
            .I(N__11844));
    LocalMux I__1939 (
            .O(N__11844),
            .I(N__11841));
    Odrv12 I__1938 (
            .O(N__11841),
            .I(\uu2.mem0.w_addr_4 ));
    CascadeMux I__1937 (
            .O(N__11838),
            .I(N__11835));
    InMux I__1936 (
            .O(N__11835),
            .I(N__11832));
    LocalMux I__1935 (
            .O(N__11832),
            .I(N__11829));
    Odrv12 I__1934 (
            .O(N__11829),
            .I(\uu2.mem0.w_addr_5 ));
    CascadeMux I__1933 (
            .O(N__11826),
            .I(N__11823));
    InMux I__1932 (
            .O(N__11823),
            .I(N__11820));
    LocalMux I__1931 (
            .O(N__11820),
            .I(N__11817));
    Odrv12 I__1930 (
            .O(N__11817),
            .I(\uu2.mem0.w_addr_7 ));
    InMux I__1929 (
            .O(N__11814),
            .I(N__11811));
    LocalMux I__1928 (
            .O(N__11811),
            .I(\Lab_UT.dictrl.g1_0Z0Z_5 ));
    CascadeMux I__1927 (
            .O(N__11808),
            .I(\Lab_UT.dictrl.g1_0_4_0_cascade_ ));
    InMux I__1926 (
            .O(N__11805),
            .I(N__11802));
    LocalMux I__1925 (
            .O(N__11802),
            .I(\Lab_UT.dictrl.g0_5_4_0 ));
    CascadeMux I__1924 (
            .O(N__11799),
            .I(\Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ));
    CascadeMux I__1923 (
            .O(N__11796),
            .I(\Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ));
    InMux I__1922 (
            .O(N__11793),
            .I(N__11790));
    LocalMux I__1921 (
            .O(N__11790),
            .I(\Lab_UT.dictrl.g0_5_3_0 ));
    CascadeMux I__1920 (
            .O(N__11787),
            .I(\Lab_UT.dictrl.G_25_i_o3_3_cascade_ ));
    InMux I__1919 (
            .O(N__11784),
            .I(N__11781));
    LocalMux I__1918 (
            .O(N__11781),
            .I(\Lab_UT.dictrl.alarmstate8Z0Z_3 ));
    CEMux I__1917 (
            .O(N__11778),
            .I(N__11775));
    LocalMux I__1916 (
            .O(N__11775),
            .I(N__11772));
    Odrv4 I__1915 (
            .O(N__11772),
            .I(\Lab_UT.didp.regrce2.LdAStens_0 ));
    CascadeMux I__1914 (
            .O(N__11769),
            .I(N__11765));
    CascadeMux I__1913 (
            .O(N__11768),
            .I(N__11762));
    InMux I__1912 (
            .O(N__11765),
            .I(N__11757));
    InMux I__1911 (
            .O(N__11762),
            .I(N__11757));
    LocalMux I__1910 (
            .O(N__11757),
            .I(N__11754));
    Span4Mux_v I__1909 (
            .O(N__11754),
            .I(N__11750));
    InMux I__1908 (
            .O(N__11753),
            .I(N__11747));
    Odrv4 I__1907 (
            .O(N__11750),
            .I(\Lab_UT.dictrl.alarmstateZ0Z8 ));
    LocalMux I__1906 (
            .O(N__11747),
            .I(\Lab_UT.dictrl.alarmstateZ0Z8 ));
    CascadeMux I__1905 (
            .O(N__11742),
            .I(N__11739));
    InMux I__1904 (
            .O(N__11739),
            .I(N__11736));
    LocalMux I__1903 (
            .O(N__11736),
            .I(N__11733));
    Odrv4 I__1902 (
            .O(N__11733),
            .I(\Lab_UT.dictrl.m37_N_2LZ0Z1 ));
    CascadeMux I__1901 (
            .O(N__11730),
            .I(\Lab_UT.didp.countrce4.q_5_3_cascade_ ));
    InMux I__1900 (
            .O(N__11727),
            .I(N__11724));
    LocalMux I__1899 (
            .O(N__11724),
            .I(N__11721));
    Odrv4 I__1898 (
            .O(N__11721),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_2 ));
    InMux I__1897 (
            .O(N__11718),
            .I(N__11715));
    LocalMux I__1896 (
            .O(N__11715),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_2_2 ));
    CascadeMux I__1895 (
            .O(N__11712),
            .I(\Lab_UT.didp.countrce4.q_5_0_cascade_ ));
    CascadeMux I__1894 (
            .O(N__11709),
            .I(N__11705));
    CascadeMux I__1893 (
            .O(N__11708),
            .I(N__11694));
    InMux I__1892 (
            .O(N__11705),
            .I(N__11690));
    InMux I__1891 (
            .O(N__11704),
            .I(N__11685));
    InMux I__1890 (
            .O(N__11703),
            .I(N__11685));
    InMux I__1889 (
            .O(N__11702),
            .I(N__11680));
    InMux I__1888 (
            .O(N__11701),
            .I(N__11680));
    InMux I__1887 (
            .O(N__11700),
            .I(N__11671));
    InMux I__1886 (
            .O(N__11699),
            .I(N__11671));
    InMux I__1885 (
            .O(N__11698),
            .I(N__11671));
    InMux I__1884 (
            .O(N__11697),
            .I(N__11671));
    InMux I__1883 (
            .O(N__11694),
            .I(N__11666));
    InMux I__1882 (
            .O(N__11693),
            .I(N__11666));
    LocalMux I__1881 (
            .O(N__11690),
            .I(G_181));
    LocalMux I__1880 (
            .O(N__11685),
            .I(G_181));
    LocalMux I__1879 (
            .O(N__11680),
            .I(G_181));
    LocalMux I__1878 (
            .O(N__11671),
            .I(G_181));
    LocalMux I__1877 (
            .O(N__11666),
            .I(G_181));
    InMux I__1876 (
            .O(N__11655),
            .I(N__11638));
    InMux I__1875 (
            .O(N__11654),
            .I(N__11638));
    InMux I__1874 (
            .O(N__11653),
            .I(N__11638));
    InMux I__1873 (
            .O(N__11652),
            .I(N__11633));
    InMux I__1872 (
            .O(N__11651),
            .I(N__11633));
    InMux I__1871 (
            .O(N__11650),
            .I(N__11630));
    InMux I__1870 (
            .O(N__11649),
            .I(N__11625));
    InMux I__1869 (
            .O(N__11648),
            .I(N__11625));
    InMux I__1868 (
            .O(N__11647),
            .I(N__11622));
    InMux I__1867 (
            .O(N__11646),
            .I(N__11619));
    InMux I__1866 (
            .O(N__11645),
            .I(N__11616));
    LocalMux I__1865 (
            .O(N__11638),
            .I(G_179));
    LocalMux I__1864 (
            .O(N__11633),
            .I(G_179));
    LocalMux I__1863 (
            .O(N__11630),
            .I(G_179));
    LocalMux I__1862 (
            .O(N__11625),
            .I(G_179));
    LocalMux I__1861 (
            .O(N__11622),
            .I(G_179));
    LocalMux I__1860 (
            .O(N__11619),
            .I(G_179));
    LocalMux I__1859 (
            .O(N__11616),
            .I(G_179));
    CascadeMux I__1858 (
            .O(N__11601),
            .I(N__11598));
    InMux I__1857 (
            .O(N__11598),
            .I(N__11595));
    LocalMux I__1856 (
            .O(N__11595),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0 ));
    CascadeMux I__1855 (
            .O(N__11592),
            .I(N__11588));
    CascadeMux I__1854 (
            .O(N__11591),
            .I(N__11584));
    InMux I__1853 (
            .O(N__11588),
            .I(N__11574));
    InMux I__1852 (
            .O(N__11587),
            .I(N__11574));
    InMux I__1851 (
            .O(N__11584),
            .I(N__11574));
    InMux I__1850 (
            .O(N__11583),
            .I(N__11571));
    InMux I__1849 (
            .O(N__11582),
            .I(N__11568));
    InMux I__1848 (
            .O(N__11581),
            .I(N__11565));
    LocalMux I__1847 (
            .O(N__11574),
            .I(N__11562));
    LocalMux I__1846 (
            .O(N__11571),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    LocalMux I__1845 (
            .O(N__11568),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    LocalMux I__1844 (
            .O(N__11565),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    Odrv4 I__1843 (
            .O(N__11562),
            .I(\Lab_UT.dispString.un42_dOutP_1 ));
    CascadeMux I__1842 (
            .O(N__11553),
            .I(N__11548));
    InMux I__1841 (
            .O(N__11552),
            .I(N__11545));
    InMux I__1840 (
            .O(N__11551),
            .I(N__11541));
    InMux I__1839 (
            .O(N__11548),
            .I(N__11538));
    LocalMux I__1838 (
            .O(N__11545),
            .I(N__11535));
    InMux I__1837 (
            .O(N__11544),
            .I(N__11532));
    LocalMux I__1836 (
            .O(N__11541),
            .I(\Lab_UT.dispString.N_95 ));
    LocalMux I__1835 (
            .O(N__11538),
            .I(\Lab_UT.dispString.N_95 ));
    Odrv4 I__1834 (
            .O(N__11535),
            .I(\Lab_UT.dispString.N_95 ));
    LocalMux I__1833 (
            .O(N__11532),
            .I(\Lab_UT.dispString.N_95 ));
    CascadeMux I__1832 (
            .O(N__11523),
            .I(N__11520));
    InMux I__1831 (
            .O(N__11520),
            .I(N__11517));
    LocalMux I__1830 (
            .O(N__11517),
            .I(\Lab_UT.dispString.N_140 ));
    CascadeMux I__1829 (
            .O(N__11514),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_ ));
    InMux I__1828 (
            .O(N__11511),
            .I(N__11508));
    LocalMux I__1827 (
            .O(N__11508),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2 ));
    InMux I__1826 (
            .O(N__11505),
            .I(N__11502));
    LocalMux I__1825 (
            .O(N__11502),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ));
    CascadeMux I__1824 (
            .O(N__11499),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ));
    InMux I__1823 (
            .O(N__11496),
            .I(N__11490));
    InMux I__1822 (
            .O(N__11495),
            .I(N__11483));
    InMux I__1821 (
            .O(N__11494),
            .I(N__11483));
    InMux I__1820 (
            .O(N__11493),
            .I(N__11483));
    LocalMux I__1819 (
            .O(N__11490),
            .I(N__11478));
    LocalMux I__1818 (
            .O(N__11483),
            .I(N__11478));
    Span4Mux_h I__1817 (
            .O(N__11478),
            .I(N__11475));
    Odrv4 I__1816 (
            .O(N__11475),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ));
    CascadeMux I__1815 (
            .O(N__11472),
            .I(N__11469));
    InMux I__1814 (
            .O(N__11469),
            .I(N__11466));
    LocalMux I__1813 (
            .O(N__11466),
            .I(\Lab_UT.didp.countrce1.un20_qPone ));
    CascadeMux I__1812 (
            .O(N__11463),
            .I(\Lab_UT.didp.countrce1.q_5_3_cascade_ ));
    InMux I__1811 (
            .O(N__11460),
            .I(N__11457));
    LocalMux I__1810 (
            .O(N__11457),
            .I(N__11454));
    Span4Mux_h I__1809 (
            .O(N__11454),
            .I(N__11451));
    Odrv4 I__1808 (
            .O(N__11451),
            .I(\Lab_UT.dispString.N_137 ));
    InMux I__1807 (
            .O(N__11448),
            .I(N__11445));
    LocalMux I__1806 (
            .O(N__11445),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ));
    InMux I__1805 (
            .O(N__11442),
            .I(N__11439));
    LocalMux I__1804 (
            .O(N__11439),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ));
    InMux I__1803 (
            .O(N__11436),
            .I(N__11430));
    InMux I__1802 (
            .O(N__11435),
            .I(N__11430));
    LocalMux I__1801 (
            .O(N__11430),
            .I(N__11425));
    InMux I__1800 (
            .O(N__11429),
            .I(N__11420));
    InMux I__1799 (
            .O(N__11428),
            .I(N__11420));
    Odrv4 I__1798 (
            .O(N__11425),
            .I(\Lab_UT.didp.ce_12_1 ));
    LocalMux I__1797 (
            .O(N__11420),
            .I(\Lab_UT.didp.ce_12_1 ));
    CascadeMux I__1796 (
            .O(N__11415),
            .I(\Lab_UT.didp.ce_12_1_cascade_ ));
    CascadeMux I__1795 (
            .O(N__11412),
            .I(\Lab_UT.didp.ce_12_3_cascade_ ));
    InMux I__1794 (
            .O(N__11409),
            .I(N__11406));
    LocalMux I__1793 (
            .O(N__11406),
            .I(N__11403));
    Span4Mux_h I__1792 (
            .O(N__11403),
            .I(N__11400));
    Odrv4 I__1791 (
            .O(N__11400),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_1 ));
    CascadeMux I__1790 (
            .O(N__11397),
            .I(N__11389));
    InMux I__1789 (
            .O(N__11396),
            .I(N__11385));
    InMux I__1788 (
            .O(N__11395),
            .I(N__11382));
    InMux I__1787 (
            .O(N__11394),
            .I(N__11371));
    InMux I__1786 (
            .O(N__11393),
            .I(N__11371));
    InMux I__1785 (
            .O(N__11392),
            .I(N__11371));
    InMux I__1784 (
            .O(N__11389),
            .I(N__11371));
    InMux I__1783 (
            .O(N__11388),
            .I(N__11371));
    LocalMux I__1782 (
            .O(N__11385),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__1781 (
            .O(N__11382),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    LocalMux I__1780 (
            .O(N__11371),
            .I(\uu2.w_addr_displaying_1_repZ0Z1 ));
    CascadeMux I__1779 (
            .O(N__11364),
            .I(\uu2.N_24_cascade_ ));
    InMux I__1778 (
            .O(N__11361),
            .I(N__11358));
    LocalMux I__1777 (
            .O(N__11358),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__1776 (
            .O(N__11355),
            .I(N__11352));
    InMux I__1775 (
            .O(N__11352),
            .I(N__11349));
    LocalMux I__1774 (
            .O(N__11349),
            .I(\uu2.bitmapZ0Z_221 ));
    InMux I__1773 (
            .O(N__11346),
            .I(N__11342));
    InMux I__1772 (
            .O(N__11345),
            .I(N__11339));
    LocalMux I__1771 (
            .O(N__11342),
            .I(\uu2.N_31_i ));
    LocalMux I__1770 (
            .O(N__11339),
            .I(\uu2.N_31_i ));
    CascadeMux I__1769 (
            .O(N__11334),
            .I(\uu2.N_26_cascade_ ));
    InMux I__1768 (
            .O(N__11331),
            .I(N__11328));
    LocalMux I__1767 (
            .O(N__11328),
            .I(\uu2.bitmap_pmux_27_ns_1 ));
    InMux I__1766 (
            .O(N__11325),
            .I(N__11322));
    LocalMux I__1765 (
            .O(N__11322),
            .I(\uu2.N_404 ));
    CascadeMux I__1764 (
            .O(N__11319),
            .I(N__11315));
    CascadeMux I__1763 (
            .O(N__11318),
            .I(N__11312));
    InMux I__1762 (
            .O(N__11315),
            .I(N__11306));
    InMux I__1761 (
            .O(N__11312),
            .I(N__11306));
    InMux I__1760 (
            .O(N__11311),
            .I(N__11303));
    LocalMux I__1759 (
            .O(N__11306),
            .I(N__11298));
    LocalMux I__1758 (
            .O(N__11303),
            .I(N__11298));
    Odrv4 I__1757 (
            .O(N__11298),
            .I(\uu2.un51_w_data_displaying_i_a2_1 ));
    CascadeMux I__1756 (
            .O(N__11295),
            .I(\uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ));
    InMux I__1755 (
            .O(N__11292),
            .I(N__11286));
    InMux I__1754 (
            .O(N__11291),
            .I(N__11286));
    LocalMux I__1753 (
            .O(N__11286),
            .I(N__11283));
    Odrv4 I__1752 (
            .O(N__11283),
            .I(\uu2.w_data_displaying_2_i_a2_i_a3_2_0 ));
    InMux I__1751 (
            .O(N__11280),
            .I(N__11276));
    InMux I__1750 (
            .O(N__11279),
            .I(N__11273));
    LocalMux I__1749 (
            .O(N__11276),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    LocalMux I__1748 (
            .O(N__11273),
            .I(\uu2.bitmap_pmux_sn_N_33 ));
    InMux I__1747 (
            .O(N__11268),
            .I(N__11265));
    LocalMux I__1746 (
            .O(N__11265),
            .I(N__11262));
    Odrv4 I__1745 (
            .O(N__11262),
            .I(\uu2.w_addr_displaying_RNI03P31Z0Z_4 ));
    CascadeMux I__1744 (
            .O(N__11259),
            .I(\uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ));
    InMux I__1743 (
            .O(N__11256),
            .I(N__11253));
    LocalMux I__1742 (
            .O(N__11253),
            .I(N__11250));
    Odrv4 I__1741 (
            .O(N__11250),
            .I(\uu2.bitmap_pmux_sn_i7_mux_0 ));
    InMux I__1740 (
            .O(N__11247),
            .I(N__11229));
    InMux I__1739 (
            .O(N__11246),
            .I(N__11229));
    InMux I__1738 (
            .O(N__11245),
            .I(N__11229));
    InMux I__1737 (
            .O(N__11244),
            .I(N__11229));
    InMux I__1736 (
            .O(N__11243),
            .I(N__11229));
    InMux I__1735 (
            .O(N__11242),
            .I(N__11229));
    LocalMux I__1734 (
            .O(N__11229),
            .I(\uu2.un28_w_addr_user_i ));
    InMux I__1733 (
            .O(N__11226),
            .I(N__11223));
    LocalMux I__1732 (
            .O(N__11223),
            .I(G_180));
    CascadeMux I__1731 (
            .O(N__11220),
            .I(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ));
    InMux I__1730 (
            .O(N__11217),
            .I(N__11210));
    InMux I__1729 (
            .O(N__11216),
            .I(N__11210));
    InMux I__1728 (
            .O(N__11215),
            .I(N__11207));
    LocalMux I__1727 (
            .O(N__11210),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    LocalMux I__1726 (
            .O(N__11207),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    CascadeMux I__1725 (
            .O(N__11202),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ));
    InMux I__1724 (
            .O(N__11199),
            .I(N__11195));
    InMux I__1723 (
            .O(N__11198),
            .I(N__11192));
    LocalMux I__1722 (
            .O(N__11195),
            .I(G_184));
    LocalMux I__1721 (
            .O(N__11192),
            .I(G_184));
    CascadeMux I__1720 (
            .O(N__11187),
            .I(\resetGen.escKeyZ0Z_5_cascade_ ));
    InMux I__1719 (
            .O(N__11184),
            .I(N__11178));
    InMux I__1718 (
            .O(N__11183),
            .I(N__11178));
    LocalMux I__1717 (
            .O(N__11178),
            .I(N__11172));
    InMux I__1716 (
            .O(N__11177),
            .I(N__11165));
    InMux I__1715 (
            .O(N__11176),
            .I(N__11165));
    InMux I__1714 (
            .O(N__11175),
            .I(N__11165));
    Span4Mux_v I__1713 (
            .O(N__11172),
            .I(N__11160));
    LocalMux I__1712 (
            .O(N__11165),
            .I(N__11160));
    Span4Mux_h I__1711 (
            .O(N__11160),
            .I(N__11157));
    Odrv4 I__1710 (
            .O(N__11157),
            .I(\resetGen.escKeyZ0 ));
    InMux I__1709 (
            .O(N__11154),
            .I(N__11151));
    LocalMux I__1708 (
            .O(N__11151),
            .I(\resetGen.escKeyZ0Z_4 ));
    InMux I__1707 (
            .O(N__11148),
            .I(N__11143));
    InMux I__1706 (
            .O(N__11147),
            .I(N__11140));
    InMux I__1705 (
            .O(N__11146),
            .I(N__11137));
    LocalMux I__1704 (
            .O(N__11143),
            .I(N__11134));
    LocalMux I__1703 (
            .O(N__11140),
            .I(G_186));
    LocalMux I__1702 (
            .O(N__11137),
            .I(G_186));
    Odrv4 I__1701 (
            .O(N__11134),
            .I(G_186));
    InMux I__1700 (
            .O(N__11127),
            .I(N__11124));
    LocalMux I__1699 (
            .O(N__11124),
            .I(N__11120));
    CascadeMux I__1698 (
            .O(N__11123),
            .I(N__11117));
    Span4Mux_v I__1697 (
            .O(N__11120),
            .I(N__11113));
    InMux I__1696 (
            .O(N__11117),
            .I(N__11110));
    InMux I__1695 (
            .O(N__11116),
            .I(N__11107));
    Odrv4 I__1694 (
            .O(N__11113),
            .I(L3_tx_data_6));
    LocalMux I__1693 (
            .O(N__11110),
            .I(L3_tx_data_6));
    LocalMux I__1692 (
            .O(N__11107),
            .I(L3_tx_data_6));
    SRMux I__1691 (
            .O(N__11100),
            .I(N__11097));
    LocalMux I__1690 (
            .O(N__11097),
            .I(N__11091));
    CascadeMux I__1689 (
            .O(N__11096),
            .I(N__11088));
    IoInMux I__1688 (
            .O(N__11095),
            .I(N__11085));
    InMux I__1687 (
            .O(N__11094),
            .I(N__11082));
    Span4Mux_s3_h I__1686 (
            .O(N__11091),
            .I(N__11079));
    InMux I__1685 (
            .O(N__11088),
            .I(N__11076));
    LocalMux I__1684 (
            .O(N__11085),
            .I(N__11073));
    LocalMux I__1683 (
            .O(N__11082),
            .I(N__11070));
    Span4Mux_v I__1682 (
            .O(N__11079),
            .I(N__11065));
    LocalMux I__1681 (
            .O(N__11076),
            .I(N__11065));
    Span12Mux_s5_v I__1680 (
            .O(N__11073),
            .I(N__11062));
    Span4Mux_v I__1679 (
            .O(N__11070),
            .I(N__11059));
    Span4Mux_v I__1678 (
            .O(N__11065),
            .I(N__11056));
    Odrv12 I__1677 (
            .O(N__11062),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1676 (
            .O(N__11059),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1675 (
            .O(N__11056),
            .I(CONSTANT_ONE_NET));
    InMux I__1674 (
            .O(N__11049),
            .I(N__11045));
    InMux I__1673 (
            .O(N__11048),
            .I(N__11042));
    LocalMux I__1672 (
            .O(N__11045),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0 ));
    LocalMux I__1671 (
            .O(N__11042),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0 ));
    CascadeMux I__1670 (
            .O(N__11037),
            .I(\Lab_UT.un1_idle_4_0_iclkZ0_cascade_ ));
    InMux I__1669 (
            .O(N__11034),
            .I(N__11031));
    LocalMux I__1668 (
            .O(N__11031),
            .I(G_185));
    CascadeMux I__1667 (
            .O(N__11028),
            .I(G_185_cascade_));
    CascadeMux I__1666 (
            .O(N__11025),
            .I(\Lab_UT.dispString.N_117_cascade_ ));
    InMux I__1665 (
            .O(N__11022),
            .I(N__11019));
    LocalMux I__1664 (
            .O(N__11019),
            .I(N__11016));
    Span4Mux_s1_v I__1663 (
            .O(N__11016),
            .I(N__11013));
    Span4Mux_v I__1662 (
            .O(N__11013),
            .I(N__11008));
    InMux I__1661 (
            .O(N__11012),
            .I(N__11003));
    InMux I__1660 (
            .O(N__11011),
            .I(N__11003));
    Odrv4 I__1659 (
            .O(N__11008),
            .I(L3_tx_data_1));
    LocalMux I__1658 (
            .O(N__11003),
            .I(L3_tx_data_1));
    InMux I__1657 (
            .O(N__10998),
            .I(N__10995));
    LocalMux I__1656 (
            .O(N__10995),
            .I(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ));
    CascadeMux I__1655 (
            .O(N__10992),
            .I(G_180_cascade_));
    CascadeMux I__1654 (
            .O(N__10989),
            .I(G_181_cascade_));
    CEMux I__1653 (
            .O(N__10986),
            .I(N__10983));
    LocalMux I__1652 (
            .O(N__10983),
            .I(N__10980));
    Span4Mux_v I__1651 (
            .O(N__10980),
            .I(N__10977));
    Odrv4 I__1650 (
            .O(N__10977),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    CascadeMux I__1649 (
            .O(N__10974),
            .I(N__10971));
    InMux I__1648 (
            .O(N__10971),
            .I(N__10968));
    LocalMux I__1647 (
            .O(N__10968),
            .I(\uu2.un1_w_user_lfZ0Z_4 ));
    InMux I__1646 (
            .O(N__10965),
            .I(N__10961));
    CascadeMux I__1645 (
            .O(N__10964),
            .I(N__10958));
    LocalMux I__1644 (
            .O(N__10961),
            .I(N__10954));
    InMux I__1643 (
            .O(N__10958),
            .I(N__10949));
    InMux I__1642 (
            .O(N__10957),
            .I(N__10949));
    Odrv12 I__1641 (
            .O(N__10954),
            .I(L3_tx_data_5));
    LocalMux I__1640 (
            .O(N__10949),
            .I(L3_tx_data_5));
    CascadeMux I__1639 (
            .O(N__10944),
            .I(N__10940));
    InMux I__1638 (
            .O(N__10943),
            .I(N__10936));
    InMux I__1637 (
            .O(N__10940),
            .I(N__10931));
    InMux I__1636 (
            .O(N__10939),
            .I(N__10931));
    LocalMux I__1635 (
            .O(N__10936),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    LocalMux I__1634 (
            .O(N__10931),
            .I(\uu2.un1_w_user_crZ0Z_4 ));
    InMux I__1633 (
            .O(N__10926),
            .I(N__10923));
    LocalMux I__1632 (
            .O(N__10923),
            .I(N__10920));
    Odrv12 I__1631 (
            .O(N__10920),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_3 ));
    InMux I__1630 (
            .O(N__10917),
            .I(N__10914));
    LocalMux I__1629 (
            .O(N__10914),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_1_3 ));
    InMux I__1628 (
            .O(N__10911),
            .I(N__10908));
    LocalMux I__1627 (
            .O(N__10908),
            .I(\uu2.un1_w_user_lfZ0Z_3 ));
    InMux I__1626 (
            .O(N__10905),
            .I(N__10902));
    LocalMux I__1625 (
            .O(N__10902),
            .I(N__10899));
    Span4Mux_s3_v I__1624 (
            .O(N__10899),
            .I(N__10894));
    InMux I__1623 (
            .O(N__10898),
            .I(N__10889));
    InMux I__1622 (
            .O(N__10897),
            .I(N__10889));
    Odrv4 I__1621 (
            .O(N__10894),
            .I(L3_tx_data_3));
    LocalMux I__1620 (
            .O(N__10889),
            .I(L3_tx_data_3));
    InMux I__1619 (
            .O(N__10884),
            .I(N__10881));
    LocalMux I__1618 (
            .O(N__10881),
            .I(N__10878));
    Span4Mux_s3_v I__1617 (
            .O(N__10878),
            .I(N__10873));
    InMux I__1616 (
            .O(N__10877),
            .I(N__10868));
    InMux I__1615 (
            .O(N__10876),
            .I(N__10868));
    Odrv4 I__1614 (
            .O(N__10873),
            .I(L3_tx_data_0));
    LocalMux I__1613 (
            .O(N__10868),
            .I(L3_tx_data_0));
    InMux I__1612 (
            .O(N__10863),
            .I(N__10858));
    InMux I__1611 (
            .O(N__10862),
            .I(N__10853));
    InMux I__1610 (
            .O(N__10861),
            .I(N__10853));
    LocalMux I__1609 (
            .O(N__10858),
            .I(\uu2.un1_w_user_crZ0Z_3 ));
    LocalMux I__1608 (
            .O(N__10853),
            .I(\uu2.un1_w_user_crZ0Z_3 ));
    InMux I__1607 (
            .O(N__10848),
            .I(N__10845));
    LocalMux I__1606 (
            .O(N__10845),
            .I(\Lab_UT.dispString.dOutP_1_iv_i_1_4 ));
    InMux I__1605 (
            .O(N__10842),
            .I(N__10839));
    LocalMux I__1604 (
            .O(N__10839),
            .I(N__10836));
    Span4Mux_v I__1603 (
            .O(N__10836),
            .I(N__10831));
    InMux I__1602 (
            .O(N__10835),
            .I(N__10826));
    InMux I__1601 (
            .O(N__10834),
            .I(N__10826));
    Odrv4 I__1600 (
            .O(N__10831),
            .I(L3_tx_data_4));
    LocalMux I__1599 (
            .O(N__10826),
            .I(L3_tx_data_4));
    InMux I__1598 (
            .O(N__10821),
            .I(N__10815));
    InMux I__1597 (
            .O(N__10820),
            .I(N__10815));
    LocalMux I__1596 (
            .O(N__10815),
            .I(\Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ));
    CascadeMux I__1595 (
            .O(N__10812),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ));
    InMux I__1594 (
            .O(N__10809),
            .I(N__10803));
    InMux I__1593 (
            .O(N__10808),
            .I(N__10803));
    LocalMux I__1592 (
            .O(N__10803),
            .I(N__10800));
    Odrv12 I__1591 (
            .O(N__10800),
            .I(\uu2.un20_w_addr_userZ0Z_1 ));
    InMux I__1590 (
            .O(N__10797),
            .I(N__10793));
    InMux I__1589 (
            .O(N__10796),
            .I(N__10789));
    LocalMux I__1588 (
            .O(N__10793),
            .I(N__10786));
    InMux I__1587 (
            .O(N__10792),
            .I(N__10783));
    LocalMux I__1586 (
            .O(N__10789),
            .I(L3_tx_data_rdy));
    Odrv12 I__1585 (
            .O(N__10786),
            .I(L3_tx_data_rdy));
    LocalMux I__1584 (
            .O(N__10783),
            .I(L3_tx_data_rdy));
    CascadeMux I__1583 (
            .O(N__10776),
            .I(\Lab_UT.dispString.N_124_cascade_ ));
    CascadeMux I__1582 (
            .O(N__10773),
            .I(\Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ));
    InMux I__1581 (
            .O(N__10770),
            .I(N__10767));
    LocalMux I__1580 (
            .O(N__10767),
            .I(\uu2.bitmap_pmux_sn_i5_mux ));
    InMux I__1579 (
            .O(N__10764),
            .I(N__10761));
    LocalMux I__1578 (
            .O(N__10761),
            .I(\uu2.bitmap_pmux_u_1 ));
    InMux I__1577 (
            .O(N__10758),
            .I(N__10754));
    InMux I__1576 (
            .O(N__10757),
            .I(N__10751));
    LocalMux I__1575 (
            .O(N__10754),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    LocalMux I__1574 (
            .O(N__10751),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    InMux I__1573 (
            .O(N__10746),
            .I(N__10743));
    LocalMux I__1572 (
            .O(N__10743),
            .I(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ));
    InMux I__1571 (
            .O(N__10740),
            .I(N__10737));
    LocalMux I__1570 (
            .O(N__10737),
            .I(\uu2.w_addr_displaying_RNI0NG56Z0Z_4 ));
    InMux I__1569 (
            .O(N__10734),
            .I(N__10730));
    InMux I__1568 (
            .O(N__10733),
            .I(N__10727));
    LocalMux I__1567 (
            .O(N__10730),
            .I(N__10724));
    LocalMux I__1566 (
            .O(N__10727),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__1565 (
            .O(N__10724),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__1564 (
            .O(N__10719),
            .I(N__10716));
    LocalMux I__1563 (
            .O(N__10716),
            .I(N__10713));
    Odrv12 I__1562 (
            .O(N__10713),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__1561 (
            .O(N__10710),
            .I(N__10707));
    LocalMux I__1560 (
            .O(N__10707),
            .I(\uu2.N_401 ));
    CascadeMux I__1559 (
            .O(N__10704),
            .I(\uu2.N_406_cascade_ ));
    InMux I__1558 (
            .O(N__10701),
            .I(N__10695));
    InMux I__1557 (
            .O(N__10700),
            .I(N__10695));
    LocalMux I__1556 (
            .O(N__10695),
            .I(\uu2.bitmap_pmux ));
    CascadeMux I__1555 (
            .O(N__10692),
            .I(\uu2.N_383_cascade_ ));
    CascadeMux I__1554 (
            .O(N__10689),
            .I(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ));
    InMux I__1553 (
            .O(N__10686),
            .I(N__10683));
    LocalMux I__1552 (
            .O(N__10683),
            .I(\uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ));
    CEMux I__1551 (
            .O(N__10680),
            .I(N__10677));
    LocalMux I__1550 (
            .O(N__10677),
            .I(N__10674));
    Odrv4 I__1549 (
            .O(N__10674),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    CascadeMux I__1548 (
            .O(N__10671),
            .I(\uu2.un28_w_addr_user_i_cascade_ ));
    CascadeMux I__1547 (
            .O(N__10668),
            .I(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ));
    CascadeMux I__1546 (
            .O(N__10665),
            .I(\uu2.bitmap_pmux_sn_N_15_cascade_ ));
    CascadeMux I__1545 (
            .O(N__10662),
            .I(G_182_cascade_));
    InMux I__1544 (
            .O(N__10659),
            .I(N__10654));
    InMux I__1543 (
            .O(N__10658),
            .I(N__10649));
    InMux I__1542 (
            .O(N__10657),
            .I(N__10649));
    LocalMux I__1541 (
            .O(N__10654),
            .I(G_187));
    LocalMux I__1540 (
            .O(N__10649),
            .I(G_187));
    CascadeMux I__1539 (
            .O(N__10644),
            .I(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ));
    InMux I__1538 (
            .O(N__10641),
            .I(N__10632));
    InMux I__1537 (
            .O(N__10640),
            .I(N__10632));
    InMux I__1536 (
            .O(N__10639),
            .I(N__10632));
    LocalMux I__1535 (
            .O(N__10632),
            .I(G_183));
    InMux I__1534 (
            .O(N__10629),
            .I(N__10623));
    InMux I__1533 (
            .O(N__10628),
            .I(N__10623));
    LocalMux I__1532 (
            .O(N__10623),
            .I(G_182));
    InMux I__1531 (
            .O(N__10620),
            .I(N__10611));
    InMux I__1530 (
            .O(N__10619),
            .I(N__10611));
    InMux I__1529 (
            .O(N__10618),
            .I(N__10606));
    InMux I__1528 (
            .O(N__10617),
            .I(N__10606));
    InMux I__1527 (
            .O(N__10616),
            .I(N__10603));
    LocalMux I__1526 (
            .O(N__10611),
            .I(N__10600));
    LocalMux I__1525 (
            .O(N__10606),
            .I(N__10596));
    LocalMux I__1524 (
            .O(N__10603),
            .I(N__10593));
    Span4Mux_s3_h I__1523 (
            .O(N__10600),
            .I(N__10590));
    InMux I__1522 (
            .O(N__10599),
            .I(N__10587));
    Span12Mux_s5_v I__1521 (
            .O(N__10596),
            .I(N__10582));
    Span12Mux_s3_h I__1520 (
            .O(N__10593),
            .I(N__10582));
    Span4Mux_v I__1519 (
            .O(N__10590),
            .I(N__10579));
    LocalMux I__1518 (
            .O(N__10587),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv12 I__1517 (
            .O(N__10582),
            .I(\uu2.l_countZ0Z_0 ));
    Odrv4 I__1516 (
            .O(N__10579),
            .I(\uu2.l_countZ0Z_0 ));
    InMux I__1515 (
            .O(N__10572),
            .I(N__10569));
    LocalMux I__1514 (
            .O(N__10569),
            .I(N__10566));
    Span4Mux_h I__1513 (
            .O(N__10566),
            .I(N__10563));
    Odrv4 I__1512 (
            .O(N__10563),
            .I(vbuf_tx_data_6));
    InMux I__1511 (
            .O(N__10560),
            .I(N__10557));
    LocalMux I__1510 (
            .O(N__10557),
            .I(N__10554));
    Span4Mux_h I__1509 (
            .O(N__10554),
            .I(N__10551));
    Odrv4 I__1508 (
            .O(N__10551),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    InMux I__1507 (
            .O(N__10548),
            .I(N__10545));
    LocalMux I__1506 (
            .O(N__10545),
            .I(N__10542));
    Odrv12 I__1505 (
            .O(N__10542),
            .I(vbuf_tx_data_7));
    InMux I__1504 (
            .O(N__10539),
            .I(N__10536));
    LocalMux I__1503 (
            .O(N__10536),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CascadeMux I__1502 (
            .O(N__10533),
            .I(N__10530));
    InMux I__1501 (
            .O(N__10530),
            .I(N__10527));
    LocalMux I__1500 (
            .O(N__10527),
            .I(N__10524));
    Odrv4 I__1499 (
            .O(N__10524),
            .I(\uu2.mem0.w_addr_8 ));
    SRMux I__1498 (
            .O(N__10521),
            .I(N__10518));
    LocalMux I__1497 (
            .O(N__10518),
            .I(N__10514));
    CEMux I__1496 (
            .O(N__10517),
            .I(N__10511));
    Span4Mux_s3_v I__1495 (
            .O(N__10514),
            .I(N__10508));
    LocalMux I__1494 (
            .O(N__10511),
            .I(N__10505));
    Span4Mux_h I__1493 (
            .O(N__10508),
            .I(N__10500));
    Span4Mux_s3_v I__1492 (
            .O(N__10505),
            .I(N__10500));
    Odrv4 I__1491 (
            .O(N__10500),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    InMux I__1490 (
            .O(N__10497),
            .I(N__10494));
    LocalMux I__1489 (
            .O(N__10494),
            .I(G_188));
    CascadeMux I__1488 (
            .O(N__10491),
            .I(G_188_cascade_));
    InMux I__1487 (
            .O(N__10488),
            .I(N__10485));
    LocalMux I__1486 (
            .O(N__10485),
            .I(\Lab_UT.un1_rst_0_iclkZ0 ));
    CascadeMux I__1485 (
            .O(N__10482),
            .I(N__10479));
    InMux I__1484 (
            .O(N__10479),
            .I(N__10473));
    InMux I__1483 (
            .O(N__10478),
            .I(N__10468));
    InMux I__1482 (
            .O(N__10477),
            .I(N__10468));
    CascadeMux I__1481 (
            .O(N__10476),
            .I(N__10465));
    LocalMux I__1480 (
            .O(N__10473),
            .I(N__10462));
    LocalMux I__1479 (
            .O(N__10468),
            .I(N__10459));
    InMux I__1478 (
            .O(N__10465),
            .I(N__10456));
    Span4Mux_s3_h I__1477 (
            .O(N__10462),
            .I(N__10451));
    Span4Mux_s1_v I__1476 (
            .O(N__10459),
            .I(N__10451));
    LocalMux I__1475 (
            .O(N__10456),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv4 I__1474 (
            .O(N__10451),
            .I(\uu2.r_addrZ0Z_5 ));
    InMux I__1473 (
            .O(N__10446),
            .I(N__10443));
    LocalMux I__1472 (
            .O(N__10443),
            .I(N__10436));
    InMux I__1471 (
            .O(N__10442),
            .I(N__10433));
    InMux I__1470 (
            .O(N__10441),
            .I(N__10426));
    InMux I__1469 (
            .O(N__10440),
            .I(N__10426));
    InMux I__1468 (
            .O(N__10439),
            .I(N__10426));
    Odrv4 I__1467 (
            .O(N__10436),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__1466 (
            .O(N__10433),
            .I(\uu2.l_countZ0Z_6 ));
    LocalMux I__1465 (
            .O(N__10426),
            .I(\uu2.l_countZ0Z_6 ));
    CascadeMux I__1464 (
            .O(N__10419),
            .I(N__10416));
    InMux I__1463 (
            .O(N__10416),
            .I(N__10412));
    CascadeMux I__1462 (
            .O(N__10415),
            .I(N__10409));
    LocalMux I__1461 (
            .O(N__10412),
            .I(N__10406));
    InMux I__1460 (
            .O(N__10409),
            .I(N__10403));
    Odrv4 I__1459 (
            .O(N__10406),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    LocalMux I__1458 (
            .O(N__10403),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    InMux I__1457 (
            .O(N__10398),
            .I(N__10395));
    LocalMux I__1456 (
            .O(N__10395),
            .I(N__10392));
    Span4Mux_h I__1455 (
            .O(N__10392),
            .I(N__10385));
    InMux I__1454 (
            .O(N__10391),
            .I(N__10376));
    InMux I__1453 (
            .O(N__10390),
            .I(N__10376));
    InMux I__1452 (
            .O(N__10389),
            .I(N__10376));
    InMux I__1451 (
            .O(N__10388),
            .I(N__10376));
    Odrv4 I__1450 (
            .O(N__10385),
            .I(\uu2.un306_ci ));
    LocalMux I__1449 (
            .O(N__10376),
            .I(\uu2.un306_ci ));
    InMux I__1448 (
            .O(N__10371),
            .I(N__10367));
    InMux I__1447 (
            .O(N__10370),
            .I(N__10364));
    LocalMux I__1446 (
            .O(N__10367),
            .I(N__10360));
    LocalMux I__1445 (
            .O(N__10364),
            .I(N__10357));
    InMux I__1444 (
            .O(N__10363),
            .I(N__10354));
    Span4Mux_s2_h I__1443 (
            .O(N__10360),
            .I(N__10349));
    Span4Mux_v I__1442 (
            .O(N__10357),
            .I(N__10349));
    LocalMux I__1441 (
            .O(N__10354),
            .I(\uu2.l_countZ0Z_7 ));
    Odrv4 I__1440 (
            .O(N__10349),
            .I(\uu2.l_countZ0Z_7 ));
    InMux I__1439 (
            .O(N__10344),
            .I(N__10338));
    InMux I__1438 (
            .O(N__10343),
            .I(N__10338));
    LocalMux I__1437 (
            .O(N__10338),
            .I(N__10335));
    Span4Mux_v I__1436 (
            .O(N__10335),
            .I(N__10332));
    Odrv4 I__1435 (
            .O(N__10332),
            .I(\uu2.un284_ci ));
    CascadeMux I__1434 (
            .O(N__10329),
            .I(N__10324));
    InMux I__1433 (
            .O(N__10328),
            .I(N__10320));
    InMux I__1432 (
            .O(N__10327),
            .I(N__10315));
    InMux I__1431 (
            .O(N__10324),
            .I(N__10315));
    CascadeMux I__1430 (
            .O(N__10323),
            .I(N__10312));
    LocalMux I__1429 (
            .O(N__10320),
            .I(N__10306));
    LocalMux I__1428 (
            .O(N__10315),
            .I(N__10306));
    InMux I__1427 (
            .O(N__10312),
            .I(N__10301));
    InMux I__1426 (
            .O(N__10311),
            .I(N__10301));
    Span4Mux_s3_h I__1425 (
            .O(N__10306),
            .I(N__10298));
    LocalMux I__1424 (
            .O(N__10301),
            .I(\uu2.l_countZ0Z_1 ));
    Odrv4 I__1423 (
            .O(N__10298),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__1422 (
            .O(N__10293),
            .I(N__10287));
    InMux I__1421 (
            .O(N__10292),
            .I(N__10287));
    LocalMux I__1420 (
            .O(N__10287),
            .I(\uu2.N_31 ));
    CascadeMux I__1419 (
            .O(N__10284),
            .I(\uu2.N_31_cascade_ ));
    InMux I__1418 (
            .O(N__10281),
            .I(N__10278));
    LocalMux I__1417 (
            .O(N__10278),
            .I(\uu2.mem0.w_data_0 ));
    CascadeMux I__1416 (
            .O(N__10275),
            .I(N__10270));
    InMux I__1415 (
            .O(N__10274),
            .I(N__10264));
    InMux I__1414 (
            .O(N__10273),
            .I(N__10264));
    InMux I__1413 (
            .O(N__10270),
            .I(N__10261));
    InMux I__1412 (
            .O(N__10269),
            .I(N__10258));
    LocalMux I__1411 (
            .O(N__10264),
            .I(N__10255));
    LocalMux I__1410 (
            .O(N__10261),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__1409 (
            .O(N__10258),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__1408 (
            .O(N__10255),
            .I(\uu2.r_addrZ0Z_2 ));
    CascadeMux I__1407 (
            .O(N__10248),
            .I(N__10244));
    CascadeMux I__1406 (
            .O(N__10247),
            .I(N__10239));
    InMux I__1405 (
            .O(N__10244),
            .I(N__10235));
    InMux I__1404 (
            .O(N__10243),
            .I(N__10230));
    InMux I__1403 (
            .O(N__10242),
            .I(N__10230));
    InMux I__1402 (
            .O(N__10239),
            .I(N__10225));
    InMux I__1401 (
            .O(N__10238),
            .I(N__10225));
    LocalMux I__1400 (
            .O(N__10235),
            .I(N__10220));
    LocalMux I__1399 (
            .O(N__10230),
            .I(N__10220));
    LocalMux I__1398 (
            .O(N__10225),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv4 I__1397 (
            .O(N__10220),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__1396 (
            .O(N__10215),
            .I(N__10210));
    InMux I__1395 (
            .O(N__10214),
            .I(N__10202));
    InMux I__1394 (
            .O(N__10213),
            .I(N__10202));
    InMux I__1393 (
            .O(N__10210),
            .I(N__10199));
    InMux I__1392 (
            .O(N__10209),
            .I(N__10192));
    InMux I__1391 (
            .O(N__10208),
            .I(N__10192));
    InMux I__1390 (
            .O(N__10207),
            .I(N__10192));
    LocalMux I__1389 (
            .O(N__10202),
            .I(N__10189));
    LocalMux I__1388 (
            .O(N__10199),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__1387 (
            .O(N__10192),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv4 I__1386 (
            .O(N__10189),
            .I(\uu2.r_addrZ0Z_0 ));
    CEMux I__1385 (
            .O(N__10182),
            .I(N__10179));
    LocalMux I__1384 (
            .O(N__10179),
            .I(N__10176));
    Span4Mux_s1_v I__1383 (
            .O(N__10176),
            .I(N__10173));
    Odrv4 I__1382 (
            .O(N__10173),
            .I(\uu2.trig_rd_is_det_0 ));
    InMux I__1381 (
            .O(N__10170),
            .I(N__10164));
    InMux I__1380 (
            .O(N__10169),
            .I(N__10161));
    InMux I__1379 (
            .O(N__10168),
            .I(N__10156));
    InMux I__1378 (
            .O(N__10167),
            .I(N__10156));
    LocalMux I__1377 (
            .O(N__10164),
            .I(N__10153));
    LocalMux I__1376 (
            .O(N__10161),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__1375 (
            .O(N__10156),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv4 I__1374 (
            .O(N__10153),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__1373 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__1372 (
            .O(N__10143),
            .I(N__10135));
    InMux I__1371 (
            .O(N__10142),
            .I(N__10124));
    InMux I__1370 (
            .O(N__10141),
            .I(N__10124));
    InMux I__1369 (
            .O(N__10140),
            .I(N__10124));
    InMux I__1368 (
            .O(N__10139),
            .I(N__10124));
    InMux I__1367 (
            .O(N__10138),
            .I(N__10124));
    Span4Mux_v I__1366 (
            .O(N__10135),
            .I(N__10119));
    LocalMux I__1365 (
            .O(N__10124),
            .I(N__10119));
    Odrv4 I__1364 (
            .O(N__10119),
            .I(\uu2.trig_rd_is_det ));
    CascadeMux I__1363 (
            .O(N__10116),
            .I(N__10110));
    InMux I__1362 (
            .O(N__10115),
            .I(N__10107));
    InMux I__1361 (
            .O(N__10114),
            .I(N__10101));
    InMux I__1360 (
            .O(N__10113),
            .I(N__10101));
    InMux I__1359 (
            .O(N__10110),
            .I(N__10098));
    LocalMux I__1358 (
            .O(N__10107),
            .I(N__10095));
    InMux I__1357 (
            .O(N__10106),
            .I(N__10092));
    LocalMux I__1356 (
            .O(N__10101),
            .I(N__10089));
    LocalMux I__1355 (
            .O(N__10098),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1354 (
            .O(N__10095),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__1353 (
            .O(N__10092),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__1352 (
            .O(N__10089),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__1351 (
            .O(N__10080),
            .I(N__10077));
    LocalMux I__1350 (
            .O(N__10077),
            .I(N__10073));
    InMux I__1349 (
            .O(N__10076),
            .I(N__10070));
    Span4Mux_v I__1348 (
            .O(N__10073),
            .I(N__10063));
    LocalMux I__1347 (
            .O(N__10070),
            .I(N__10063));
    InMux I__1346 (
            .O(N__10069),
            .I(N__10058));
    InMux I__1345 (
            .O(N__10068),
            .I(N__10058));
    Odrv4 I__1344 (
            .O(N__10063),
            .I(\uu2.un404_ci_0 ));
    LocalMux I__1343 (
            .O(N__10058),
            .I(\uu2.un404_ci_0 ));
    CascadeMux I__1342 (
            .O(N__10053),
            .I(\uu2.un404_ci_0_cascade_ ));
    CascadeMux I__1341 (
            .O(N__10050),
            .I(N__10047));
    InMux I__1340 (
            .O(N__10047),
            .I(N__10042));
    InMux I__1339 (
            .O(N__10046),
            .I(N__10039));
    InMux I__1338 (
            .O(N__10045),
            .I(N__10036));
    LocalMux I__1337 (
            .O(N__10042),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1336 (
            .O(N__10039),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__1335 (
            .O(N__10036),
            .I(\uu2.r_addrZ0Z_7 ));
    CascadeMux I__1334 (
            .O(N__10029),
            .I(N__10025));
    CascadeMux I__1333 (
            .O(N__10028),
            .I(N__10021));
    InMux I__1332 (
            .O(N__10025),
            .I(N__10017));
    InMux I__1331 (
            .O(N__10024),
            .I(N__10010));
    InMux I__1330 (
            .O(N__10021),
            .I(N__10010));
    InMux I__1329 (
            .O(N__10020),
            .I(N__10010));
    LocalMux I__1328 (
            .O(N__10017),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__1327 (
            .O(N__10010),
            .I(\uu2.r_addrZ0Z_6 ));
    InMux I__1326 (
            .O(N__10005),
            .I(N__10002));
    LocalMux I__1325 (
            .O(N__10002),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    InMux I__1324 (
            .O(N__9999),
            .I(N__9996));
    LocalMux I__1323 (
            .O(N__9996),
            .I(\uu2.mem0.w_data_6 ));
    InMux I__1322 (
            .O(N__9993),
            .I(N__9990));
    LocalMux I__1321 (
            .O(N__9990),
            .I(\uu2.mem0.w_data_5 ));
    InMux I__1320 (
            .O(N__9987),
            .I(N__9984));
    LocalMux I__1319 (
            .O(N__9984),
            .I(\uu2.N_34 ));
    CascadeMux I__1318 (
            .O(N__9981),
            .I(\uu2.N_34_cascade_ ));
    InMux I__1317 (
            .O(N__9978),
            .I(N__9975));
    LocalMux I__1316 (
            .O(N__9975),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__1315 (
            .O(N__9972),
            .I(N__9969));
    LocalMux I__1314 (
            .O(N__9969),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__1313 (
            .O(N__9966),
            .I(N__9963));
    LocalMux I__1312 (
            .O(N__9963),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__1311 (
            .O(N__9960),
            .I(N__9955));
    InMux I__1310 (
            .O(N__9959),
            .I(N__9952));
    InMux I__1309 (
            .O(N__9958),
            .I(N__9949));
    LocalMux I__1308 (
            .O(N__9955),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1307 (
            .O(N__9952),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__1306 (
            .O(N__9949),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    InMux I__1305 (
            .O(N__9942),
            .I(N__9939));
    LocalMux I__1304 (
            .O(N__9939),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__1303 (
            .O(N__9936),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1302 (
            .O(N__9933),
            .I(N__9929));
    InMux I__1301 (
            .O(N__9932),
            .I(N__9926));
    LocalMux I__1300 (
            .O(N__9929),
            .I(N__9923));
    LocalMux I__1299 (
            .O(N__9926),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    Odrv4 I__1298 (
            .O(N__9923),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    InMux I__1297 (
            .O(N__9918),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    CascadeMux I__1296 (
            .O(N__9915),
            .I(N__9912));
    InMux I__1295 (
            .O(N__9912),
            .I(N__9907));
    InMux I__1294 (
            .O(N__9911),
            .I(N__9904));
    InMux I__1293 (
            .O(N__9910),
            .I(N__9901));
    LocalMux I__1292 (
            .O(N__9907),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1291 (
            .O(N__9904),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__1290 (
            .O(N__9901),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__1289 (
            .O(N__9894),
            .I(N__9891));
    LocalMux I__1288 (
            .O(N__9891),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    InMux I__1287 (
            .O(N__9888),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__1286 (
            .O(N__9885),
            .I(N__9879));
    InMux I__1285 (
            .O(N__9884),
            .I(N__9872));
    InMux I__1284 (
            .O(N__9883),
            .I(N__9872));
    InMux I__1283 (
            .O(N__9882),
            .I(N__9872));
    LocalMux I__1282 (
            .O(N__9879),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__1281 (
            .O(N__9872),
            .I(\buart.Z_rx.ser_clk ));
    CascadeMux I__1280 (
            .O(N__9867),
            .I(N__9861));
    InMux I__1279 (
            .O(N__9866),
            .I(N__9855));
    InMux I__1278 (
            .O(N__9865),
            .I(N__9852));
    InMux I__1277 (
            .O(N__9864),
            .I(N__9849));
    InMux I__1276 (
            .O(N__9861),
            .I(N__9841));
    InMux I__1275 (
            .O(N__9860),
            .I(N__9838));
    InMux I__1274 (
            .O(N__9859),
            .I(N__9833));
    InMux I__1273 (
            .O(N__9858),
            .I(N__9833));
    LocalMux I__1272 (
            .O(N__9855),
            .I(N__9826));
    LocalMux I__1271 (
            .O(N__9852),
            .I(N__9826));
    LocalMux I__1270 (
            .O(N__9849),
            .I(N__9826));
    InMux I__1269 (
            .O(N__9848),
            .I(N__9815));
    InMux I__1268 (
            .O(N__9847),
            .I(N__9815));
    InMux I__1267 (
            .O(N__9846),
            .I(N__9815));
    InMux I__1266 (
            .O(N__9845),
            .I(N__9815));
    InMux I__1265 (
            .O(N__9844),
            .I(N__9815));
    LocalMux I__1264 (
            .O(N__9841),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__1263 (
            .O(N__9838),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__1262 (
            .O(N__9833),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__1261 (
            .O(N__9826),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__1260 (
            .O(N__9815),
            .I(\buart.Z_rx.startbit ));
    InMux I__1259 (
            .O(N__9804),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    CascadeMux I__1258 (
            .O(N__9801),
            .I(N__9797));
    CascadeMux I__1257 (
            .O(N__9800),
            .I(N__9794));
    InMux I__1256 (
            .O(N__9797),
            .I(N__9791));
    InMux I__1255 (
            .O(N__9794),
            .I(N__9788));
    LocalMux I__1254 (
            .O(N__9791),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__1253 (
            .O(N__9788),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__1252 (
            .O(N__9783),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__1251 (
            .O(N__9780),
            .I(N__9777));
    InMux I__1250 (
            .O(N__9777),
            .I(N__9773));
    InMux I__1249 (
            .O(N__9776),
            .I(N__9770));
    LocalMux I__1248 (
            .O(N__9773),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__1247 (
            .O(N__9770),
            .I(\uu2.r_addrZ0Z_8 ));
    InMux I__1246 (
            .O(N__9765),
            .I(N__9762));
    LocalMux I__1245 (
            .O(N__9762),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__1244 (
            .O(N__9759),
            .I(N__9754));
    CascadeMux I__1243 (
            .O(N__9758),
            .I(N__9751));
    CascadeMux I__1242 (
            .O(N__9757),
            .I(N__9748));
    InMux I__1241 (
            .O(N__9754),
            .I(N__9745));
    InMux I__1240 (
            .O(N__9751),
            .I(N__9740));
    InMux I__1239 (
            .O(N__9748),
            .I(N__9740));
    LocalMux I__1238 (
            .O(N__9745),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__1237 (
            .O(N__9740),
            .I(\uu2.r_addrZ0Z_3 ));
    InMux I__1236 (
            .O(N__9735),
            .I(N__9732));
    LocalMux I__1235 (
            .O(N__9732),
            .I(N__9729));
    Odrv4 I__1234 (
            .O(N__9729),
            .I(\buart.Z_rx.un1_sample_0 ));
    InMux I__1233 (
            .O(N__9726),
            .I(N__9720));
    InMux I__1232 (
            .O(N__9725),
            .I(N__9716));
    InMux I__1231 (
            .O(N__9724),
            .I(N__9711));
    InMux I__1230 (
            .O(N__9723),
            .I(N__9711));
    LocalMux I__1229 (
            .O(N__9720),
            .I(N__9708));
    InMux I__1228 (
            .O(N__9719),
            .I(N__9705));
    LocalMux I__1227 (
            .O(N__9716),
            .I(N__9700));
    LocalMux I__1226 (
            .O(N__9711),
            .I(N__9700));
    Odrv4 I__1225 (
            .O(N__9708),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__1224 (
            .O(N__9705),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    Odrv4 I__1223 (
            .O(N__9700),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    IoInMux I__1222 (
            .O(N__9693),
            .I(N__9690));
    LocalMux I__1221 (
            .O(N__9690),
            .I(N__9687));
    Span4Mux_s2_v I__1220 (
            .O(N__9687),
            .I(N__9684));
    Span4Mux_h I__1219 (
            .O(N__9684),
            .I(N__9681));
    Odrv4 I__1218 (
            .O(N__9681),
            .I(\buart.Z_rx.sample ));
    CascadeMux I__1217 (
            .O(N__9678),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    CascadeMux I__1216 (
            .O(N__9675),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    CascadeMux I__1215 (
            .O(N__9672),
            .I(N__9669));
    InMux I__1214 (
            .O(N__9669),
            .I(N__9664));
    InMux I__1213 (
            .O(N__9668),
            .I(N__9659));
    InMux I__1212 (
            .O(N__9667),
            .I(N__9659));
    LocalMux I__1211 (
            .O(N__9664),
            .I(\buart.Z_rx.idle ));
    LocalMux I__1210 (
            .O(N__9659),
            .I(\buart.Z_rx.idle ));
    CEMux I__1209 (
            .O(N__9654),
            .I(N__9648));
    CEMux I__1208 (
            .O(N__9653),
            .I(N__9645));
    CEMux I__1207 (
            .O(N__9652),
            .I(N__9642));
    CEMux I__1206 (
            .O(N__9651),
            .I(N__9639));
    LocalMux I__1205 (
            .O(N__9648),
            .I(N__9634));
    LocalMux I__1204 (
            .O(N__9645),
            .I(N__9634));
    LocalMux I__1203 (
            .O(N__9642),
            .I(N__9631));
    LocalMux I__1202 (
            .O(N__9639),
            .I(N__9628));
    Odrv4 I__1201 (
            .O(N__9634),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv12 I__1200 (
            .O(N__9631),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv4 I__1199 (
            .O(N__9628),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__1198 (
            .O(N__9621),
            .I(N__9616));
    InMux I__1197 (
            .O(N__9620),
            .I(N__9611));
    InMux I__1196 (
            .O(N__9619),
            .I(N__9611));
    LocalMux I__1195 (
            .O(N__9616),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__1194 (
            .O(N__9611),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__1193 (
            .O(N__9606),
            .I(N__9602));
    CascadeMux I__1192 (
            .O(N__9605),
            .I(N__9599));
    InMux I__1191 (
            .O(N__9602),
            .I(N__9594));
    InMux I__1190 (
            .O(N__9599),
            .I(N__9587));
    InMux I__1189 (
            .O(N__9598),
            .I(N__9587));
    InMux I__1188 (
            .O(N__9597),
            .I(N__9587));
    LocalMux I__1187 (
            .O(N__9594),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__1186 (
            .O(N__9587),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__1185 (
            .O(N__9582),
            .I(N__9579));
    InMux I__1184 (
            .O(N__9579),
            .I(N__9576));
    LocalMux I__1183 (
            .O(N__9576),
            .I(N__9573));
    Span12Mux_s9_v I__1182 (
            .O(N__9573),
            .I(N__9570));
    Odrv12 I__1181 (
            .O(N__9570),
            .I(\uu2.mem0.w_addr_0 ));
    InMux I__1180 (
            .O(N__9567),
            .I(N__9563));
    InMux I__1179 (
            .O(N__9566),
            .I(N__9560));
    LocalMux I__1178 (
            .O(N__9563),
            .I(N__9557));
    LocalMux I__1177 (
            .O(N__9560),
            .I(N__9552));
    Span4Mux_v I__1176 (
            .O(N__9557),
            .I(N__9552));
    Odrv4 I__1175 (
            .O(N__9552),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    CascadeMux I__1174 (
            .O(N__9549),
            .I(N__9546));
    InMux I__1173 (
            .O(N__9546),
            .I(N__9542));
    CascadeMux I__1172 (
            .O(N__9545),
            .I(N__9537));
    LocalMux I__1171 (
            .O(N__9542),
            .I(N__9533));
    InMux I__1170 (
            .O(N__9541),
            .I(N__9530));
    InMux I__1169 (
            .O(N__9540),
            .I(N__9527));
    InMux I__1168 (
            .O(N__9537),
            .I(N__9522));
    InMux I__1167 (
            .O(N__9536),
            .I(N__9522));
    Odrv4 I__1166 (
            .O(N__9533),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1165 (
            .O(N__9530),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1164 (
            .O(N__9527),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__1163 (
            .O(N__9522),
            .I(\buart.Z_rx.N_27_0_i ));
    CascadeMux I__1162 (
            .O(N__9513),
            .I(\resetGen.un241_ci_cascade_ ));
    InMux I__1161 (
            .O(N__9510),
            .I(N__9505));
    InMux I__1160 (
            .O(N__9509),
            .I(N__9500));
    InMux I__1159 (
            .O(N__9508),
            .I(N__9500));
    LocalMux I__1158 (
            .O(N__9505),
            .I(\resetGen.reset_countZ0Z_1 ));
    LocalMux I__1157 (
            .O(N__9500),
            .I(\resetGen.reset_countZ0Z_1 ));
    CascadeMux I__1156 (
            .O(N__9495),
            .I(N__9492));
    InMux I__1155 (
            .O(N__9492),
            .I(N__9484));
    InMux I__1154 (
            .O(N__9491),
            .I(N__9484));
    InMux I__1153 (
            .O(N__9490),
            .I(N__9479));
    InMux I__1152 (
            .O(N__9489),
            .I(N__9479));
    LocalMux I__1151 (
            .O(N__9484),
            .I(\resetGen.reset_countZ0Z_0 ));
    LocalMux I__1150 (
            .O(N__9479),
            .I(\resetGen.reset_countZ0Z_0 ));
    CascadeMux I__1149 (
            .O(N__9474),
            .I(\resetGen.un252_ci_cascade_ ));
    InMux I__1148 (
            .O(N__9471),
            .I(N__9465));
    InMux I__1147 (
            .O(N__9470),
            .I(N__9465));
    LocalMux I__1146 (
            .O(N__9465),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__1145 (
            .O(N__9462),
            .I(N__9453));
    InMux I__1144 (
            .O(N__9461),
            .I(N__9453));
    InMux I__1143 (
            .O(N__9460),
            .I(N__9453));
    LocalMux I__1142 (
            .O(N__9453),
            .I(\resetGen.reset_countZ0Z_2 ));
    InMux I__1141 (
            .O(N__9450),
            .I(N__9447));
    LocalMux I__1140 (
            .O(N__9447),
            .I(\resetGen.un241_ci ));
    CascadeMux I__1139 (
            .O(N__9444),
            .I(\resetGen.reset_count_2_0_4_cascade_ ));
    InMux I__1138 (
            .O(N__9441),
            .I(N__9431));
    InMux I__1137 (
            .O(N__9440),
            .I(N__9431));
    InMux I__1136 (
            .O(N__9439),
            .I(N__9424));
    InMux I__1135 (
            .O(N__9438),
            .I(N__9424));
    InMux I__1134 (
            .O(N__9437),
            .I(N__9424));
    InMux I__1133 (
            .O(N__9436),
            .I(N__9421));
    LocalMux I__1132 (
            .O(N__9431),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__1131 (
            .O(N__9424),
            .I(\resetGen.reset_countZ0Z_4 ));
    LocalMux I__1130 (
            .O(N__9421),
            .I(\resetGen.reset_countZ0Z_4 ));
    InMux I__1129 (
            .O(N__9414),
            .I(N__9410));
    InMux I__1128 (
            .O(N__9413),
            .I(N__9407));
    LocalMux I__1127 (
            .O(N__9410),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__1126 (
            .O(N__9407),
            .I(\uu0.l_countZ0Z_18 ));
    CascadeMux I__1125 (
            .O(N__9402),
            .I(N__9399));
    InMux I__1124 (
            .O(N__9399),
            .I(N__9394));
    InMux I__1123 (
            .O(N__9398),
            .I(N__9391));
    InMux I__1122 (
            .O(N__9397),
            .I(N__9388));
    LocalMux I__1121 (
            .O(N__9394),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__1120 (
            .O(N__9391),
            .I(\uu0.l_countZ0Z_15 ));
    LocalMux I__1119 (
            .O(N__9388),
            .I(\uu0.l_countZ0Z_15 ));
    CascadeMux I__1118 (
            .O(N__9381),
            .I(\uu0.un4_l_count_11_cascade_ ));
    InMux I__1117 (
            .O(N__9378),
            .I(N__9368));
    InMux I__1116 (
            .O(N__9377),
            .I(N__9368));
    InMux I__1115 (
            .O(N__9376),
            .I(N__9368));
    InMux I__1114 (
            .O(N__9375),
            .I(N__9365));
    LocalMux I__1113 (
            .O(N__9368),
            .I(\uu0.l_countZ0Z_6 ));
    LocalMux I__1112 (
            .O(N__9365),
            .I(\uu0.l_countZ0Z_6 ));
    InMux I__1111 (
            .O(N__9360),
            .I(N__9357));
    LocalMux I__1110 (
            .O(N__9357),
            .I(\uu0.un4_l_count_16 ));
    InMux I__1109 (
            .O(N__9354),
            .I(N__9347));
    InMux I__1108 (
            .O(N__9353),
            .I(N__9340));
    InMux I__1107 (
            .O(N__9352),
            .I(N__9340));
    InMux I__1106 (
            .O(N__9351),
            .I(N__9340));
    InMux I__1105 (
            .O(N__9350),
            .I(N__9336));
    LocalMux I__1104 (
            .O(N__9347),
            .I(N__9331));
    LocalMux I__1103 (
            .O(N__9340),
            .I(N__9331));
    InMux I__1102 (
            .O(N__9339),
            .I(N__9328));
    LocalMux I__1101 (
            .O(N__9336),
            .I(N__9325));
    Odrv12 I__1100 (
            .O(N__9331),
            .I(\uu0.l_precountZ0Z_0 ));
    LocalMux I__1099 (
            .O(N__9328),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__1098 (
            .O(N__9325),
            .I(\uu0.l_precountZ0Z_0 ));
    CascadeMux I__1097 (
            .O(N__9318),
            .I(N__9314));
    InMux I__1096 (
            .O(N__9317),
            .I(N__9308));
    InMux I__1095 (
            .O(N__9314),
            .I(N__9301));
    InMux I__1094 (
            .O(N__9313),
            .I(N__9301));
    InMux I__1093 (
            .O(N__9312),
            .I(N__9301));
    InMux I__1092 (
            .O(N__9311),
            .I(N__9298));
    LocalMux I__1091 (
            .O(N__9308),
            .I(\uu0.l_precountZ0Z_1 ));
    LocalMux I__1090 (
            .O(N__9301),
            .I(\uu0.l_precountZ0Z_1 ));
    LocalMux I__1089 (
            .O(N__9298),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__1088 (
            .O(N__9291),
            .I(CONSTANT_ONE_NET_cascade_));
    InMux I__1087 (
            .O(N__9288),
            .I(N__9285));
    LocalMux I__1086 (
            .O(N__9285),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1085 (
            .O(N__9282),
            .I(N__9272));
    InMux I__1084 (
            .O(N__9281),
            .I(N__9272));
    InMux I__1083 (
            .O(N__9280),
            .I(N__9272));
    InMux I__1082 (
            .O(N__9279),
            .I(N__9269));
    LocalMux I__1081 (
            .O(N__9272),
            .I(N__9265));
    LocalMux I__1080 (
            .O(N__9269),
            .I(N__9262));
    InMux I__1079 (
            .O(N__9268),
            .I(N__9259));
    Span4Mux_v I__1078 (
            .O(N__9265),
            .I(N__9256));
    Odrv4 I__1077 (
            .O(N__9262),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1076 (
            .O(N__9259),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    Odrv4 I__1075 (
            .O(N__9256),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    InMux I__1074 (
            .O(N__9249),
            .I(N__9246));
    LocalMux I__1073 (
            .O(N__9246),
            .I(N__9243));
    Odrv4 I__1072 (
            .O(N__9243),
            .I(\uu0.delay_lineZ0Z_1 ));
    InMux I__1071 (
            .O(N__9240),
            .I(N__9236));
    InMux I__1070 (
            .O(N__9239),
            .I(N__9233));
    LocalMux I__1069 (
            .O(N__9236),
            .I(N__9230));
    LocalMux I__1068 (
            .O(N__9233),
            .I(\uu0.delay_lineZ0Z_0 ));
    Odrv4 I__1067 (
            .O(N__9230),
            .I(\uu0.delay_lineZ0Z_0 ));
    InMux I__1066 (
            .O(N__9225),
            .I(N__9210));
    InMux I__1065 (
            .O(N__9224),
            .I(N__9203));
    InMux I__1064 (
            .O(N__9223),
            .I(N__9203));
    InMux I__1063 (
            .O(N__9222),
            .I(N__9203));
    InMux I__1062 (
            .O(N__9221),
            .I(N__9200));
    InMux I__1061 (
            .O(N__9220),
            .I(N__9197));
    InMux I__1060 (
            .O(N__9219),
            .I(N__9192));
    InMux I__1059 (
            .O(N__9218),
            .I(N__9192));
    InMux I__1058 (
            .O(N__9217),
            .I(N__9189));
    InMux I__1057 (
            .O(N__9216),
            .I(N__9186));
    InMux I__1056 (
            .O(N__9215),
            .I(N__9183));
    InMux I__1055 (
            .O(N__9214),
            .I(N__9178));
    InMux I__1054 (
            .O(N__9213),
            .I(N__9178));
    LocalMux I__1053 (
            .O(N__9210),
            .I(N__9175));
    LocalMux I__1052 (
            .O(N__9203),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1051 (
            .O(N__9200),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1050 (
            .O(N__9197),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1049 (
            .O(N__9192),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1048 (
            .O(N__9189),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1047 (
            .O(N__9186),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1046 (
            .O(N__9183),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1045 (
            .O(N__9178),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1044 (
            .O(N__9175),
            .I(\uu0.un4_l_count_0 ));
    IoInMux I__1043 (
            .O(N__9156),
            .I(N__9153));
    LocalMux I__1042 (
            .O(N__9153),
            .I(N__9150));
    Span4Mux_s1_h I__1041 (
            .O(N__9150),
            .I(N__9147));
    Odrv4 I__1040 (
            .O(N__9147),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__1039 (
            .O(N__9144),
            .I(\uu0.un143_ci_0_cascade_ ));
    CascadeMux I__1038 (
            .O(N__9141),
            .I(N__9131));
    CascadeMux I__1037 (
            .O(N__9140),
            .I(N__9128));
    CascadeMux I__1036 (
            .O(N__9139),
            .I(N__9125));
    InMux I__1035 (
            .O(N__9138),
            .I(N__9118));
    InMux I__1034 (
            .O(N__9137),
            .I(N__9118));
    InMux I__1033 (
            .O(N__9136),
            .I(N__9109));
    InMux I__1032 (
            .O(N__9135),
            .I(N__9109));
    InMux I__1031 (
            .O(N__9134),
            .I(N__9109));
    InMux I__1030 (
            .O(N__9131),
            .I(N__9109));
    InMux I__1029 (
            .O(N__9128),
            .I(N__9100));
    InMux I__1028 (
            .O(N__9125),
            .I(N__9100));
    InMux I__1027 (
            .O(N__9124),
            .I(N__9100));
    InMux I__1026 (
            .O(N__9123),
            .I(N__9100));
    LocalMux I__1025 (
            .O(N__9118),
            .I(\uu0.un110_ci ));
    LocalMux I__1024 (
            .O(N__9109),
            .I(\uu0.un110_ci ));
    LocalMux I__1023 (
            .O(N__9100),
            .I(\uu0.un110_ci ));
    InMux I__1022 (
            .O(N__9093),
            .I(N__9085));
    InMux I__1021 (
            .O(N__9092),
            .I(N__9074));
    InMux I__1020 (
            .O(N__9091),
            .I(N__9074));
    InMux I__1019 (
            .O(N__9090),
            .I(N__9074));
    InMux I__1018 (
            .O(N__9089),
            .I(N__9074));
    InMux I__1017 (
            .O(N__9088),
            .I(N__9074));
    LocalMux I__1016 (
            .O(N__9085),
            .I(\uu0.l_countZ0Z_8 ));
    LocalMux I__1015 (
            .O(N__9074),
            .I(\uu0.l_countZ0Z_8 ));
    CEMux I__1014 (
            .O(N__9069),
            .I(N__9057));
    CEMux I__1013 (
            .O(N__9068),
            .I(N__9057));
    CEMux I__1012 (
            .O(N__9067),
            .I(N__9057));
    CEMux I__1011 (
            .O(N__9066),
            .I(N__9057));
    GlobalMux I__1010 (
            .O(N__9057),
            .I(N__9054));
    gio2CtrlBuf I__1009 (
            .O(N__9054),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__1008 (
            .O(N__9051),
            .I(N__9046));
    CascadeMux I__1007 (
            .O(N__9050),
            .I(N__9042));
    InMux I__1006 (
            .O(N__9049),
            .I(N__9039));
    InMux I__1005 (
            .O(N__9046),
            .I(N__9032));
    InMux I__1004 (
            .O(N__9045),
            .I(N__9032));
    InMux I__1003 (
            .O(N__9042),
            .I(N__9032));
    LocalMux I__1002 (
            .O(N__9039),
            .I(N__9029));
    LocalMux I__1001 (
            .O(N__9032),
            .I(\uu0.l_countZ0Z_16 ));
    Odrv4 I__1000 (
            .O(N__9029),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__999 (
            .O(N__9024),
            .I(N__9020));
    InMux I__998 (
            .O(N__9023),
            .I(N__9016));
    InMux I__997 (
            .O(N__9020),
            .I(N__9013));
    InMux I__996 (
            .O(N__9019),
            .I(N__9010));
    LocalMux I__995 (
            .O(N__9016),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__994 (
            .O(N__9013),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__993 (
            .O(N__9010),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__992 (
            .O(N__9003),
            .I(N__8996));
    CascadeMux I__991 (
            .O(N__9002),
            .I(N__8993));
    InMux I__990 (
            .O(N__9001),
            .I(N__8984));
    InMux I__989 (
            .O(N__9000),
            .I(N__8984));
    InMux I__988 (
            .O(N__8999),
            .I(N__8984));
    InMux I__987 (
            .O(N__8996),
            .I(N__8984));
    InMux I__986 (
            .O(N__8993),
            .I(N__8981));
    LocalMux I__985 (
            .O(N__8984),
            .I(\uu0.l_countZ0Z_0 ));
    LocalMux I__984 (
            .O(N__8981),
            .I(\uu0.l_countZ0Z_0 ));
    InMux I__983 (
            .O(N__8976),
            .I(N__8973));
    LocalMux I__982 (
            .O(N__8973),
            .I(\uu0.un4_l_count_12 ));
    InMux I__981 (
            .O(N__8970),
            .I(N__8967));
    LocalMux I__980 (
            .O(N__8967),
            .I(\uu0.un4_l_count_18 ));
    CascadeMux I__979 (
            .O(N__8964),
            .I(\uu0.un4_l_count_13_cascade_ ));
    CascadeMux I__978 (
            .O(N__8961),
            .I(N__8957));
    InMux I__977 (
            .O(N__8960),
            .I(N__8946));
    InMux I__976 (
            .O(N__8957),
            .I(N__8946));
    InMux I__975 (
            .O(N__8956),
            .I(N__8946));
    InMux I__974 (
            .O(N__8955),
            .I(N__8946));
    LocalMux I__973 (
            .O(N__8946),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__972 (
            .O(N__8943),
            .I(N__8936));
    InMux I__971 (
            .O(N__8942),
            .I(N__8936));
    InMux I__970 (
            .O(N__8941),
            .I(N__8933));
    LocalMux I__969 (
            .O(N__8936),
            .I(\uu0.l_countZ0Z_5 ));
    LocalMux I__968 (
            .O(N__8933),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__967 (
            .O(N__8928),
            .I(N__8923));
    CascadeMux I__966 (
            .O(N__8927),
            .I(N__8920));
    InMux I__965 (
            .O(N__8926),
            .I(N__8913));
    InMux I__964 (
            .O(N__8923),
            .I(N__8913));
    InMux I__963 (
            .O(N__8920),
            .I(N__8913));
    LocalMux I__962 (
            .O(N__8913),
            .I(\uu0.l_precountZ0Z_3 ));
    InMux I__961 (
            .O(N__8910),
            .I(N__8900));
    InMux I__960 (
            .O(N__8909),
            .I(N__8900));
    InMux I__959 (
            .O(N__8908),
            .I(N__8900));
    InMux I__958 (
            .O(N__8907),
            .I(N__8897));
    LocalMux I__957 (
            .O(N__8900),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__956 (
            .O(N__8897),
            .I(\uu0.l_countZ0Z_1 ));
    InMux I__955 (
            .O(N__8892),
            .I(N__8889));
    LocalMux I__954 (
            .O(N__8889),
            .I(\uu0.un187_ci_1 ));
    InMux I__953 (
            .O(N__8886),
            .I(N__8877));
    InMux I__952 (
            .O(N__8885),
            .I(N__8877));
    InMux I__951 (
            .O(N__8884),
            .I(N__8877));
    LocalMux I__950 (
            .O(N__8877),
            .I(\uu2.l_countZ0Z_3 ));
    InMux I__949 (
            .O(N__8874),
            .I(N__8863));
    InMux I__948 (
            .O(N__8873),
            .I(N__8863));
    InMux I__947 (
            .O(N__8872),
            .I(N__8863));
    InMux I__946 (
            .O(N__8871),
            .I(N__8858));
    InMux I__945 (
            .O(N__8870),
            .I(N__8858));
    LocalMux I__944 (
            .O(N__8863),
            .I(N__8855));
    LocalMux I__943 (
            .O(N__8858),
            .I(\uu2.l_countZ0Z_2 ));
    Odrv4 I__942 (
            .O(N__8855),
            .I(\uu2.l_countZ0Z_2 ));
    CascadeMux I__941 (
            .O(N__8850),
            .I(N__8847));
    InMux I__940 (
            .O(N__8847),
            .I(N__8841));
    InMux I__939 (
            .O(N__8846),
            .I(N__8838));
    InMux I__938 (
            .O(N__8845),
            .I(N__8833));
    InMux I__937 (
            .O(N__8844),
            .I(N__8833));
    LocalMux I__936 (
            .O(N__8841),
            .I(N__8828));
    LocalMux I__935 (
            .O(N__8838),
            .I(N__8828));
    LocalMux I__934 (
            .O(N__8833),
            .I(\uu0.l_countZ0Z_2 ));
    Odrv4 I__933 (
            .O(N__8828),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__932 (
            .O(N__8823),
            .I(\uu0.un4_l_count_14_cascade_ ));
    CascadeMux I__931 (
            .O(N__8820),
            .I(N__8816));
    InMux I__930 (
            .O(N__8819),
            .I(N__8811));
    InMux I__929 (
            .O(N__8816),
            .I(N__8804));
    InMux I__928 (
            .O(N__8815),
            .I(N__8804));
    InMux I__927 (
            .O(N__8814),
            .I(N__8804));
    LocalMux I__926 (
            .O(N__8811),
            .I(N__8801));
    LocalMux I__925 (
            .O(N__8804),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__924 (
            .O(N__8801),
            .I(\uu0.l_countZ0Z_4 ));
    CascadeMux I__923 (
            .O(N__8796),
            .I(N__8790));
    InMux I__922 (
            .O(N__8795),
            .I(N__8787));
    InMux I__921 (
            .O(N__8794),
            .I(N__8784));
    InMux I__920 (
            .O(N__8793),
            .I(N__8779));
    InMux I__919 (
            .O(N__8790),
            .I(N__8779));
    LocalMux I__918 (
            .O(N__8787),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__917 (
            .O(N__8784),
            .I(\uu0.un154_ci_9 ));
    LocalMux I__916 (
            .O(N__8779),
            .I(\uu0.un154_ci_9 ));
    InMux I__915 (
            .O(N__8772),
            .I(N__8764));
    InMux I__914 (
            .O(N__8771),
            .I(N__8764));
    InMux I__913 (
            .O(N__8770),
            .I(N__8759));
    InMux I__912 (
            .O(N__8769),
            .I(N__8759));
    LocalMux I__911 (
            .O(N__8764),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__910 (
            .O(N__8759),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__909 (
            .O(N__8754),
            .I(\uu0.un154_ci_9_cascade_ ));
    CascadeMux I__908 (
            .O(N__8751),
            .I(N__8745));
    InMux I__907 (
            .O(N__8750),
            .I(N__8742));
    InMux I__906 (
            .O(N__8749),
            .I(N__8739));
    InMux I__905 (
            .O(N__8748),
            .I(N__8736));
    InMux I__904 (
            .O(N__8745),
            .I(N__8733));
    LocalMux I__903 (
            .O(N__8742),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__902 (
            .O(N__8739),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__901 (
            .O(N__8736),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__900 (
            .O(N__8733),
            .I(\uu0.l_countZ0Z_14 ));
    CascadeMux I__899 (
            .O(N__8724),
            .I(N__8721));
    InMux I__898 (
            .O(N__8721),
            .I(N__8710));
    InMux I__897 (
            .O(N__8720),
            .I(N__8710));
    InMux I__896 (
            .O(N__8719),
            .I(N__8710));
    InMux I__895 (
            .O(N__8718),
            .I(N__8705));
    InMux I__894 (
            .O(N__8717),
            .I(N__8705));
    LocalMux I__893 (
            .O(N__8710),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__892 (
            .O(N__8705),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__891 (
            .O(N__8700),
            .I(N__8688));
    InMux I__890 (
            .O(N__8699),
            .I(N__8688));
    InMux I__889 (
            .O(N__8698),
            .I(N__8688));
    InMux I__888 (
            .O(N__8697),
            .I(N__8688));
    LocalMux I__887 (
            .O(N__8688),
            .I(\uu0.l_countZ0Z_10 ));
    CascadeMux I__886 (
            .O(N__8685),
            .I(\uu2.vbuf_count.un328_ci_3_cascade_ ));
    CascadeMux I__885 (
            .O(N__8682),
            .I(N__8677));
    InMux I__884 (
            .O(N__8681),
            .I(N__8674));
    InMux I__883 (
            .O(N__8680),
            .I(N__8669));
    InMux I__882 (
            .O(N__8677),
            .I(N__8669));
    LocalMux I__881 (
            .O(N__8674),
            .I(\uu2.l_countZ0Z_9 ));
    LocalMux I__880 (
            .O(N__8669),
            .I(\uu2.l_countZ0Z_9 ));
    CascadeMux I__879 (
            .O(N__8664),
            .I(N__8658));
    InMux I__878 (
            .O(N__8663),
            .I(N__8646));
    InMux I__877 (
            .O(N__8662),
            .I(N__8646));
    InMux I__876 (
            .O(N__8661),
            .I(N__8646));
    InMux I__875 (
            .O(N__8658),
            .I(N__8646));
    InMux I__874 (
            .O(N__8657),
            .I(N__8646));
    LocalMux I__873 (
            .O(N__8646),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__872 (
            .O(N__8643),
            .I(N__8636));
    InMux I__871 (
            .O(N__8642),
            .I(N__8636));
    InMux I__870 (
            .O(N__8641),
            .I(N__8633));
    LocalMux I__869 (
            .O(N__8636),
            .I(\uu2.l_countZ0Z_5 ));
    LocalMux I__868 (
            .O(N__8633),
            .I(\uu2.l_countZ0Z_5 ));
    CascadeMux I__867 (
            .O(N__8628),
            .I(N__8625));
    InMux I__866 (
            .O(N__8625),
            .I(N__8620));
    InMux I__865 (
            .O(N__8624),
            .I(N__8617));
    InMux I__864 (
            .O(N__8623),
            .I(N__8614));
    LocalMux I__863 (
            .O(N__8620),
            .I(N__8611));
    LocalMux I__862 (
            .O(N__8617),
            .I(\uu2.l_countZ0Z_8 ));
    LocalMux I__861 (
            .O(N__8614),
            .I(\uu2.l_countZ0Z_8 ));
    Odrv4 I__860 (
            .O(N__8611),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__859 (
            .O(N__8604),
            .I(\uu2.un1_l_count_1_3_cascade_ ));
    InMux I__858 (
            .O(N__8601),
            .I(N__8598));
    LocalMux I__857 (
            .O(N__8598),
            .I(\uu2.un1_l_count_1_2_0 ));
    InMux I__856 (
            .O(N__8595),
            .I(N__8591));
    InMux I__855 (
            .O(N__8594),
            .I(N__8588));
    LocalMux I__854 (
            .O(N__8591),
            .I(N__8585));
    LocalMux I__853 (
            .O(N__8588),
            .I(N__8582));
    Odrv4 I__852 (
            .O(N__8585),
            .I(\uu2.un1_l_count_1_0 ));
    Odrv4 I__851 (
            .O(N__8582),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__850 (
            .O(N__8577),
            .I(N__8568));
    InMux I__849 (
            .O(N__8576),
            .I(N__8568));
    InMux I__848 (
            .O(N__8575),
            .I(N__8568));
    LocalMux I__847 (
            .O(N__8568),
            .I(N__8565));
    Odrv4 I__846 (
            .O(N__8565),
            .I(\uu0.un198_ci_2 ));
    InMux I__845 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__844 (
            .O(N__8559),
            .I(\uu2.un1_l_count_1_3 ));
    CascadeMux I__843 (
            .O(N__8556),
            .I(N__8553));
    InMux I__842 (
            .O(N__8553),
            .I(N__8550));
    LocalMux I__841 (
            .O(N__8550),
            .I(\uu2.un1_l_count_2_2 ));
    InMux I__840 (
            .O(N__8547),
            .I(N__8542));
    InMux I__839 (
            .O(N__8546),
            .I(N__8537));
    InMux I__838 (
            .O(N__8545),
            .I(N__8537));
    LocalMux I__837 (
            .O(N__8542),
            .I(N__8534));
    LocalMux I__836 (
            .O(N__8537),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__835 (
            .O(N__8534),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__834 (
            .O(N__8529),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__833 (
            .O(N__8526),
            .I(N__8522));
    InMux I__832 (
            .O(N__8525),
            .I(N__8519));
    LocalMux I__831 (
            .O(N__8522),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    LocalMux I__830 (
            .O(N__8519),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    InMux I__829 (
            .O(N__8514),
            .I(N__8511));
    LocalMux I__828 (
            .O(N__8511),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__827 (
            .O(N__8508),
            .I(N__8505));
    LocalMux I__826 (
            .O(N__8505),
            .I(\uu2.un350_ci ));
    CascadeMux I__825 (
            .O(N__8502),
            .I(\uu2.un350_ci_cascade_ ));
    InMux I__824 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__823 (
            .O(N__8496),
            .I(vbuf_tx_data_0));
    InMux I__822 (
            .O(N__8493),
            .I(N__8490));
    LocalMux I__821 (
            .O(N__8490),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__820 (
            .O(N__8487),
            .I(N__8484));
    LocalMux I__819 (
            .O(N__8484),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__818 (
            .O(N__8481),
            .I(N__8478));
    LocalMux I__817 (
            .O(N__8478),
            .I(N__8475));
    Span12Mux_s1_h I__816 (
            .O(N__8475),
            .I(N__8472));
    Odrv12 I__815 (
            .O(N__8472),
            .I(o_serial_data_c));
    InMux I__814 (
            .O(N__8469),
            .I(N__8466));
    LocalMux I__813 (
            .O(N__8466),
            .I(vbuf_tx_data_1));
    InMux I__812 (
            .O(N__8463),
            .I(N__8460));
    LocalMux I__811 (
            .O(N__8460),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__810 (
            .O(N__8457),
            .I(N__8454));
    LocalMux I__809 (
            .O(N__8454),
            .I(vbuf_tx_data_2));
    InMux I__808 (
            .O(N__8451),
            .I(N__8448));
    LocalMux I__807 (
            .O(N__8448),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__806 (
            .O(N__8445),
            .I(N__8442));
    LocalMux I__805 (
            .O(N__8442),
            .I(vbuf_tx_data_3));
    InMux I__804 (
            .O(N__8439),
            .I(N__8436));
    LocalMux I__803 (
            .O(N__8436),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__802 (
            .O(N__8433),
            .I(N__8430));
    LocalMux I__801 (
            .O(N__8430),
            .I(vbuf_tx_data_4));
    InMux I__800 (
            .O(N__8427),
            .I(N__8424));
    LocalMux I__799 (
            .O(N__8424),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__798 (
            .O(N__8421),
            .I(N__8418));
    LocalMux I__797 (
            .O(N__8418),
            .I(vbuf_tx_data_5));
    InMux I__796 (
            .O(N__8415),
            .I(N__8412));
    LocalMux I__795 (
            .O(N__8412),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    InMux I__794 (
            .O(N__8409),
            .I(N__8406));
    LocalMux I__793 (
            .O(N__8406),
            .I(N__8403));
    Odrv4 I__792 (
            .O(N__8403),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__791 (
            .O(N__8400),
            .I(N__8396));
    InMux I__790 (
            .O(N__8399),
            .I(N__8390));
    LocalMux I__789 (
            .O(N__8396),
            .I(N__8387));
    InMux I__788 (
            .O(N__8395),
            .I(N__8380));
    InMux I__787 (
            .O(N__8394),
            .I(N__8380));
    InMux I__786 (
            .O(N__8393),
            .I(N__8380));
    LocalMux I__785 (
            .O(N__8390),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    Odrv4 I__784 (
            .O(N__8387),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__783 (
            .O(N__8380),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    InMux I__782 (
            .O(N__8373),
            .I(N__8370));
    LocalMux I__781 (
            .O(N__8370),
            .I(\uu2.r_data_wire_0 ));
    InMux I__780 (
            .O(N__8367),
            .I(N__8364));
    LocalMux I__779 (
            .O(N__8364),
            .I(\uu2.r_data_wire_1 ));
    InMux I__778 (
            .O(N__8361),
            .I(N__8358));
    LocalMux I__777 (
            .O(N__8358),
            .I(\uu2.r_data_wire_2 ));
    InMux I__776 (
            .O(N__8355),
            .I(N__8352));
    LocalMux I__775 (
            .O(N__8352),
            .I(\uu2.r_data_wire_3 ));
    InMux I__774 (
            .O(N__8349),
            .I(N__8346));
    LocalMux I__773 (
            .O(N__8346),
            .I(\uu2.r_data_wire_4 ));
    InMux I__772 (
            .O(N__8343),
            .I(N__8340));
    LocalMux I__771 (
            .O(N__8340),
            .I(\uu2.r_data_wire_5 ));
    InMux I__770 (
            .O(N__8337),
            .I(N__8334));
    LocalMux I__769 (
            .O(N__8334),
            .I(\uu2.r_data_wire_6 ));
    InMux I__768 (
            .O(N__8331),
            .I(N__8328));
    LocalMux I__767 (
            .O(N__8328),
            .I(\uu2.r_data_wire_7 ));
    InMux I__766 (
            .O(N__8325),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__765 (
            .O(N__8322),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__764 (
            .O(N__8319),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    CascadeMux I__763 (
            .O(N__8316),
            .I(\buart.Z_rx.valid_0_cascade_ ));
    CascadeMux I__762 (
            .O(N__8313),
            .I(N__8310));
    InMux I__761 (
            .O(N__8310),
            .I(N__8304));
    InMux I__760 (
            .O(N__8309),
            .I(N__8297));
    InMux I__759 (
            .O(N__8308),
            .I(N__8297));
    InMux I__758 (
            .O(N__8307),
            .I(N__8297));
    LocalMux I__757 (
            .O(N__8304),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__756 (
            .O(N__8297),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__755 (
            .O(N__8292),
            .I(\buart.Z_rx.idle_0_cascade_ ));
    InMux I__754 (
            .O(N__8289),
            .I(N__8286));
    LocalMux I__753 (
            .O(N__8286),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__752 (
            .O(N__8283),
            .I(N__8278));
    InMux I__751 (
            .O(N__8282),
            .I(N__8273));
    InMux I__750 (
            .O(N__8281),
            .I(N__8264));
    InMux I__749 (
            .O(N__8278),
            .I(N__8264));
    InMux I__748 (
            .O(N__8277),
            .I(N__8264));
    InMux I__747 (
            .O(N__8276),
            .I(N__8264));
    LocalMux I__746 (
            .O(N__8273),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__745 (
            .O(N__8264),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    CascadeMux I__744 (
            .O(N__8259),
            .I(N__8254));
    InMux I__743 (
            .O(N__8258),
            .I(N__8251));
    InMux I__742 (
            .O(N__8257),
            .I(N__8248));
    InMux I__741 (
            .O(N__8254),
            .I(N__8245));
    LocalMux I__740 (
            .O(N__8251),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__739 (
            .O(N__8248),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__738 (
            .O(N__8245),
            .I(\uu0.l_countZ0Z_3 ));
    CascadeMux I__737 (
            .O(N__8238),
            .I(\uu0.un66_ci_cascade_ ));
    CascadeMux I__736 (
            .O(N__8235),
            .I(N__8231));
    InMux I__735 (
            .O(N__8234),
            .I(N__8226));
    InMux I__734 (
            .O(N__8231),
            .I(N__8221));
    InMux I__733 (
            .O(N__8230),
            .I(N__8221));
    InMux I__732 (
            .O(N__8229),
            .I(N__8218));
    LocalMux I__731 (
            .O(N__8226),
            .I(N__8213));
    LocalMux I__730 (
            .O(N__8221),
            .I(N__8213));
    LocalMux I__729 (
            .O(N__8218),
            .I(\uu0.un66_ci ));
    Odrv4 I__728 (
            .O(N__8213),
            .I(\uu0.un66_ci ));
    CascadeMux I__727 (
            .O(N__8208),
            .I(N__8203));
    InMux I__726 (
            .O(N__8207),
            .I(N__8196));
    InMux I__725 (
            .O(N__8206),
            .I(N__8196));
    InMux I__724 (
            .O(N__8203),
            .I(N__8196));
    LocalMux I__723 (
            .O(N__8196),
            .I(N__8193));
    Odrv4 I__722 (
            .O(N__8193),
            .I(\uu0.un88_ci_3 ));
    InMux I__721 (
            .O(N__8190),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__720 (
            .O(N__8187),
            .I(N__8178));
    InMux I__719 (
            .O(N__8186),
            .I(N__8178));
    InMux I__718 (
            .O(N__8185),
            .I(N__8178));
    LocalMux I__717 (
            .O(N__8178),
            .I(\uu0.l_countZ0Z_17 ));
    CascadeMux I__716 (
            .O(N__8175),
            .I(\uu0.un220_ci_cascade_ ));
    CascadeMux I__715 (
            .O(N__8172),
            .I(N__8169));
    InMux I__714 (
            .O(N__8169),
            .I(N__8166));
    LocalMux I__713 (
            .O(N__8166),
            .I(\uu0.un99_ci_0 ));
    InMux I__712 (
            .O(N__8163),
            .I(N__8158));
    InMux I__711 (
            .O(N__8162),
            .I(N__8153));
    InMux I__710 (
            .O(N__8161),
            .I(N__8153));
    LocalMux I__709 (
            .O(N__8158),
            .I(\uu0.l_countZ0Z_7 ));
    LocalMux I__708 (
            .O(N__8153),
            .I(\uu0.l_countZ0Z_7 ));
    InMux I__707 (
            .O(N__8148),
            .I(N__8145));
    LocalMux I__706 (
            .O(N__8145),
            .I(\uu0.un44_ci ));
    CascadeMux I__705 (
            .O(N__8142),
            .I(\uu0.un44_ci_cascade_ ));
    CascadeMux I__704 (
            .O(N__8139),
            .I(\uu0.un165_ci_0_cascade_ ));
    InMux I__703 (
            .O(N__8136),
            .I(N__8130));
    InMux I__702 (
            .O(N__8135),
            .I(N__8130));
    LocalMux I__701 (
            .O(N__8130),
            .I(\uu0.l_countZ0Z_13 ));
    CascadeMux I__700 (
            .O(N__8127),
            .I(\uu0.un110_ci_cascade_ ));
    InMux I__699 (
            .O(N__8124),
            .I(N__8115));
    InMux I__698 (
            .O(N__8123),
            .I(N__8115));
    InMux I__697 (
            .O(N__8122),
            .I(N__8115));
    LocalMux I__696 (
            .O(N__8115),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__695 (
            .O(N__8112),
            .I(N__8109));
    LocalMux I__694 (
            .O(N__8109),
            .I(N__8106));
    IoSpan4Mux I__693 (
            .O(N__8106),
            .I(N__8103));
    IoSpan4Mux I__692 (
            .O(N__8103),
            .I(N__8100));
    Odrv4 I__691 (
            .O(N__8100),
            .I(uart_RXD));
    IoInMux I__690 (
            .O(N__8097),
            .I(N__8094));
    LocalMux I__689 (
            .O(N__8094),
            .I(N__8091));
    Span12Mux_s5_v I__688 (
            .O(N__8091),
            .I(N__8088));
    Odrv12 I__687 (
            .O(N__8088),
            .I(\latticehx1k_pll_inst.clk ));
    IoInMux I__686 (
            .O(N__8085),
            .I(N__8082));
    LocalMux I__685 (
            .O(N__8082),
            .I(N__8079));
    IoSpan4Mux I__684 (
            .O(N__8079),
            .I(N__8076));
    Odrv4 I__683 (
            .O(N__8076),
            .I(clk_in_c));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__22262));
    INV \INVuu2.w_addr_displaying_7C  (
            .O(\INVuu2.w_addr_displaying_7C_net ),
            .I(N__22266));
    INV \INVuu2.w_addr_user_nesr_3C  (
            .O(\INVuu2.w_addr_user_nesr_3C_net ),
            .I(N__22270));
    INV \INVuu2.bitmap_215C  (
            .O(\INVuu2.bitmap_215C_net ),
            .I(N__22248));
    INV \INVuu2.bitmap_290C  (
            .O(\INVuu2.bitmap_290C_net ),
            .I(N__22261));
    INV \INVuu2.w_addr_displaying_fast_8C  (
            .O(\INVuu2.w_addr_displaying_fast_8C_net ),
            .I(N__22265));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__22240));
    INV \INVuu2.bitmap_197C  (
            .O(\INVuu2.bitmap_197C_net ),
            .I(N__22247));
    INV \INVuu2.bitmap_168C  (
            .O(\INVuu2.bitmap_168C_net ),
            .I(N__22255));
    INV \INVuu2.w_addr_displaying_ness_6C  (
            .O(\INVuu2.w_addr_displaying_ness_6C_net ),
            .I(N__22260));
    INV \INVuu2.bitmap_93C  (
            .O(\INVuu2.bitmap_93C_net ),
            .I(N__22235));
    INV \INVuu2.w_addr_displaying_nesr_3C  (
            .O(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .I(N__22243));
    INV \INVuu2.w_addr_user_2C  (
            .O(\INVuu2.w_addr_user_2C_net ),
            .I(N__22250));
    INV \INVuu2.vram_rd_clk_det_1C  (
            .O(\INVuu2.vram_rd_clk_det_1C_net ),
            .I(N__22239));
    INV \INVuu2.w_addr_displaying_1_rep1_nesrC  (
            .O(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .I(N__22254));
    INV \INVuu2.vram_rd_clk_det_0C  (
            .O(\INVuu2.vram_rd_clk_det_0C_net ),
            .I(N__22246));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__22272));
    defparam IN_MUX_bfv_12_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_2_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_2_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_13_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__8097),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__9693),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__9156),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__14914),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \buart.Z_rx.hh_0_LC_1_6_4 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_6_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8112),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22251),
            .ce(),
            .sr(N__20679));
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_7_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_7_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_1_7_0  (
            .in0(_gnd_net_),
            .in1(N__8135),
            .in2(_gnd_net_),
            .in3(N__8122),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_7_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_7_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_1_7_1  (
            .in0(N__9377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8206),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_7_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_7_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_7_2  (
            .in0(_gnd_net_),
            .in1(N__8794),
            .in2(_gnd_net_),
            .in3(N__8123),
            .lcout(),
            .ltout(\uu0.un165_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_13_LC_1_7_3 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_7_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_7_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_13_LC_1_7_3  (
            .in0(N__8136),
            .in1(N__9137),
            .in2(N__8139),
            .in3(N__9223),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__9068),
            .sr(N__20677));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_7_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_7_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_1_7_4  (
            .in0(N__8230),
            .in1(N__9376),
            .in2(N__8208),
            .in3(N__8163),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_12_LC_1_7_5 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_7_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_7_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_12_LC_1_7_5  (
            .in0(N__8124),
            .in1(N__8795),
            .in2(N__8127),
            .in3(N__9222),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__9068),
            .sr(N__20677));
    defparam \uu0.l_count_6_LC_1_7_6 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_1_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_1_7_6 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_6_LC_1_7_6  (
            .in0(N__8207),
            .in1(N__9216),
            .in2(N__8235),
            .in3(N__9378),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__9068),
            .sr(N__20677));
    defparam \uu0.l_count_15_LC_1_7_7 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_7_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_7_7 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \uu0.l_count_15_LC_1_7_7  (
            .in0(N__8892),
            .in1(N__9138),
            .in2(N__9402),
            .in3(N__9224),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22244),
            .ce(N__9068),
            .sr(N__20677));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_8_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_1_8_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_1_8_0  (
            .in0(N__8717),
            .in1(N__8161),
            .in2(N__8259),
            .in3(N__8185),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_16_LC_1_8_1 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_1_8_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_1_8_1 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uu0.l_count_16_LC_1_8_1  (
            .in0(N__9214),
            .in1(N__9124),
            .in2(N__9051),
            .in3(N__8576),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.l_count_17_LC_1_8_2 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_1_8_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu0.l_count_17_LC_1_8_2  (
            .in0(N__8577),
            .in1(N__9045),
            .in2(N__9139),
            .in3(N__8187),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_8_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_1_8_3  (
            .in0(N__8186),
            .in1(N__9123),
            .in2(N__9050),
            .in3(N__8575),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_1_8_4 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_1_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_1_8_4 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uu0.l_count_18_LC_1_8_4  (
            .in0(_gnd_net_),
            .in1(N__9213),
            .in2(N__8175),
            .in3(N__9414),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.l_count_3_LC_1_8_5 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_8_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_8_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_3_LC_1_8_5  (
            .in0(N__8258),
            .in1(N__8148),
            .in2(N__8850),
            .in3(N__9219),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.l_count_9_LC_1_8_6 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_1_8_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu0.l_count_9_LC_1_8_6  (
            .in0(N__8718),
            .in1(_gnd_net_),
            .in2(N__9140),
            .in3(N__9093),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.l_count_7_LC_1_8_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_1_8_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_7_LC_1_8_7  (
            .in0(N__8162),
            .in1(N__8234),
            .in2(N__8172),
            .in3(N__9218),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22236),
            .ce(N__9067),
            .sr(N__20675));
    defparam \uu0.l_count_0_LC_1_9_0 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_9_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_9_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_9_0  (
            .in0(N__9000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9221),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(N__9066),
            .sr(N__20678));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_9_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_9_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_1_LC_1_9_1  (
            .in0(N__8909),
            .in1(N__8999),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.un44_ci ),
            .ltout(\uu0.un44_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_9_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \uu0.l_count_2_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8142),
            .in3(N__8845),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(N__9066),
            .sr(N__20678));
    defparam \uu0.l_count_1_LC_1_9_3 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_9_3 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \uu0.l_count_1_LC_1_9_3  (
            .in0(N__8910),
            .in1(N__9001),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(N__9066),
            .sr(N__20678));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_9_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_9_4  (
            .in0(N__8257),
            .in1(N__8844),
            .in2(N__9003),
            .in3(N__8908),
            .lcout(\uu0.un66_ci ),
            .ltout(\uu0.un66_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_4_LC_1_9_5 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_9_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uu0.l_count_4_LC_1_9_5  (
            .in0(_gnd_net_),
            .in1(N__9215),
            .in2(N__8238),
            .in3(N__8815),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(N__9066),
            .sr(N__20678));
    defparam \uu0.l_count_5_LC_1_9_6 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_1_9_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_1_9_6 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \uu0.l_count_5_LC_1_9_6  (
            .in0(N__8943),
            .in1(_gnd_net_),
            .in2(N__8820),
            .in3(N__8229),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(N__9066),
            .sr(N__20678));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_7 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(N__8814),
            .in2(_gnd_net_),
            .in3(N__8942),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_1_10_0 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_1_10_0 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_1_10_0 .LUT_INIT=16'b0100010100010000;
    LogicCell40 \resetGen.reset_count_1_LC_1_10_0  (
            .in0(N__11184),
            .in1(N__9441),
            .in2(N__9495),
            .in3(N__9510),
            .lcout(\resetGen.reset_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22224),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_1_10_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_1_10_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_1_10_1 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \resetGen.reset_count_0_LC_1_10_1  (
            .in0(N__9440),
            .in1(N__9491),
            .in2(_gnd_net_),
            .in3(N__11183),
            .lcout(\resetGen.reset_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22224),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_1_10_5 .C_ON=1'b0;
    defparam \resetGen.rst_LC_1_10_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_1_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9436),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22224),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_11_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_1_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__9719),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_11_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__8400),
            .in2(_gnd_net_),
            .in3(N__8190),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_11_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__9268),
            .in2(_gnd_net_),
            .in3(N__8325),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_11_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__8282),
            .in2(_gnd_net_),
            .in3(N__8322),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_1_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_11_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_1_11_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_1_11_4  (
            .in0(N__9540),
            .in1(N__9860),
            .in2(N__8313),
            .in3(N__8319),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22216),
            .ce(N__9653),
            .sr(N__20682));
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_1_12_0  (
            .in0(N__8308),
            .in1(N__9281),
            .in2(N__8283),
            .in3(N__8394),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOUCP_4_LC_1_12_1  (
            .in0(_gnd_net_),
            .in1(N__8307),
            .in2(_gnd_net_),
            .in3(N__9723),
            .lcout(),
            .ltout(\buart.Z_rx.valid_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_12_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_1_LC_1_12_2  (
            .in0(N__8277),
            .in1(N__9280),
            .in2(N__8316),
            .in3(N__8393),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_12_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIR1DP_4_LC_1_12_3  (
            .in0(_gnd_net_),
            .in1(N__8276),
            .in2(_gnd_net_),
            .in3(N__8309),
            .lcout(),
            .ltout(\buart.Z_rx.idle_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_12_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_1_12_4  (
            .in0(N__9724),
            .in1(N__9282),
            .in2(N__8292),
            .in3(N__8395),
            .lcout(\buart.Z_rx.idle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_1_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_12_6 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_1_12_6 .LUT_INIT=16'b0001110100101110;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_1_12_6  (
            .in0(N__8281),
            .in1(N__9541),
            .in2(N__9867),
            .in3(N__8289),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22209),
            .ce(N__9651),
            .sr(N__20685));
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_1_13_4 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_1_13_4  (
            .in0(N__9864),
            .in1(N__8409),
            .in2(N__9549),
            .in3(N__8399),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22202),
            .ce(N__9654),
            .sr(N__20687));
    defparam \uu2.r_data_reg_0_LC_2_1_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_2_1_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_0_LC_2_1_0  (
            .in0(N__8373),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_2_1_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_2_1_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_1_LC_2_1_1  (
            .in0(N__8367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_2_1_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_2_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_2_LC_2_1_2  (
            .in0(N__8361),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_2_1_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_2_1_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.r_data_reg_3_LC_2_1_3  (
            .in0(N__8355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_2_1_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_2_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8349),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_2_1_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_2_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_2_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8343),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_2_1_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_2_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_2_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8337),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_2_1_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_2_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_2_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8331),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__10680),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_2_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_2_2_0  (
            .in0(N__20418),
            .in1(N__8463),
            .in2(_gnd_net_),
            .in3(N__8499),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_2_2_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__8493),
            .in2(_gnd_net_),
            .in3(N__20424),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_2_2_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_2_2_2  (
            .in0(N__20417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8487),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_2_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_2_2_3  (
            .in0(N__8451),
            .in1(N__20421),
            .in2(_gnd_net_),
            .in3(N__8469),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_2_2_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_2_2_4  (
            .in0(N__20419),
            .in1(N__8439),
            .in2(_gnd_net_),
            .in3(N__8457),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_2_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_2_2_5  (
            .in0(N__8427),
            .in1(N__20422),
            .in2(_gnd_net_),
            .in3(N__8445),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_2_2_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_2_2_6  (
            .in0(N__20420),
            .in1(N__8415),
            .in2(_gnd_net_),
            .in3(N__8433),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_2_2_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_2_2_7  (
            .in0(N__10560),
            .in1(N__20423),
            .in2(_gnd_net_),
            .in3(N__8421),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22267),
            .ce(N__20376),
            .sr(N__20689));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_3_0 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_2_3_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(N__8514),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_2_3_4 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_2_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_2_3_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_2_3_4  (
            .in0(N__10169),
            .in1(N__8595),
            .in2(N__20438),
            .in3(N__20763),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22263),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_8_LC_2_4_1 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_2_4_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_2_4_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__8623),
            .in2(_gnd_net_),
            .in3(N__8508),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22258),
            .ce(),
            .sr(N__20658));
    defparam \uu2.vram_rd_clk_LC_2_4_2 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_2_4_2 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_2_4_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.vram_rd_clk_LC_2_4_2  (
            .in0(N__10168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8547),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22258),
            .ce(),
            .sr(N__20658));
    defparam \uu2.trig_rd_det_0_LC_2_4_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_2_4_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__10167),
            .in2(_gnd_net_),
            .in3(N__8594),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22258),
            .ce(),
            .sr(N__20658));
    defparam \uu2.trig_rd_det_1_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_2_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_2_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8526),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22258),
            .ce(),
            .sr(N__20658));
    defparam \uu0.l_precount_0_LC_2_4_6 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_2_4_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu0.l_precount_0_LC_2_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9339),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22258),
            .ce(),
            .sr(N__20658));
    defparam \uu2.l_count_5_LC_2_5_0 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_2_5_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_5_LC_2_5_0  (
            .in0(N__10391),
            .in1(N__8663),
            .in2(_gnd_net_),
            .in3(N__8643),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(N__20686));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_5_1  (
            .in0(N__10442),
            .in1(N__10371),
            .in2(N__10415),
            .in3(N__10388),
            .lcout(\uu2.un350_ci ),
            .ltout(\uu2.un350_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_2_5_2 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \uu2.l_count_9_LC_2_5_2  (
            .in0(N__8546),
            .in1(N__8624),
            .in2(N__8502),
            .in3(N__8681),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(N__20686));
    defparam \uu2.l_count_4_LC_2_5_3 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_2_5_3 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_2_5_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \uu2.l_count_4_LC_2_5_3  (
            .in0(N__8662),
            .in1(N__10390),
            .in2(_gnd_net_),
            .in3(N__8545),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(N__20686));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_4 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_2_5_4  (
            .in0(_gnd_net_),
            .in1(N__8661),
            .in2(_gnd_net_),
            .in3(N__8642),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(\uu2.vbuf_count.un328_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_6_LC_2_5_5 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_2_5_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_2_5_5 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \uu2.l_count_6_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__10441),
            .in2(N__8685),
            .in3(N__10389),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22252),
            .ce(),
            .sr(N__20686));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_2_5_6  (
            .in0(N__10439),
            .in1(N__8657),
            .in2(N__8682),
            .in3(N__10619),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_5_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_2_5_7  (
            .in0(N__10620),
            .in1(N__8680),
            .in2(N__8664),
            .in3(N__10440),
            .lcout(\uu2.un1_l_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_6_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_2_6_0  (
            .in0(N__10370),
            .in1(N__8641),
            .in2(N__8628),
            .in3(N__8884),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(\uu2.un1_l_count_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_6_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_2_6_1  (
            .in0(N__10328),
            .in1(N__8873),
            .in2(N__8604),
            .in3(N__8601),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_2_6_2  (
            .in0(N__9398),
            .in1(N__8748),
            .in2(N__8796),
            .in3(N__8771),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_2_6_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_2_6_3  (
            .in0(N__8870),
            .in1(N__8562),
            .in2(N__8556),
            .in3(N__10327),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_3_LC_2_6_4 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_2_6_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \uu2.l_count_3_LC_2_6_4  (
            .in0(N__10344),
            .in1(N__8871),
            .in2(N__8529),
            .in3(N__8886),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22245),
            .ce(),
            .sr(N__20684));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_6_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_6_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_2_6_5  (
            .in0(N__8772),
            .in1(N__8793),
            .in2(_gnd_net_),
            .in3(N__8749),
            .lcout(\uu0.un187_ci_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_6_6  (
            .in0(N__8872),
            .in1(N__10616),
            .in2(N__10329),
            .in3(N__8885),
            .lcout(\uu2.un306_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_2_6_7 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_2_6_7 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_2_6_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__10343),
            .in2(_gnd_net_),
            .in3(N__8874),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22245),
            .ce(),
            .sr(N__20684));
    defparam \uu0.l_count_RNI04591_10_LC_2_7_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI04591_10_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI04591_10_LC_2_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_count_RNI04591_10_LC_2_7_0  (
            .in0(N__8697),
            .in1(N__9088),
            .in2(N__8751),
            .in3(N__8846),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2GS72_4_LC_2_7_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2GS72_4_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2GS72_4_LC_2_7_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNI2GS72_4_LC_2_7_1  (
            .in0(N__9350),
            .in1(N__8769),
            .in2(N__8823),
            .in3(N__8819),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_10_LC_2_7_2 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_2_7_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_2_7_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_10_LC_2_7_2  (
            .in0(N__8700),
            .in1(N__9092),
            .in2(N__8724),
            .in3(N__9136),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22237),
            .ce(N__9069),
            .sr(N__20680));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_7_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_2_7_3  (
            .in0(N__9089),
            .in1(N__8719),
            .in2(N__9024),
            .in3(N__8698),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_2_7_4 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_2_7_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_2_7_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_count_14_LC_2_7_4  (
            .in0(N__8770),
            .in1(N__8750),
            .in2(N__8754),
            .in3(N__9135),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22237),
            .ce(N__9069),
            .sr(N__20680));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_7_5 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_7_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_2_7_5  (
            .in0(N__9090),
            .in1(N__8720),
            .in2(_gnd_net_),
            .in3(N__8699),
            .lcout(),
            .ltout(\uu0.un143_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_11_LC_2_7_6 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_2_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_2_7_6 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_11_LC_2_7_6  (
            .in0(N__9023),
            .in1(N__9134),
            .in2(N__9144),
            .in3(N__9217),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22237),
            .ce(N__9069),
            .sr(N__20680));
    defparam \uu0.l_count_8_LC_2_7_7 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_2_7_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu0.l_count_8_LC_2_7_7  (
            .in0(N__9091),
            .in1(_gnd_net_),
            .in2(N__9141),
            .in3(_gnd_net_),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22237),
            .ce(N__9069),
            .sr(N__20680));
    defparam \uu0.delay_line_0_LC_2_8_0 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_2_8_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_2_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_2_8_0  (
            .in0(N__8956),
            .in1(N__9312),
            .in2(N__8928),
            .in3(N__9351),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(),
            .sr(N__20676));
    defparam \uu0.l_count_RNI2CNU_11_LC_2_8_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2CNU_11_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2CNU_11_LC_2_8_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uu0.l_count_RNI2CNU_11_LC_2_8_1  (
            .in0(N__9049),
            .in1(N__9019),
            .in2(N__9002),
            .in3(N__8955),
            .lcout(),
            .ltout(\uu0.un4_l_count_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_8_2 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_11_LC_2_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_11_LC_2_8_2  (
            .in0(N__8976),
            .in1(N__8970),
            .in2(N__8964),
            .in3(N__9360),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_precount_2_LC_2_8_4 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_2_8_4 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \uu0.l_precount_2_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__9313),
            .in2(N__8961),
            .in3(N__9352),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(),
            .sr(N__20676));
    defparam \uu0.l_precount_3_LC_2_8_5 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_2_8_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_2_8_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_2_8_5  (
            .in0(N__9353),
            .in1(N__8926),
            .in2(N__9318),
            .in3(N__8960),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(),
            .sr(N__20676));
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_8_6 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_2_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_2_8_6  (
            .in0(N__9311),
            .in1(N__8941),
            .in2(N__8927),
            .in3(N__8907),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI96A32_18_LC_2_8_7 .C_ON=1'b0;
    defparam \uu0.l_count_RNI96A32_18_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI96A32_18_LC_2_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI96A32_18_LC_2_8_7  (
            .in0(N__9413),
            .in1(N__9397),
            .in2(N__9381),
            .in3(N__9375),
            .lcout(\uu0.un4_l_count_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_1_LC_2_9_0 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_2_9_0 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_2_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9239),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22225),
            .ce(),
            .sr(N__20681));
    defparam \buart.Z_rx.hh_1_LC_2_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_2_9_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_2_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9566),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22225),
            .ce(),
            .sr(N__20681));
    defparam \uu0.l_precount_1_LC_2_9_3 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_2_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_2_9_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.l_precount_1_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__9354),
            .in2(_gnd_net_),
            .in3(N__9317),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22225),
            .ce(),
            .sr(N__20681));
    defparam \uu0.sec_clk_LC_2_9_6 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_2_9_6 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_2_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__17512),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22225),
            .ce(),
            .sr(N__20681));
    defparam CONSTANT_ONE_LUT4_LC_2_10_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_10_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_10_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(CONSTANT_ONE_NET_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_2_10_1 .LUT_INIT=16'b0011001101011010;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_2_10_1  (
            .in0(N__9726),
            .in1(N__9859),
            .in2(N__9291),
            .in3(N__9536),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22217),
            .ce(N__9652),
            .sr(N__20683));
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_2_10_2 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_2_10_2  (
            .in0(N__9858),
            .in1(N__9288),
            .in2(N__9545),
            .in3(N__9279),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22217),
            .ce(N__9652),
            .sr(N__20683));
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_2_10_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_2_10_6  (
            .in0(N__9249),
            .in1(N__9240),
            .in2(_gnd_net_),
            .in3(N__9225),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_2_10_7  (
            .in0(N__16245),
            .in1(N__12111),
            .in2(_gnd_net_),
            .in3(N__21772),
            .lcout(\uu2.mem0.w_addr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_2_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_2_11_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_2_11_0  (
            .in0(N__13016),
            .in1(N__9567),
            .in2(_gnd_net_),
            .in3(N__9667),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_2_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_2_11_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_2_11_1  (
            .in0(N__9668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14961),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_11_2 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_2__un241_ci_LC_2_11_2  (
            .in0(N__9508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9489),
            .lcout(\resetGen.un241_ci ),
            .ltout(\resetGen.un241_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_2_11_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_2_11_3 .LUT_INIT=16'b0000000010011010;
    LogicCell40 \resetGen.reset_count_2_LC_2_11_3  (
            .in0(N__9462),
            .in1(N__9438),
            .in2(N__9513),
            .in3(N__11175),
            .lcout(\resetGen.reset_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22210),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_4 .C_ON=1'b0;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \resetGen.uu0.counter_gen_label_3__un252_ci_LC_2_11_4  (
            .in0(N__9509),
            .in1(N__9490),
            .in2(_gnd_net_),
            .in3(N__9461),
            .lcout(),
            .ltout(\resetGen.un252_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_2_11_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_2_11_5 .LUT_INIT=16'b0000000010011010;
    LogicCell40 \resetGen.reset_count_3_LC_2_11_5  (
            .in0(N__9471),
            .in1(N__9439),
            .in2(N__9474),
            .in3(N__11176),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22210),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_RNO_0_4_LC_2_11_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \resetGen.reset_count_RNO_0_4_LC_2_11_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \resetGen.reset_count_RNO_0_4_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__9470),
            .in2(_gnd_net_),
            .in3(N__9460),
            .lcout(),
            .ltout(\resetGen.reset_count_2_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_2_11_7 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_2_11_7 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \resetGen.reset_count_4_LC_2_11_7  (
            .in0(N__9450),
            .in1(N__9437),
            .in2(N__9444),
            .in3(N__11177),
            .lcout(\resetGen.reset_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22210),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_2_12_0  (
            .in0(N__9735),
            .in1(N__9882),
            .in2(_gnd_net_),
            .in3(N__9725),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__9847),
            .in2(_gnd_net_),
            .in3(N__9598),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_2_12_2  (
            .in0(N__9910),
            .in1(N__9933),
            .in2(N__9800),
            .in3(N__9619),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__9958),
            .in2(N__9678),
            .in3(N__9597),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_2_12_4  (
            .in0(N__9846),
            .in1(N__9942),
            .in2(N__9675),
            .in3(N__9960),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_5 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_5 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_2_12_5  (
            .in0(N__9884),
            .in1(N__9848),
            .in2(N__9915),
            .in3(N__9894),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_2_12_6  (
            .in0(N__9845),
            .in1(_gnd_net_),
            .in2(N__9605),
            .in3(N__9620),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22203),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_2_12_7  (
            .in0(N__9883),
            .in1(N__9844),
            .in2(N__9672),
            .in3(N__14962),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(N__9621),
            .in2(N__9606),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_13_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_2_13_1  (
            .in0(_gnd_net_),
            .in1(N__9959),
            .in2(_gnd_net_),
            .in3(N__9936),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_2_13_2  (
            .in0(N__9866),
            .in1(N__9932),
            .in2(_gnd_net_),
            .in3(N__9918),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__22197),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(N__9911),
            .in2(_gnd_net_),
            .in3(N__9888),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_2_13_4  (
            .in0(N__9885),
            .in1(N__9865),
            .in2(N__9801),
            .in3(N__9804),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22197),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_4_1_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_4_1_0  (
            .in0(N__10274),
            .in1(N__10243),
            .in2(N__9758),
            .in3(N__10214),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__10182),
            .sr(N__20674));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_4_1_1  (
            .in0(_gnd_net_),
            .in1(N__10477),
            .in2(_gnd_net_),
            .in3(N__10113),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_4_1_2 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_8_LC_4_1_2  (
            .in0(N__9776),
            .in1(N__10005),
            .in2(N__9783),
            .in3(N__10068),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__10182),
            .sr(N__20674));
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_4_1_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_4_1_3  (
            .in0(N__10069),
            .in1(N__10046),
            .in2(N__10028),
            .in3(N__9765),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__10182),
            .sr(N__20674));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_4_1_4  (
            .in0(N__10273),
            .in1(N__10242),
            .in2(N__9757),
            .in3(N__10213),
            .lcout(\uu2.un404_ci_0 ),
            .ltout(\uu2.un404_ci_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_4_1_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.r_addr_esr_6_LC_4_1_5  (
            .in0(N__10024),
            .in1(N__10478),
            .in2(N__10053),
            .in3(N__10114),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22264),
            .ce(N__10182),
            .sr(N__20674));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_6 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_4_1_6  (
            .in0(_gnd_net_),
            .in1(N__10045),
            .in2(_gnd_net_),
            .in3(N__10020),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_7_LC_4_1_7  (
            .in0(N__13197),
            .in1(N__13304),
            .in2(N__13431),
            .in3(N__13384),
            .lcout(\uu2.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0 .LUT_INIT=16'b1011101000010000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_4_2_0  (
            .in0(N__21766),
            .in1(N__12993),
            .in2(N__11319),
            .in3(N__11127),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_4_2_1  (
            .in0(N__9987),
            .in1(N__10965),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(\uu2.mem0.w_data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uu2.w_addr_displaying_RNI4E8U4_8_LC_4_2_2  (
            .in0(N__11291),
            .in1(N__11311),
            .in2(_gnd_net_),
            .in3(N__12991),
            .lcout(\uu2.N_34 ),
            .ltout(\uu2.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3 .LUT_INIT=16'b1011101110111000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_4_2_3  (
            .in0(N__10905),
            .in1(N__21768),
            .in2(N__9981),
            .in3(N__10700),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_4_2_4  (
            .in0(N__10701),
            .in1(N__10293),
            .in2(N__21787),
            .in3(N__11022),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_4_2_5  (
            .in0(N__10292),
            .in1(N__10842),
            .in2(_gnd_net_),
            .in3(N__21764),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6 .LUT_INIT=16'b0010001000110010;
    LogicCell40 \uu2.w_addr_displaying_RNIQN495_0_LC_4_2_6  (
            .in0(N__11292),
            .in1(N__12992),
            .in2(N__11318),
            .in3(N__12107),
            .lcout(\uu2.N_31 ),
            .ltout(\uu2.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(N__21767),
            .in2(N__10284),
            .in3(N__10884),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_2_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_4_3_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_2_LC_4_3_0  (
            .in0(N__10142),
            .in1(N__10269),
            .in2(N__10247),
            .in3(N__10209),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22253),
            .ce(),
            .sr(N__20668));
    defparam \uu2.r_addr_1_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_4_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_4_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uu2.r_addr_1_LC_4_3_1  (
            .in0(N__10208),
            .in1(N__10238),
            .in2(_gnd_net_),
            .in3(N__10140),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22253),
            .ce(),
            .sr(N__20668));
    defparam \uu2.r_addr_0_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_4_3_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.r_addr_0_LC_4_3_2  (
            .in0(N__10139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10207),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22253),
            .ce(),
            .sr(N__20668));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__10138),
            .in2(_gnd_net_),
            .in3(N__20761),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_4_LC_4_3_7 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_4_3_7 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_4_3_7  (
            .in0(N__10106),
            .in1(N__10076),
            .in2(_gnd_net_),
            .in3(N__10141),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22253),
            .ce(),
            .sr(N__20668));
    defparam \uu2.vram_rd_clk_det_0_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_4_4_0 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_4_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10170),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.vram_rd_clk_det_0C_net ),
            .ce(),
            .sr(N__20629));
    defparam \uu2.r_addr_5_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_4_5_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_5_LC_4_5_0  (
            .in0(N__10146),
            .in1(N__10115),
            .in2(N__10476),
            .in3(N__10080),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22238),
            .ce(),
            .sr(N__20661));
    defparam \uu2.l_count_7_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_4_5_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_4_5_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.l_count_7_LC_4_5_1  (
            .in0(N__10446),
            .in1(N__10363),
            .in2(N__10419),
            .in3(N__10398),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22238),
            .ce(),
            .sr(N__20661));
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_4_5_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_4_5_2  (
            .in0(N__11436),
            .in1(_gnd_net_),
            .in2(N__12279),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22238),
            .ce(),
            .sr(N__20661));
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_4_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__12275),
            .in2(_gnd_net_),
            .in3(N__11435),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22238),
            .ce(),
            .sr(N__20661));
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_ctle_3_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__14811),
            .in2(_gnd_net_),
            .in3(N__20754),
            .lcout(\Lab_UT.didp.regrce3.LdAMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_5_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_5_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__10311),
            .in2(_gnd_net_),
            .in3(N__10617),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_1_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_4_5_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_4_5_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.l_count_1_LC_4_5_6  (
            .in0(N__10618),
            .in1(_gnd_net_),
            .in2(N__10323),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22238),
            .ce(),
            .sr(N__20661));
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_4_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_4_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_0_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20050),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(N__10986),
            .sr(N__20659));
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_4_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_4_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_1_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21390),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(N__10986),
            .sr(N__20659));
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_4_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_4_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_2_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20956),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(N__10986),
            .sr(N__20659));
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_4_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_4_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_3_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21140),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22231),
            .ce(N__10986),
            .sr(N__20659));
    defparam \uu2.vram_wr_en_0_i_LC_4_7_7 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_4_7_7 .LUT_INIT=16'b0010111110101111;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_4_7_7  (
            .in0(N__10796),
            .in1(N__10943),
            .in2(N__22281),
            .in3(N__10863),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_8_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_8_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_4_8_2  (
            .in0(N__14293),
            .in1(N__20046),
            .in2(_gnd_net_),
            .in3(N__14361),
            .lcout(\Lab_UT.didp.countrce1.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_0 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_3_LC_4_9_0 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \Lab_UT.alarmchar_latch_3_LC_4_9_0  (
            .in0(N__11048),
            .in1(N__10497),
            .in2(N__11096),
            .in3(N__10488),
            .lcout(G_188),
            .ltout(G_188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_4_9_1 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_4_9_1  (
            .in0(N__18119),
            .in1(N__11587),
            .in2(N__10491),
            .in3(N__11460),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_4_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_4_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_4_9_2 .LUT_INIT=16'b0000010101000101;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_4_9_2  (
            .in0(N__10821),
            .in1(N__10658),
            .in2(N__11592),
            .in3(N__18121),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22211),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_9_4 .C_ON=1'b0;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_4_9_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.un1_armed_2_0_iso_i_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__11693),
            .in2(_gnd_net_),
            .in3(N__11646),
            .lcout(\Lab_UT.un1_armed_2_0_iso_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_rst_0_iclk_LC_4_9_5 .C_ON=1'b0;
    defparam \Lab_UT.un1_rst_0_iclk_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_rst_0_iclk_LC_4_9_5 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \Lab_UT.un1_rst_0_iclk_LC_4_9_5  (
            .in0(N__20749),
            .in1(_gnd_net_),
            .in2(N__11708),
            .in3(N__11647),
            .lcout(\Lab_UT.un1_rst_0_iclkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_4_9_6 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_4_9_6  (
            .in0(N__10820),
            .in1(N__10657),
            .in2(N__11591),
            .in3(N__18120),
            .lcout(\Lab_UT.dispString.dOutP_1_iv_i_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m1_LC_4_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m1_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m1_LC_4_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.m1_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(N__11701),
            .in2(_gnd_net_),
            .in3(N__11650),
            .lcout(G_182),
            .ltout(G_182_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_4_LC_4_10_1 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_4_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_4_LC_4_10_1 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \Lab_UT.alarmchar_latch_4_LC_4_10_1  (
            .in0(N__11702),
            .in1(N__20755),
            .in2(N__10662),
            .in3(N__10659),
            .lcout(G_187),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_4_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_4_10_2 .LUT_INIT=16'b0001000000110011;
    LogicCell40 \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_LC_4_10_2  (
            .in0(N__10641),
            .in1(N__11495),
            .in2(N__11769),
            .in3(N__10629),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.justentered_latch_LC_4_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.justentered_latch_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.justentered_latch_LC_4_10_3 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \Lab_UT.dictrl.justentered_latch_LC_4_10_3  (
            .in0(N__11494),
            .in1(N__10639),
            .in2(N__10644),
            .in3(N__20756),
            .lcout(G_183),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_4_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_4_10_6 .LUT_INIT=16'b1111111110001100;
    LogicCell40 \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_4_10_6  (
            .in0(N__10640),
            .in1(N__10628),
            .in2(N__11768),
            .in3(N__11493),
            .lcout(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_0_LC_4_11_7 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_4_11_7 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_4_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uu2.l_count_0_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10599),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22198),
            .ce(),
            .sr(N__20688));
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_5_1_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_5_1_0  (
            .in0(N__20451),
            .in1(N__10539),
            .in2(_gnd_net_),
            .in3(N__10572),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22259),
            .ce(N__20372),
            .sr(N__20693));
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_5_1_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(N__20452),
            .in2(_gnd_net_),
            .in3(N__10548),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22259),
            .ce(N__20372),
            .sr(N__20693));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_5_1_2  (
            .in0(N__15978),
            .in1(N__21748),
            .in2(_gnd_net_),
            .in3(N__13262),
            .lcout(\uu2.mem0.w_addr_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_5_1_3  (
            .in0(N__10734),
            .in1(N__10719),
            .in2(_gnd_net_),
            .in3(N__20747),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4 .LUT_INIT=16'b0001000110001000;
    LogicCell40 \uu2.w_addr_displaying_RNI03P31_4_LC_5_1_4  (
            .in0(N__21692),
            .in1(N__20273),
            .in2(_gnd_net_),
            .in3(N__13383),
            .lcout(\uu2.w_addr_displaying_RNI03P31Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \uu2.w_addr_user_RNI93NG7_4_LC_5_1_5  (
            .in0(N__16260),
            .in1(N__10797),
            .in2(_gnd_net_),
            .in3(N__10809),
            .lcout(\uu2.un28_w_addr_user_i ),
            .ltout(\uu2.un28_w_addr_user_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNID65PE_4_LC_5_1_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_user_RNID65PE_4_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10671),
            .in3(N__15929),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNI43E87_4_LC_5_1_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \uu2.w_addr_user_RNI43E87_4_LC_5_1_7  (
            .in0(N__16259),
            .in1(N__20746),
            .in2(_gnd_net_),
            .in3(N__10808),
            .lcout(\uu2.w_addr_user_RNI43E87Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_5_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_5_2_0 .LUT_INIT=16'b0010000111011110;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI1BE61_2_LC_5_2_0  (
            .in0(N__16554),
            .in1(N__13386),
            .in2(N__13789),
            .in3(N__12137),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_m24_0_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_5_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_5_2_1 .LUT_INIT=16'b0000100101000010;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIDDQM2_3_LC_5_2_1  (
            .in0(N__12106),
            .in1(N__16106),
            .in2(N__10668),
            .in3(N__11279),
            .lcout(\uu2.bitmap_pmux_sn_i5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_5_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_5_2_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI6DFN_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__11388),
            .in2(_gnd_net_),
            .in3(N__13385),
            .lcout(\uu2.bitmap_pmux_sn_N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_5_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_5_2_3 .LUT_INIT=16'b0001001100010010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNISF1A1_2_LC_5_2_3  (
            .in0(N__12138),
            .in1(N__16623),
            .in2(N__11397),
            .in3(N__13782),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_N_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_5_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_5_2_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNINCTH4_2_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__13743),
            .in2(N__10665),
            .in3(N__11952),
            .lcout(\uu2.N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_5_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_LC_5_2_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_LC_5_2_5  (
            .in0(N__11392),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16555),
            .lcout(\uu2.w_addr_displaying_1_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__11901),
            .sr(N__20617));
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_5_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_1_LC_5_2_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_1_LC_5_2_6  (
            .in0(N__16556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11393),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__11901),
            .sr(N__20617));
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_1_LC_5_2_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_1_LC_5_2_7  (
            .in0(N__11394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16557),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_1_rep1_nesrC_net ),
            .ce(N__11901),
            .sr(N__20617));
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNINQUSG_2_LC_5_3_0  (
            .in0(N__10686),
            .in1(N__10740),
            .in2(_gnd_net_),
            .in3(N__10710),
            .lcout(),
            .ltout(\uu2.N_406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \uu2.w_addr_displaying_RNI6SEI31_8_LC_5_3_1  (
            .in0(N__11256),
            .in1(N__10764),
            .in2(N__10704),
            .in3(N__11325),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNIO4T61_LC_5_3_2  (
            .in0(N__13777),
            .in1(N__13263),
            .in2(_gnd_net_),
            .in3(N__11395),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNICM7R_180_LC_5_3_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNICM7R_180_LC_5_3_3  (
            .in0(N__16371),
            .in1(N__12243),
            .in2(_gnd_net_),
            .in3(N__11936),
            .lcout(),
            .ltout(\uu2.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_RNI2UBA2_LC_5_3_4  (
            .in0(N__13778),
            .in1(N__16631),
            .in2(N__10692),
            .in3(N__12219),
            .lcout(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2 ),
            .ltout(\uu2.w_addr_displaying_3_rep1_nesr_RNI2UBAZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \uu2.w_addr_displaying_RNI0NG56_0_4_LC_5_3_5  (
            .in0(N__12005),
            .in1(N__10757),
            .in2(N__10689),
            .in3(N__16313),
            .lcout(\uu2.w_addr_displaying_RNI0NG56_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \uu2.w_addr_displaying_RNI8GJC3_8_LC_5_3_6  (
            .in0(N__13264),
            .in1(N__10770),
            .in2(_gnd_net_),
            .in3(N__16632),
            .lcout(\uu2.bitmap_pmux_u_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7 .LUT_INIT=16'b1101111110001111;
    LogicCell40 \uu2.w_addr_displaying_RNI0NG56_4_LC_5_3_7  (
            .in0(N__10758),
            .in1(N__16314),
            .in2(N__12009),
            .in3(N__10746),
            .lcout(\uu2.w_addr_displaying_RNI0NG56Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_1_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_5_4_5 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_5_4_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__10733),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.vram_rd_clk_det_1C_net ),
            .ce(),
            .sr(N__20630));
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_5_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_0_LC_5_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_0_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20052),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22232),
            .ce(N__14621),
            .sr(N__20664));
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_5_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_2_LC_5_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_2_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20945),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22232),
            .ce(N__14621),
            .sr(N__20664));
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_5_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_3_LC_5_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_3_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21121),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22232),
            .ce(N__14621),
            .sr(N__20664));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_6_0 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_5_6_0  (
            .in0(N__18002),
            .in1(N__17123),
            .in2(N__11523),
            .in3(N__13612),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_1_LC_5_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_5_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_5_6_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_5_6_3  (
            .in0(N__18080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18201),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22226),
            .ce(),
            .sr(N__20662));
    defparam \Lab_UT.dispString.cnt_0_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_5_6_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_5_6_4 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_5_6_4  (
            .in0(N__18003),
            .in1(N__17492),
            .in2(N__18220),
            .in3(N__18081),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22226),
            .ce(),
            .sr(N__20662));
    defparam \Lab_UT.didp.ce_0_LC_5_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_5_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_5_6_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_5_6_5  (
            .in0(N__17491),
            .in1(N__12687),
            .in2(_gnd_net_),
            .in3(N__18478),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22226),
            .ce(),
            .sr(N__20662));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_6 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_6  (
            .in0(N__14420),
            .in1(N__12173),
            .in2(N__14546),
            .in3(N__17122),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_7 .LUT_INIT=16'b1111000011111100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__12564),
            .in2(N__10812),
            .in3(N__14680),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_5_7_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_7_LC_5_7_0  (
            .in0(N__17294),
            .in1(N__13579),
            .in2(N__17087),
            .in3(N__12517),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_0_LC_5_7_1 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_0_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_0_LC_5_7_1 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \uu2.un4_w_user_data_rdy_0_LC_5_7_1  (
            .in0(N__10862),
            .in1(_gnd_net_),
            .in2(N__10944),
            .in3(N__10792),
            .lcout(\uu2.un4_w_user_data_rdyZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un20_w_addr_user_1_LC_5_7_2 .C_ON=1'b0;
    defparam \uu2.un20_w_addr_user_1_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.un20_w_addr_user_1_LC_5_7_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \uu2.un20_w_addr_user_1_LC_5_7_2  (
            .in0(N__10911),
            .in1(N__10939),
            .in2(N__10974),
            .in3(N__10861),
            .lcout(\uu2.un20_w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_5_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_5_7_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dispString.rdy_LC_5_7_4  (
            .in0(N__18197),
            .in1(N__18007),
            .in2(N__17493),
            .in3(N__18079),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22218),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_5_7_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_5_7_5  (
            .in0(N__18078),
            .in1(N__18196),
            .in2(_gnd_net_),
            .in3(N__11148),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_5_7_6 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_5_7_6  (
            .in0(N__14547),
            .in1(N__12495),
            .in2(N__10776),
            .in3(N__12401),
            .lcout(),
            .ltout(\Lab_UT.dispString.dOutP_0_iv_i_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_5_7_7 .LUT_INIT=16'b0000010100000100;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_5_7_7  (
            .in0(N__17429),
            .in1(N__11552),
            .in2(N__10773),
            .in3(N__13650),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22218),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_5_8_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_5_8_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_5_8_0  (
            .in0(N__19137),
            .in1(N__18477),
            .in2(N__20766),
            .in3(N__19511),
            .lcout(\Lab_UT.didp.regrce4.LdAMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_4_LC_5_8_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.un1_w_user_lf_4_LC_5_8_1  (
            .in0(N__10877),
            .in1(N__10835),
            .in2(N__10964),
            .in3(N__11012),
            .lcout(\uu2.un1_w_user_lfZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_8_2 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_5_8_2  (
            .in0(N__18115),
            .in1(N__11146),
            .in2(N__17430),
            .in3(N__11581),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_4_LC_5_8_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.un1_w_user_cr_4_LC_5_8_3  (
            .in0(N__10957),
            .in1(N__21869),
            .in2(N__11123),
            .in3(N__11011),
            .lcout(\uu2.un1_w_user_crZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_5_8_4 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_5_8_4  (
            .in0(N__11551),
            .in1(N__10926),
            .in2(N__13686),
            .in3(N__10917),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22212),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_lf_3_LC_5_8_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uu2.un1_w_user_lf_3_LC_5_8_5  (
            .in0(N__10898),
            .in1(N__11116),
            .in2(_gnd_net_),
            .in3(N__21868),
            .lcout(\uu2.un1_w_user_lfZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_3_LC_5_8_6 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_3_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_3_LC_5_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \uu2.un1_w_user_cr_3_LC_5_8_6  (
            .in0(N__10834),
            .in1(N__10897),
            .in2(_gnd_net_),
            .in3(N__10876),
            .lcout(\uu2.un1_w_user_crZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_5_8_7 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_5_8_7  (
            .in0(N__18012),
            .in1(N__18116),
            .in2(_gnd_net_),
            .in3(N__10848),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22212),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_5_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_1_LC_5_9_0 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIKUO21_1_LC_5_9_0  (
            .in0(N__18226),
            .in1(N__17542),
            .in2(N__17571),
            .in3(N__12542),
            .lcout(\Lab_UT.dispString.cnt_RNIKUO21Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_1 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_0_LC_5_9_1 .LUT_INIT=16'b1111110101010101;
    LogicCell40 \Lab_UT.alarmchar_latch_0_LC_5_9_1  (
            .in0(N__11651),
            .in1(N__11147),
            .in2(N__20765),
            .in3(N__11703),
            .lcout(G_186),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_5_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_5_9_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_5_9_3  (
            .in0(N__18123),
            .in1(N__11583),
            .in2(_gnd_net_),
            .in3(N__11198),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22204),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_idle_4_0_iclk_LC_5_9_4 .C_ON=1'b0;
    defparam \Lab_UT.un1_idle_4_0_iclk_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_idle_4_0_iclk_LC_5_9_4 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \Lab_UT.un1_idle_4_0_iclk_LC_5_9_4  (
            .in0(N__11704),
            .in1(N__11652),
            .in2(_gnd_net_),
            .in3(N__11215),
            .lcout(),
            .ltout(\Lab_UT.un1_idle_4_0_iclkZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_1_LC_5_9_5 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_1_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_1_LC_5_9_5 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.alarmchar_latch_1_LC_5_9_5  (
            .in0(N__11094),
            .in1(N__11049),
            .in2(N__11037),
            .in3(N__11034),
            .lcout(G_185),
            .ltout(G_185_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_5_9_6  (
            .in0(_gnd_net_),
            .in1(N__11582),
            .in2(N__11028),
            .in3(N__18122),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_117_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_5_9_7 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_5_9_7  (
            .in0(N__11544),
            .in1(N__11409),
            .in2(N__11025),
            .in3(N__17831),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22204),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_5_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_5_10_0 .LUT_INIT=16'b1011101111111111;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_5_10_0  (
            .in0(N__20764),
            .in1(N__11699),
            .in2(_gnd_net_),
            .in3(N__11654),
            .lcout(G_180),
            .ltout(G_180_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_5_10_1 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_1_LC_5_10_1  (
            .in0(N__11700),
            .in1(N__10998),
            .in2(N__10992),
            .in3(N__11217),
            .lcout(G_181),
            .ltout(G_181_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_5_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_5_10_2 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_0__m3_LC_5_10_2  (
            .in0(N__11496),
            .in1(N__11653),
            .in2(N__10989),
            .in3(N__11753),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_5_10_3 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_0_LC_5_10_3  (
            .in0(N__11655),
            .in1(N__11226),
            .in2(N__11220),
            .in3(N__11216),
            .lcout(G_179),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m59_LC_5_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m59_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m59_LC_5_10_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.m59_LC_5_10_6  (
            .in0(N__11648),
            .in1(N__14910),
            .in2(_gnd_net_),
            .in3(N__11697),
            .lcout(\Lab_UT.alarmstate_0_sqmuxa_1 ),
            .ltout(\Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_6_LC_5_10_7 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_6_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_6_LC_5_10_7 .LUT_INIT=16'b0000111000000110;
    LogicCell40 \Lab_UT.alarmchar_latch_6_LC_5_10_7  (
            .in0(N__11698),
            .in1(N__11649),
            .in2(N__11202),
            .in3(N__11199),
            .lcout(G_184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m37_LC_5_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m37_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m37_LC_5_12_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m37_LC_5_12_1  (
            .in0(N__12906),
            .in1(N__13091),
            .in2(N__11742),
            .in3(N__12811),
            .lcout(\Lab_UT.dictrl.next_state6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_5_LC_5_12_3 .C_ON=1'b0;
    defparam \resetGen.escKey_5_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_5_LC_5_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \resetGen.escKey_5_LC_5_12_3  (
            .in0(N__13093),
            .in1(N__15747),
            .in2(N__20928),
            .in3(N__12812),
            .lcout(),
            .ltout(\resetGen.escKeyZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_LC_5_12_4 .C_ON=1'b0;
    defparam \resetGen.escKey_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_LC_5_12_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \resetGen.escKey_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__11154),
            .in2(N__11187),
            .in3(N__14974),
            .lcout(\resetGen.escKeyZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.escKey_4_LC_5_12_5 .C_ON=1'b0;
    defparam \resetGen.escKey_4_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \resetGen.escKey_4_LC_5_12_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \resetGen.escKey_4_LC_5_12_5  (
            .in0(N__21313),
            .in1(N__19990),
            .in2(N__15610),
            .in3(N__21097),
            .lcout(\resetGen.escKeyZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_0_LC_5_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_0_LC_5_12_6 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g2_0_LC_5_12_6  (
            .in0(N__21096),
            .in1(N__21312),
            .in2(_gnd_net_),
            .in3(N__20904),
            .lcout(\Lab_UT.dictrl.g2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_5_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_5_LC_5_12_7 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_5_LC_5_12_7  (
            .in0(N__13092),
            .in1(N__15746),
            .in2(N__18479),
            .in3(N__15596),
            .lcout(\Lab_UT.dictrl.G_25_i_o3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_0_LC_5_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_5_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_5_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21306),
            .lcout(bu_rx_data_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22193),
            .ce(N__20794),
            .sr(N__20690));
    defparam \buart.Z_rx.shifter_1_LC_5_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_5_14_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_1_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20900),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22193),
            .ce(N__20794),
            .sr(N__20690));
    defparam \buart.Z_rx.shifter_3_LC_5_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_5_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_5_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15602),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22193),
            .ce(N__20794),
            .sr(N__20690));
    defparam \buart.Z_rx.shifter_7_LC_5_15_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_5_15_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_5_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13028),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22190),
            .ce(N__20792),
            .sr(N__20692));
    defparam \uu2.w_addr_user_2_LC_6_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_2_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_2_LC_6_1_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_2_LC_6_1_0  (
            .in0(N__21836),
            .in1(N__16231),
            .in2(N__20341),
            .in3(N__11245),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_user_1_LC_6_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_6_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_6_1_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \uu2.w_addr_user_1_LC_6_1_1  (
            .in0(N__11243),
            .in1(_gnd_net_),
            .in2(N__16238),
            .in3(N__20332),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_user_0_LC_6_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_0_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_0_LC_6_1_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_user_0_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(N__16227),
            .in2(_gnd_net_),
            .in3(N__11242),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_user_4_LC_6_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_6_1_3 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.w_addr_user_4_LC_6_1_3  (
            .in0(N__11244),
            .in1(N__16012),
            .in2(_gnd_net_),
            .in3(N__16294),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_user_5_LC_6_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_5_LC_6_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_5_LC_6_1_4 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_5_LC_6_1_4  (
            .in0(N__16295),
            .in1(N__15521),
            .in2(N__16017),
            .in3(N__11246),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_user_6_LC_6_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_6_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_6_LC_6_1_5 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_6_LC_6_1_5  (
            .in0(N__11247),
            .in1(N__16016),
            .in2(N__16039),
            .in3(N__16193),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_2C_net ),
            .ce(),
            .sr(N__15941));
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_displaying_RNI47N27_8_LC_6_1_6  (
            .in0(_gnd_net_),
            .in1(N__20748),
            .in2(_gnd_net_),
            .in3(N__15879),
            .lcout(\uu2.N_33_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_6_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_6_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIKIPH1_8_LC_6_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIKIPH1_8_LC_6_2_0  (
            .in0(N__20275),
            .in1(N__21676),
            .in2(N__16121),
            .in3(N__13266),
            .lcout(\uu2.un51_w_data_displaying_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_6_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_6_2_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4JSO_1_LC_6_2_1  (
            .in0(_gnd_net_),
            .in1(N__12079),
            .in2(_gnd_net_),
            .in3(N__20274),
            .lcout(),
            .ltout(\uu2.w_data_displaying_2_i_a2_i_a3_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_6_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_6_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIASLS1_8_LC_6_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIASLS1_8_LC_6_2_2  (
            .in0(N__21675),
            .in1(N__16113),
            .in2(N__11295),
            .in3(N__13265),
            .lcout(\uu2.w_data_displaying_2_i_a2_i_a3_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_3_LC_6_2_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_3_LC_6_2_3  (
            .in0(N__16114),
            .in1(N__20278),
            .in2(N__21688),
            .in3(N__12084),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__11890),
            .sr(N__20620));
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_6_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_3_LC_6_2_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_3_LC_6_2_4  (
            .in0(N__20276),
            .in1(N__21678),
            .in2(N__12099),
            .in3(N__11937),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__11890),
            .sr(N__20620));
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_6_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_6_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_nesr_LC_6_2_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_nesr_LC_6_2_5  (
            .in0(N__21677),
            .in1(N__20277),
            .in2(N__13790),
            .in3(N__12080),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_3C_net ),
            .ce(N__11890),
            .sr(N__20620));
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_6_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_6_2_6 .LUT_INIT=16'b1100110001001000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIO7503_3_LC_6_2_6  (
            .in0(N__21674),
            .in1(N__13161),
            .in2(N__16120),
            .in3(N__11280),
            .lcout(),
            .ltout(\uu2.w_addr_displaying_nesr_RNIO7503Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_6_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0FGN6_4_LC_6_2_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_RNI0FGN6_4_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(N__11268),
            .in2(N__11259),
            .in3(N__12015),
            .lcout(\uu2.bitmap_pmux_sn_i7_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_93_LC_6_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_6_3_0 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_93_LC_6_3_0  (
            .in0(N__16482),
            .in1(N__16451),
            .in2(N__17724),
            .in3(N__16920),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__20618));
    defparam \uu2.bitmap_221_LC_6_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_6_3_1 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_221_LC_6_3_1  (
            .in0(N__16919),
            .in1(N__17720),
            .in2(N__16452),
            .in3(N__16481),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_93C_net ),
            .ce(),
            .sr(N__20618));
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_6_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_6_3_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_1_rep1_nesr_RNI0TIL_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__16542),
            .in2(_gnd_net_),
            .in3(N__11396),
            .lcout(\uu2.N_31_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIPIHG1_75_LC_6_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPIHG1_75_LC_6_3_3 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.bitmap_RNIPIHG1_75_LC_6_3_3  (
            .in0(N__16543),
            .in1(N__11991),
            .in2(N__11985),
            .in3(N__14001),
            .lcout(),
            .ltout(\uu2.N_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_6_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_6_3_4 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI4IVU3_3_LC_6_3_4  (
            .in0(N__16116),
            .in1(N__11345),
            .in2(N__11364),
            .in3(N__12192),
            .lcout(\uu2.bitmap_pmux_27_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI6MCU1_93_LC_6_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI6MCU1_93_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI6MCU1_93_LC_6_3_5 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.bitmap_RNI6MCU1_93_LC_6_3_5  (
            .in0(N__16544),
            .in1(N__11361),
            .in2(N__11355),
            .in3(N__16491),
            .lcout(),
            .ltout(\uu2.N_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI72CH8_69_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI72CH8_69_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI72CH8_69_LC_6_3_6 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \uu2.bitmap_RNI72CH8_69_LC_6_3_6  (
            .in0(N__11346),
            .in1(N__11907),
            .in2(N__11334),
            .in3(N__11331),
            .lcout(\uu2.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_3_LC_6_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_6_5_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_6_5_0  (
            .in0(N__12273),
            .in1(N__14186),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__20669));
    defparam \Lab_UT.didp.ce_1_LC_6_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_6_5_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_6_5_1  (
            .in0(N__12185),
            .in1(N__17884),
            .in2(N__17496),
            .in3(N__13726),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__20669));
    defparam \Lab_UT.didp.reset_0_LC_6_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_6_5_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_6_5_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_6_5_2  (
            .in0(N__13727),
            .in1(N__17487),
            .in2(N__17891),
            .in3(N__12186),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__20669));
    defparam \Lab_UT.didp.reset_2_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_6_5_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_6_5_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_6_5_4  (
            .in0(N__12274),
            .in1(N__14187),
            .in2(_gnd_net_),
            .in3(N__11429),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__20669));
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_5_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNIULOK1_3_LC_6_5_5  (
            .in0(N__12184),
            .in1(N__17883),
            .in2(N__17495),
            .in3(N__13725),
            .lcout(\Lab_UT.didp.ce_12_1 ),
            .ltout(\Lab_UT.didp.ce_12_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_5_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__12262),
            .in2(N__11415),
            .in3(N__14185),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_6_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_6_5_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_6_5_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_6_5_7  (
            .in0(N__16758),
            .in1(N__17619),
            .in2(N__11412),
            .in3(N__13508),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22222),
            .ce(),
            .sr(N__20669));
    defparam \Lab_UT.didp.countrce2.q_3_LC_6_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_6_6_0 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_6_6_0  (
            .in0(N__12482),
            .in1(N__12327),
            .in2(N__12465),
            .in3(N__12305),
            .lcout(\Lab_UT.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22215),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_6_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_6_6_1 .LUT_INIT=16'b0000000010001011;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_6_6_1  (
            .in0(N__13854),
            .in1(N__12483),
            .in2(N__12321),
            .in3(N__12459),
            .lcout(\Lab_UT.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22215),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_6_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_6_6_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_6_LC_6_6_2  (
            .in0(N__16749),
            .in1(N__12397),
            .in2(N__12626),
            .in3(N__12169),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_6_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_6_6_3 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_2_LC_6_6_3  (
            .in0(N__13853),
            .in1(N__12364),
            .in2(N__12309),
            .in3(N__14579),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_6_6_4 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_6_6_4  (
            .in0(N__14559),
            .in1(N__12559),
            .in2(N__17494),
            .in3(N__14519),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_6_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_6_6_5  (
            .in0(N__17877),
            .in1(N__14346),
            .in2(_gnd_net_),
            .in3(N__16989),
            .lcout(\Lab_UT.didp.countrce1.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_6_6_7 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_6_6_7  (
            .in0(N__18194),
            .in1(N__18077),
            .in2(N__18008),
            .in3(N__12365),
            .lcout(\Lab_UT.dispString.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_7_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_LC_6_7_1  (
            .in0(N__13491),
            .in1(N__13675),
            .in2(N__13721),
            .in3(N__13534),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_6_7_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_13_LC_6_7_2  (
            .in0(N__12336),
            .in1(N__14172),
            .in2(N__11514),
            .in3(N__11511),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_6_7_3  (
            .in0(N__11505),
            .in1(N__12408),
            .in2(N__11499),
            .in3(N__11442),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_7_5 .LUT_INIT=16'b1101111000010010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_6_7_5  (
            .in0(N__13709),
            .in1(N__14292),
            .in2(N__11472),
            .in3(N__21116),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_6_7_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_6_7_6  (
            .in0(N__14251),
            .in1(N__14210),
            .in2(N__11463),
            .in3(N__13710),
            .lcout(\Lab_UT.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22208),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_3_LC_6_7_7 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_3_LC_6_7_7  (
            .in0(N__18195),
            .in1(N__12558),
            .in2(N__17480),
            .in3(N__13535),
            .lcout(\Lab_UT.dispString.N_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_2 .LUT_INIT=16'b1001000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_12_LC_6_8_2  (
            .in0(N__13631),
            .in1(N__14336),
            .in2(N__11601),
            .in3(N__11448),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_6_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_6_8_3 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_6_8_3  (
            .in0(N__17679),
            .in1(N__21117),
            .in2(N__12153),
            .in3(N__13497),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_6_8_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_6_8_4  (
            .in0(N__13498),
            .in1(N__16831),
            .in2(N__11730),
            .in3(N__16788),
            .lcout(\Lab_UT.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_6_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_6_8_5 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_6_8_5  (
            .in0(N__11727),
            .in1(N__16942),
            .in2(N__11553),
            .in3(N__11718),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_8_6 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_6_8_6  (
            .in0(N__17677),
            .in1(N__20031),
            .in2(_gnd_net_),
            .in3(N__17083),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_6_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_6_8_7 .LUT_INIT=16'b0101000001000001;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_6_8_7  (
            .in0(N__16830),
            .in1(N__16808),
            .in2(N__11712),
            .in3(N__17678),
            .lcout(\Lab_UT.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22201),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_9_1 .LUT_INIT=16'b0000100100000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_0_LC_6_9_1  (
            .in0(N__13619),
            .in1(N__16707),
            .in2(N__11709),
            .in3(N__11645),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_6_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIH15E_2_LC_6_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIH15E_2_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__17982),
            .in2(_gnd_net_),
            .in3(N__18228),
            .lcout(\Lab_UT.dispString.un42_dOutP_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_6_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_6_9_4 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \Lab_UT.dispString.cnt_RNIOG7L_2_LC_6_9_4  (
            .in0(N__18114),
            .in1(N__17997),
            .in2(_gnd_net_),
            .in3(N__18227),
            .lcout(\Lab_UT.dispString.N_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dispString.cnt_RNIG05E_2_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(N__17981),
            .in2(_gnd_net_),
            .in3(N__18113),
            .lcout(\Lab_UT.dispString.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_6_9_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_ctle_3_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(N__14844),
            .in2(_gnd_net_),
            .in3(N__20762),
            .lcout(\Lab_UT.didp.regrce2.LdAStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_10_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_0_LC_6_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_0_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20032),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22196),
            .ce(N__11778),
            .sr(N__20665));
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_10_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_1_LC_6_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_1_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21352),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22196),
            .ce(N__11778),
            .sr(N__20665));
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_10_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_2_LC_6_10_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_2_LC_6_10_2  (
            .in0(N__20957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22196),
            .ce(N__11778),
            .sr(N__20665));
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_10_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_esr_3_LC_6_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_3_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21094),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22196),
            .ce(N__11778),
            .sr(N__20665));
    defparam \Lab_UT.dictrl.alarmstate8_LC_6_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_LC_6_11_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_LC_6_11_0  (
            .in0(N__13103),
            .in1(N__15741),
            .in2(N__19036),
            .in3(N__11784),
            .lcout(\Lab_UT.dictrl.alarmstateZ0Z8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_5_LC_6_11_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_5_LC_6_11_1  (
            .in0(N__15743),
            .in1(N__12823),
            .in2(N__19774),
            .in3(N__15609),
            .lcout(\Lab_UT.dictrl.g1_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m37_N_2L1_LC_6_11_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m37_N_2L1_LC_6_11_2  (
            .in0(N__20006),
            .in1(N__15742),
            .in2(N__20927),
            .in3(N__21231),
            .lcout(\Lab_UT.dictrl.m37_N_2LZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_1_LC_6_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_1_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_1_LC_6_11_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_1_LC_6_11_4  (
            .in0(N__12824),
            .in1(N__21092),
            .in2(N__13112),
            .in3(N__15744),
            .lcout(\Lab_UT.dictrl.g0_5_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_1_LC_6_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_1_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_1_LC_6_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \Lab_UT.dictrl.g1_0_1_LC_6_11_5  (
            .in0(N__21232),
            .in1(N__13104),
            .in2(_gnd_net_),
            .in3(N__19696),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_6_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_6_11_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNII6R92_LC_6_11_6  (
            .in0(N__17239),
            .in1(N__11814),
            .in2(N__11808),
            .in3(N__21336),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_6_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_6_11_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIR0L55_1_LC_6_11_7  (
            .in0(N__11805),
            .in1(N__11793),
            .in2(N__11799),
            .in3(N__19923),
            .lcout(\Lab_UT.dictrl.N_55_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_6_1_LC_6_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.g0_6_1_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__15745),
            .in2(_gnd_net_),
            .in3(N__12807),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_6Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIC4II1_0_LC_6_12_2  (
            .in0(N__19510),
            .in1(N__15587),
            .in2(N__11796),
            .in3(N__13101),
            .lcout(\Lab_UT.dictrl.g0_6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_12_3 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNITL791_0_LC_6_12_3  (
            .in0(N__20908),
            .in1(N__19509),
            .in2(N__15603),
            .in3(N__21314),
            .lcout(\Lab_UT.dictrl.g0_5_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_12_4 .LUT_INIT=16'b1010111111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_9_LC_6_12_4  (
            .in0(N__12808),
            .in1(_gnd_net_),
            .in2(N__19929),
            .in3(N__20139),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_25_i_o3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_12_5 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_6_LC_6_12_5  (
            .in0(N__21054),
            .in1(N__21315),
            .in2(N__11787),
            .in3(N__20909),
            .lcout(\Lab_UT.dictrl.G_25_i_o3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_6_12_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_3_LC_6_12_7  (
            .in0(N__15583),
            .in1(N__12806),
            .in2(N__21213),
            .in3(N__19668),
            .lcout(\Lab_UT.dictrl.alarmstate8Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_6_13_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_6_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_LC_6_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21307),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_6_LC_6_13_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_6_13_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_6_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_LC_6_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13102),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_fast_4_LC_6_13_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_6_13_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_6_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_6_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15739),
            .lcout(buart__rx_shifter_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_0_rep1_LC_6_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_LC_6_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_rep1_LC_6_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_LC_6_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21308),
            .lcout(bu_rx_data_0_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_fast_2_LC_6_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_6_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_6_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21044),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_3_rep2_LC_6_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_LC_6_13_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep2_LC_6_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15600),
            .lcout(bu_rx_data_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_4_LC_6_13_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_6_13_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_6_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_6_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15738),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22192),
            .ce(N__20795),
            .sr(N__20691));
    defparam \buart.Z_rx.shifter_2_rep1_LC_6_14_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_6_14_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_6_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21084),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22189),
            .ce(N__20793),
            .sr(N__20694));
    defparam \buart.Z_rx.shifter_5_rep1_LC_6_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_rep1_LC_6_14_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_rep1_LC_6_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_5_rep1_LC_6_14_5  (
            .in0(N__12822),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_5_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22189),
            .ce(N__20793),
            .sr(N__20694));
    defparam \buart.Z_rx.shifter_fast_5_LC_6_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_6_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12821),
            .lcout(bu_rx_data_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22189),
            .ce(N__20793),
            .sr(N__20694));
    defparam \buart.Z_rx.shifter_fast_3_LC_6_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_6_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_6_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15601),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22189),
            .ce(N__20793),
            .sr(N__20694));
    defparam \buart.Z_rx.shifter_5_LC_6_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_6_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_6_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_5_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12825),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22188),
            .ce(N__20790),
            .sr(N__20695));
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_7_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_7_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_7_1_0 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI6VOF1_6_LC_7_1_0  (
            .in0(N__16633),
            .in1(N__13296),
            .in2(N__13193),
            .in3(N__13369),
            .lcout(\uu2.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_6_LC_7_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_7_1_1 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_7_1_1 .LUT_INIT=16'b1100101111000011;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_7_1_1  (
            .in0(N__13249),
            .in1(N__13189),
            .in2(N__13323),
            .in3(N__16635),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_ness_6C_net ),
            .ce(N__11897),
            .sr(N__20624));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_2 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_7_1_2  (
            .in0(N__13188),
            .in1(_gnd_net_),
            .in2(N__21803),
            .in3(N__16181),
            .lcout(\uu2.mem0.w_addr_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_1_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_7_1_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_7_1_3  (
            .in0(N__13370),
            .in1(N__16289),
            .in2(_gnd_net_),
            .in3(N__21788),
            .lcout(\uu2.mem0.w_addr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_4 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_7_1_4  (
            .in0(N__21789),
            .in1(N__15519),
            .in2(_gnd_net_),
            .in3(N__13297),
            .lcout(\uu2.mem0.w_addr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_1_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_1_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_6__un426_ci_3_LC_7_1_5  (
            .in0(N__15520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16290),
            .lcout(\uu2.un426_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_7_1_6  (
            .in0(N__16634),
            .in1(_gnd_net_),
            .in2(N__21804),
            .in3(N__16160),
            .lcout(\uu2.mem0.w_addr_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_1_7 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_1_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_8__un448_ci_0_LC_7_1_7  (
            .in0(N__16161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16191),
            .lcout(\uu2.vbuf_w_addr_user.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_168_LC_7_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_7_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_7_2_0 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_168_LC_7_2_0  (
            .in0(N__13908),
            .in1(N__14151),
            .in2(N__13946),
            .in3(N__13974),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__20623));
    defparam \uu2.bitmap_40_LC_7_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_7_2_1 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_40_LC_7_2_1  (
            .in0(N__13976),
            .in1(N__13941),
            .in2(N__14160),
            .in3(N__13910),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__20623));
    defparam \uu2.bitmap_75_LC_7_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_7_2_2 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.bitmap_75_LC_7_2_2  (
            .in0(N__13911),
            .in1(N__14158),
            .in2(N__13947),
            .in3(N__13977),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__20623));
    defparam \uu2.bitmap_203_LC_7_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_7_2_3 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \uu2.bitmap_203_LC_7_2_3  (
            .in0(N__13975),
            .in1(N__13940),
            .in2(N__14159),
            .in3(N__13909),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__20623));
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJS4P_162_LC_7_2_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIJS4P_162_LC_7_2_4  (
            .in0(N__11933),
            .in1(N__11976),
            .in2(_gnd_net_),
            .in3(N__13131),
            .lcout(\uu2.N_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_5 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_RNIT3TB_1_LC_7_2_5  (
            .in0(N__12127),
            .in1(N__11970),
            .in2(_gnd_net_),
            .in3(N__11935),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_sn_N_54_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \uu2.bitmap_RNI2Q8F1_111_LC_7_2_6  (
            .in0(_gnd_net_),
            .in1(N__16647),
            .in2(N__11961),
            .in3(N__11958),
            .lcout(\uu2.bitmap_RNI2Q8F1Z0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIBPBO_40_LC_7_2_7 .LUT_INIT=16'b0000011111000111;
    LogicCell40 \uu2.bitmap_RNIBPBO_40_LC_7_2_7  (
            .in0(N__11943),
            .in1(N__11934),
            .in2(N__16353),
            .in3(N__13881),
            .lcout(\uu2.bitmap_pmux_26_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_197_LC_7_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_7_3_0 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \uu2.bitmap_197_LC_7_3_0  (
            .in0(N__13563),
            .in1(N__14664),
            .in2(N__13473),
            .in3(N__14490),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20621));
    defparam \uu2.bitmap_RNITSCU1_69_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNITSCU1_69_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNITSCU1_69_LC_7_3_1 .LUT_INIT=16'b1101010110000101;
    LogicCell40 \uu2.bitmap_RNITSCU1_69_LC_7_3_1  (
            .in0(N__13137),
            .in1(N__11913),
            .in2(N__12093),
            .in3(N__13734),
            .lcout(\uu2.N_166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_0_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_7_3_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__12072),
            .in2(_gnd_net_),
            .in3(N__15889),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20621));
    defparam \uu2.w_addr_displaying_fast_2_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_7_3_3 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_7_3_3  (
            .in0(N__15891),
            .in1(N__20297),
            .in2(N__12095),
            .in3(N__12131),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20621));
    defparam \uu2.w_addr_displaying_2_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_7_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_7_3_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_displaying_2_LC_7_3_4  (
            .in0(N__20296),
            .in1(N__15890),
            .in2(N__12092),
            .in3(N__21673),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_197C_net ),
            .ce(),
            .sr(N__20621));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_7_3_5 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_4_LC_7_3_5  (
            .in0(N__21672),
            .in1(N__16099),
            .in2(N__12094),
            .in3(N__20295),
            .lcout(\uu2.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_7_3_6 .LUT_INIT=16'b1000000100000000;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI84IJ2_3_LC_7_3_6  (
            .in0(N__16098),
            .in1(N__21671),
            .in2(N__12091),
            .in3(N__13314),
            .lcout(\uu2.w_addr_displaying_nesr_RNI84IJ2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIGEPH1_4_LC_7_3_7 .LUT_INIT=16'b0110101000001000;
    LogicCell40 \uu2.w_addr_displaying_RNIGEPH1_4_LC_7_3_7  (
            .in0(N__21670),
            .in1(N__20294),
            .in2(N__16115),
            .in3(N__13382),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_7_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_7_4_0 .LUT_INIT=16'b0000011100011001;
    LogicCell40 \uu2.bitmap_308_LC_7_4_0  (
            .in0(N__14060),
            .in1(N__14388),
            .in2(N__14111),
            .in3(N__13830),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_212_LC_7_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_7_4_1 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_212_LC_7_4_1  (
            .in0(N__14387),
            .in1(N__13829),
            .in2(N__14110),
            .in3(N__14059),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_84_LC_7_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_7_4_2 .LUT_INIT=16'b0000010000111101;
    LogicCell40 \uu2.bitmap_84_LC_7_4_2  (
            .in0(N__14062),
            .in1(N__14390),
            .in2(N__14113),
            .in3(N__13832),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_180_LC_7_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_7_4_3 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_180_LC_7_4_3  (
            .in0(N__14386),
            .in1(N__13828),
            .in2(N__14109),
            .in3(N__14058),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_52_LC_7_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_7_4_4 .LUT_INIT=16'b1101111101111001;
    LogicCell40 \uu2.bitmap_52_LC_7_4_4  (
            .in0(N__14061),
            .in1(N__14389),
            .in2(N__14112),
            .in3(N__13831),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIB3QK_52_LC_7_4_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIB3QK_52_LC_7_4_5  (
            .in0(N__16349),
            .in1(N__12231),
            .in2(_gnd_net_),
            .in3(N__12225),
            .lcout(\uu2.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_87_LC_7_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_7_4_6 .LUT_INIT=16'b0001101110110111;
    LogicCell40 \uu2.bitmap_87_LC_7_4_6  (
            .in0(N__14063),
            .in1(N__14391),
            .in2(N__14114),
            .in3(N__13833),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__20619));
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIRMQA1_84_LC_7_4_7 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \uu2.bitmap_RNIRMQA1_84_LC_7_4_7  (
            .in0(N__12207),
            .in1(N__16407),
            .in2(N__12201),
            .in3(N__14025),
            .lcout(\uu2.N_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI19F76_0_LC_7_5_0  (
            .in0(N__17790),
            .in1(N__17301),
            .in2(_gnd_net_),
            .in3(N__12518),
            .lcout(\Lab_UT.min2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_7_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_7_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_7_5_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNI0JJJ_2_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(N__14355),
            .in2(_gnd_net_),
            .in3(N__16979),
            .lcout(\Lab_UT.didp.countrce1.ce_12_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_7_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_7_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI5DF76_2_LC_7_5_2  (
            .in0(N__17791),
            .in1(N__16747),
            .in2(_gnd_net_),
            .in3(N__12174),
            .lcout(\Lab_UT.min2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_5_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_5_3  (
            .in0(N__17037),
            .in1(N__17618),
            .in2(_gnd_net_),
            .in3(N__17101),
            .lcout(\Lab_UT.didp.countrce4.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_7_5_5 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_2_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12627),
            .in3(N__13865),
            .lcout(\Lab_UT.didp.countrce2.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNIVQ0O5_0_LC_7_5_6  (
            .in0(N__17792),
            .in1(N__12620),
            .in2(_gnd_net_),
            .in3(N__12402),
            .lcout(\Lab_UT.sec1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI511O5_3_LC_7_5_7  (
            .in0(N__12372),
            .in1(N__12306),
            .in2(_gnd_net_),
            .in3(N__17793),
            .lcout(\Lab_UT.sec1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_6_0 .LUT_INIT=16'b1011011110000100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_7_6_0  (
            .in0(N__14454),
            .in1(N__12655),
            .in2(N__12345),
            .in3(N__20946),
            .lcout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_7_6_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_4_LC_7_6_1  (
            .in0(N__17029),
            .in1(N__16943),
            .in2(N__16985),
            .in3(N__14515),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_6_2 .LUT_INIT=16'b0101111111111111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_3_LC_7_6_2  (
            .in0(N__14453),
            .in1(_gnd_net_),
            .in2(N__12625),
            .in3(N__13870),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.N_96_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_3 .LUT_INIT=16'b1101011110000010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_7_6_3  (
            .in0(N__12656),
            .in1(N__12308),
            .in2(N__12330),
            .in3(N__21136),
            .lcout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_4 .LUT_INIT=16'b1001100100001111;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_1_LC_7_6_4  (
            .in0(N__12615),
            .in1(N__13871),
            .in2(N__21391),
            .in3(N__12657),
            .lcout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIAE4B1_LC_7_6_5  (
            .in0(N__18473),
            .in1(N__19922),
            .in2(N__17252),
            .in3(N__18346),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_6_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_7_6_6  (
            .in0(N__14452),
            .in1(N__12307),
            .in2(N__12624),
            .in3(N__13869),
            .lcout(\Lab_UT.didp.un24_ce_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_7 .LUT_INIT=16'b0011000010111010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_7_6_7  (
            .in0(N__17124),
            .in1(N__13589),
            .in2(N__12563),
            .in3(N__12522),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI62AM_1_LC_7_7_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI62AM_1_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__12431),
            .in2(_gnd_net_),
            .in3(N__12646),
            .lcout(\Lab_UT.didp.un1_dicLdStens_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdStens_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_7_7_1 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_7_7_1  (
            .in0(N__14439),
            .in1(N__12474),
            .in2(N__12468),
            .in3(N__12464),
            .lcout(\Lab_UT.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22219),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_7_7_2 .LUT_INIT=16'b0000010101000001;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_7_7_2  (
            .in0(N__12463),
            .in1(N__12647),
            .in2(N__12579),
            .in3(N__12432),
            .lcout(\Lab_UT.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22219),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_7_7_3 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_7_7_3  (
            .in0(N__14208),
            .in1(N__12420),
            .in2(N__14258),
            .in3(N__14351),
            .lcout(\Lab_UT.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22219),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_7_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__17036),
            .in2(_gnd_net_),
            .in3(N__17077),
            .lcout(\Lab_UT.didp.countrce4.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_7_5 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_5_LC_7_7_5  (
            .in0(N__17865),
            .in1(N__14410),
            .in2(N__14450),
            .in3(N__17827),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_7_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_7_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__20757),
            .in2(_gnd_net_),
            .in3(N__18246),
            .lcout(\Lab_UT.didp.regrce1.LdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_7_7_7 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_7_7_7  (
            .in0(N__17866),
            .in1(N__14209),
            .in2(N__14259),
            .in3(N__12570),
            .lcout(\Lab_UT.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22219),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_10_esr_LC_7_8_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_10_esr_LC_7_8_0  (
            .in0(N__15069),
            .in1(N__18603),
            .in2(N__15224),
            .in3(N__15029),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(N__18514),
            .sr(N__20660));
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_7_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_11_ess_LC_7_8_1 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_ess_LC_7_8_1  (
            .in0(N__15030),
            .in1(N__15220),
            .in2(N__18611),
            .in3(N__15070),
            .lcout(\Lab_UT.LdSones_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(N__18514),
            .sr(N__20660));
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_7_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_7_8_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_7_8_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_LC_7_8_2  (
            .in0(N__15071),
            .in1(N__18607),
            .in2(N__15225),
            .in3(N__15031),
            .lcout(\Lab_UT.state_ret_8_ess ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(N__18514),
            .sr(N__20660));
    defparam \Lab_UT.didp.state_ret_1_esr_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.state_ret_1_esr_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.state_ret_1_esr_LC_7_8_3 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \Lab_UT.didp.state_ret_1_esr_LC_7_8_3  (
            .in0(N__15032),
            .in1(_gnd_net_),
            .in2(N__18612),
            .in3(N__15072),
            .lcout(\Lab_UT.didp.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22213),
            .ce(N__18514),
            .sr(N__20660));
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIFQ9K_0_LC_7_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.didp.ce_RNIFQ9K_0_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__12675),
            .in2(_gnd_net_),
            .in3(N__12669),
            .lcout(\Lab_UT.didp.un1_dicLdSones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_7_8_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_0_LC_7_8_6  (
            .in0(N__12645),
            .in1(N__20030),
            .in2(_gnd_net_),
            .in3(N__12616),
            .lcout(\Lab_UT.didp.countrce2.q_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_8_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_7_8_7  (
            .in0(N__21377),
            .in1(N__14347),
            .in2(N__14294),
            .in3(N__17881),
            .lcout(\Lab_UT.didp.countrce1.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_1_LC_7_9_1  (
            .in0(N__21378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22205),
            .ce(N__12705),
            .sr(N__20666));
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_2_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20958),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22205),
            .ce(N__12705),
            .sr(N__20666));
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_3_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21141),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22205),
            .ce(N__12705),
            .sr(N__20666));
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_7_9_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_7_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_7_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_0_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20033),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22205),
            .ce(N__12705),
            .sr(N__20666));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_10_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m21_LC_7_10_0  (
            .in0(N__18987),
            .in1(N__15494),
            .in2(N__17248),
            .in3(N__19865),
            .lcout(\Lab_UT.dictrl.N_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_2_LC_7_10_1  (
            .in0(N__19227),
            .in1(N__14978),
            .in2(N__14919),
            .in3(N__18628),
            .lcout(\Lab_UT.dictrl.G_25_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_4_LC_7_10_2 .LUT_INIT=16'b0001101111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_4_LC_7_10_2  (
            .in0(N__18339),
            .in1(N__15774),
            .in2(N__12918),
            .in3(N__18441),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_25_i_a5_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_3 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_1_LC_7_10_3  (
            .in0(N__19228),
            .in1(N__14724),
            .in2(N__12693),
            .in3(N__14979),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_25_i_a5_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_13_LC_7_10_4 .LUT_INIT=16'b0100010100000101;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_LC_7_10_4  (
            .in0(N__12729),
            .in1(N__18590),
            .in2(N__12690),
            .in3(N__15073),
            .lcout(\Lab_UT.un1_next_state66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22199),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_7_10_5 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNIK3GV_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(N__19581),
            .in2(N__19256),
            .in3(N__19120),
            .lcout(\Lab_UT.dictrl.G_14_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIH8JQ_2_LC_7_10_6  (
            .in0(N__18340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19596),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIH8JQZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g2_LC_7_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g2_LC_7_10_7  (
            .in0(_gnd_net_),
            .in1(N__18708),
            .in2(_gnd_net_),
            .in3(N__18338),
            .lcout(\Lab_UT.dictrl.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_11_0 .LUT_INIT=16'b0101110011111100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_mb_LC_7_11_0  (
            .in0(N__15264),
            .in1(N__12744),
            .in2(N__12762),
            .in3(N__12939),
            .lcout(),
            .ltout(\Lab_UT.i8_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_11_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_2_1_LC_7_11_1 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \Lab_UT.didp.g0_0_2_1_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__12750),
            .in2(N__12765),
            .in3(N__18341),
            .lcout(\Lab_UT.didp.g0_0_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_sn_LC_7_11_2  (
            .in0(N__18550),
            .in1(N__21229),
            .in2(N__17247),
            .in3(N__19695),
            .lcout(\Lab_UT.dictrl.g0_0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_11_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_1_0_LC_7_11_3  (
            .in0(N__19886),
            .in1(_gnd_net_),
            .in2(N__18469),
            .in3(N__20135),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_11_4 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g1_LC_7_11_4  (
            .in0(N__21481),
            .in1(N__19029),
            .in2(N__12753),
            .in3(N__21230),
            .lcout(\Lab_UT.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_11_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_rn_LC_7_11_5  (
            .in0(N__19600),
            .in1(N__17231),
            .in2(_gnd_net_),
            .in3(N__18549),
            .lcout(\Lab_UT.dictrl.g0_0_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_11_7 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_0_LC_7_11_7  (
            .in0(N__12738),
            .in1(N__14996),
            .in2(N__19281),
            .in3(N__12834),
            .lcout(\Lab_UT.dictrl.G_25_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_12_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNISV3C5_1_LC_7_12_0  (
            .in0(N__19919),
            .in1(N__12723),
            .in2(N__12714),
            .in3(N__12924),
            .lcout(\Lab_UT.dictrl.N_57_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_1_LC_7_12_1 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_1_LC_7_12_1  (
            .in0(N__20183),
            .in1(N__19400),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.m13_out ),
            .ltout(\Lab_UT.dictrl.m13_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_12_2 .LUT_INIT=16'b1000000010001000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_LC_7_12_2  (
            .in0(N__21468),
            .in1(N__20152),
            .in2(N__12858),
            .in3(N__21212),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_18_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_12_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_4_LC_7_12_3  (
            .in0(N__17243),
            .in1(N__12954),
            .in2(N__12855),
            .in3(N__19918),
            .lcout(\Lab_UT.dictrl.N_22_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKTFH_LC_7_12_5  (
            .in0(N__19985),
            .in1(_gnd_net_),
            .in2(N__20157),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.g1_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_12_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_7_LC_7_12_6  (
            .in0(N__17238),
            .in1(N__19607),
            .in2(N__18561),
            .in3(N__15681),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_13_RNOZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_12_7 .LUT_INIT=16'b1110111000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_3_LC_7_12_7  (
            .in0(N__12852),
            .in1(N__12846),
            .in2(N__12837),
            .in3(N__18348),
            .lcout(\Lab_UT.dictrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m34_1_LC_7_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m34_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m34_1_LC_7_13_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m34_1_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__15398),
            .in2(_gnd_net_),
            .in3(N__19401),
            .lcout(\Lab_UT.dictrl.m34Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.m34Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m34_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m34_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m34_LC_7_13_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m34_LC_7_13_2  (
            .in0(N__12810),
            .in1(N__13111),
            .in2(N__12828),
            .in3(N__15737),
            .lcout(\Lab_UT.dictrl.N_67_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_7_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_7_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_7_LC_7_13_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.g1_7_LC_7_13_3  (
            .in0(N__15736),
            .in1(N__12809),
            .in2(N__13113),
            .in3(N__15589),
            .lcout(\Lab_UT.dictrl.g1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_1_LC_7_13_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.m22_1_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__19740),
            .in2(_gnd_net_),
            .in3(N__19359),
            .lcout(\Lab_UT.dictrl.m22Z0Z_1 ),
            .ltout(\Lab_UT.dictrl.m22Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_8_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_8_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_8_LC_7_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_8_LC_7_13_5  (
            .in0(N__19989),
            .in1(N__15262),
            .in2(N__12957),
            .in3(N__21223),
            .lcout(\Lab_UT.dictrl.N_72_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJ5AG2_LC_7_13_6  (
            .in0(N__15263),
            .in1(N__21104),
            .in2(N__12948),
            .in3(N__12938),
            .lcout(\Lab_UT.dictrl.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_4_LC_7_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_4_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_4_LC_7_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.m22_4_LC_7_14_0  (
            .in0(N__15665),
            .in1(N__15367),
            .in2(N__15645),
            .in3(N__15399),
            .lcout(\Lab_UT.dictrl.m22Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_7_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_8_LC_7_14_1 .LUT_INIT=16'b0101111100110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_8_LC_7_14_1  (
            .in0(N__15351),
            .in1(N__15320),
            .in2(N__15342),
            .in3(N__19921),
            .lcout(\Lab_UT.dictrl.g1_rn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_7_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_7_14_2 .LUT_INIT=16'b0111000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI61IM_0_LC_7_14_2  (
            .in0(N__19739),
            .in1(N__19347),
            .in2(N__15439),
            .in3(N__15588),
            .lcout(\Lab_UT.dictrl.g0_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m5_LC_7_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m5_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m5_LC_7_14_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.m5_LC_7_14_3  (
            .in0(N__15400),
            .in1(N__13001),
            .in2(N__15376),
            .in3(N__15827),
            .lcout(N_63_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_0_x1_LC_7_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_0_x1_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_0_x1_LC_7_14_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.g1_0_x1_LC_7_14_4  (
            .in0(N__15641),
            .in1(N__12899),
            .in2(N__12887),
            .in3(N__12869),
            .lcout(\Lab_UT.dictrl.g1_0_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_1_5_LC_7_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_5_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_5_LC_7_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.g1_1_5_LC_7_14_5  (
            .in0(N__15401),
            .in1(N__15815),
            .in2(N__12888),
            .in3(N__20192),
            .lcout(\Lab_UT.dictrl.g1_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_7_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_7_14_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI43D01_0_LC_7_14_6  (
            .in0(N__13002),
            .in1(_gnd_net_),
            .in2(N__15440),
            .in3(N__12870),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_7_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_7_14_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI9GK03_0_LC_7_14_7  (
            .in0(N__19348),
            .in1(N__15666),
            .in2(N__13125),
            .in3(N__13122),
            .lcout(\Lab_UT.dictrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_rep1_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_6_rep1_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13099),
            .lcout(bu_rx_data_6_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22191),
            .ce(N__20789),
            .sr(N__20696));
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_15_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_15_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13034),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22191),
            .ce(N__20789),
            .sr(N__20696));
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_7_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_7_15_5  (
            .in0(N__13100),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22191),
            .ce(N__20789),
            .sr(N__20696));
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_7_15_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_7_15_6  (
            .in0(N__13035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22191),
            .ce(N__20789),
            .sr(N__20696));
    defparam \uu2.w_addr_displaying_fast_8_LC_8_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_8_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_8_LC_8_1_0 .LUT_INIT=16'b1111000010110100;
    LogicCell40 \uu2.w_addr_displaying_fast_8_LC_8_1_0  (
            .in0(N__12982),
            .in1(N__15878),
            .in2(N__16348),
            .in3(N__13422),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20627));
    defparam \uu2.w_addr_displaying_8_LC_8_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_8_1_1 .LUT_INIT=16'b1111110100000010;
    LogicCell40 \uu2.w_addr_displaying_8_LC_8_1_1  (
            .in0(N__15877),
            .in1(N__12981),
            .in2(N__13427),
            .in3(N__13242),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20627));
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_8_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0ES07_8_LC_8_1_2 .LUT_INIT=16'b0000001011111111;
    LogicCell40 \uu2.w_addr_displaying_RNI0ES07_8_LC_8_1_2  (
            .in0(N__13241),
            .in1(N__13413),
            .in2(N__12990),
            .in3(N__21785),
            .lcout(\uu2.w_addr_displaying_RNI0ES07Z0Z_8 ),
            .ltout(\uu2.w_addr_displaying_RNI0ES07Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_4_LC_8_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_4_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_4_LC_8_1_3 .LUT_INIT=16'b1010111101010000;
    LogicCell40 \uu2.w_addr_displaying_4_LC_8_1_3  (
            .in0(N__13417),
            .in1(_gnd_net_),
            .in2(N__12960),
            .in3(N__13372),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20627));
    defparam \uu2.w_addr_displaying_5_LC_8_1_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_8_1_4 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \uu2.w_addr_displaying_5_LC_8_1_4  (
            .in0(N__13373),
            .in1(N__15876),
            .in2(N__13305),
            .in3(N__13418),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_8C_net ),
            .ce(),
            .sr(N__20627));
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_8_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNO_0_6_LC_8_1_5 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNO_0_6_LC_8_1_5  (
            .in0(N__13295),
            .in1(_gnd_net_),
            .in2(N__13426),
            .in3(N__13371),
            .lcout(\uu2.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_8_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_8_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_8_1_6 .LUT_INIT=16'b0001010000011000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_0_6_LC_8_1_6  (
            .in0(N__13183),
            .in1(N__16603),
            .in2(N__13256),
            .in3(N__13293),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_8_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_8_1_7 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNIA3PF1_6_LC_8_1_7  (
            .in0(N__13294),
            .in1(N__13240),
            .in2(N__16617),
            .in3(N__13184),
            .lcout(\uu2.bitmap_pmux_sn_N_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_290_LC_8_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_8_2_0 .LUT_INIT=16'b0000011000011101;
    LogicCell40 \uu2.bitmap_290_LC_8_2_0  (
            .in0(N__14657),
            .in1(N__14482),
            .in2(N__13468),
            .in3(N__13559),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \uu2.bitmap_194_LC_8_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_8_2_1 .LUT_INIT=16'b0001000000010101;
    LogicCell40 \uu2.bitmap_194_LC_8_2_1  (
            .in0(N__13558),
            .in1(N__13455),
            .in2(N__14491),
            .in3(N__14656),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \uu2.bitmap_66_LC_8_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_8_2_2 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \uu2.bitmap_66_LC_8_2_2  (
            .in0(N__14659),
            .in1(N__14486),
            .in2(N__13469),
            .in3(N__13561),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \uu2.bitmap_RNIPDM31_66_LC_8_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIPDM31_66_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIPDM31_66_LC_8_2_3 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \uu2.bitmap_RNIPDM31_66_LC_8_2_3  (
            .in0(N__13149),
            .in1(N__16602),
            .in2(N__16541),
            .in3(N__13143),
            .lcout(\uu2.bitmap_pmux_20_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_8_2_4 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_8_2_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_162_LC_8_2_4  (
            .in0(N__14655),
            .in1(N__14478),
            .in2(N__13467),
            .in3(N__13557),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \uu2.bitmap_34_LC_8_2_5 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_8_2_5 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_34_LC_8_2_5  (
            .in0(N__13560),
            .in1(N__13459),
            .in2(N__14492),
            .in3(N__14658),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \uu2.bitmap_RNIP2JO1_34_LC_8_2_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIP2JO1_34_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIP2JO1_34_LC_8_2_6 .LUT_INIT=16'b0000110011111010;
    LogicCell40 \uu2.bitmap_RNIP2JO1_34_LC_8_2_6  (
            .in0(N__13803),
            .in1(N__13797),
            .in2(N__13791),
            .in3(N__13749),
            .lcout(\uu2.bitmap_RNIP2JO1Z0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_69_LC_8_2_7 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_8_2_7 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_69_LC_8_2_7  (
            .in0(N__13562),
            .in1(N__13463),
            .in2(N__14493),
            .in3(N__14660),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_290C_net ),
            .ce(),
            .sr(N__20625));
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_2_LC_8_3_0 .LUT_INIT=16'b0100010011000000;
    LogicCell40 \Lab_UT.dictrl.next_state_2_LC_8_3_0  (
            .in0(N__14787),
            .in1(N__18480),
            .in2(N__14760),
            .in3(N__18347),
            .lcout(\Lab_UT.dictrl.next_state_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22256),
            .ce(N__18771),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNI3JI86_3_LC_8_3_1  (
            .in0(N__17797),
            .in1(N__13728),
            .in2(_gnd_net_),
            .in3(N__13682),
            .lcout(\Lab_UT.sec2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNITCI86_0_LC_8_3_2  (
            .in0(N__13649),
            .in1(N__14360),
            .in2(_gnd_net_),
            .in3(N__17798),
            .lcout(\Lab_UT.sec2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI7FF76_3_LC_8_3_3  (
            .in0(N__17801),
            .in1(N__16697),
            .in2(_gnd_net_),
            .in3(N__13620),
            .lcout(\Lab_UT.min2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI3NT66_0_LC_8_3_4  (
            .in0(N__13590),
            .in1(N__17100),
            .in2(_gnd_net_),
            .in3(N__17800),
            .lcout(\Lab_UT.min1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI9TT66_3_LC_8_3_6  (
            .in0(N__13536),
            .in1(N__13509),
            .in2(_gnd_net_),
            .in3(N__17799),
            .lcout(\Lab_UT.min1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_215_LC_8_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_8_4_0 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_215_LC_8_4_0  (
            .in0(N__13827),
            .in1(N__14372),
            .in2(N__14115),
            .in3(N__14064),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIOPSS_212_LC_8_4_1 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \uu2.bitmap_RNIOPSS_212_LC_8_4_1  (
            .in0(N__14037),
            .in1(N__16405),
            .in2(N__14019),
            .in3(N__14031),
            .lcout(\uu2.bitmap_pmux_17_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_0_LC_8_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_8_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__15880),
            .in2(_gnd_net_),
            .in3(N__14017),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \uu2.bitmap_RNI65TM_72_LC_8_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI65TM_72_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI65TM_72_LC_8_4_3 .LUT_INIT=16'b0011000100111101;
    LogicCell40 \uu2.bitmap_RNI65TM_72_LC_8_4_3  (
            .in0(N__13983),
            .in1(N__16404),
            .in2(N__14018),
            .in3(N__13989),
            .lcout(\uu2.bitmap_pmux_16_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_7_LC_8_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_7_LC_8_4_4 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \uu2.w_addr_displaying_fast_7_LC_8_4_4  (
            .in0(N__16406),
            .in1(N__15881),
            .in2(_gnd_net_),
            .in3(N__15917),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \uu2.bitmap_72_LC_8_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_8_4_5 .LUT_INIT=16'b0001001100001101;
    LogicCell40 \uu2.bitmap_72_LC_8_4_5  (
            .in0(N__13964),
            .in1(N__13936),
            .in2(N__14150),
            .in3(N__13898),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \uu2.bitmap_200_LC_8_4_6 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_8_4_6 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_200_LC_8_4_6  (
            .in0(N__13896),
            .in1(N__14133),
            .in2(N__13945),
            .in3(N__13962),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \uu2.bitmap_296_LC_8_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_8_4_7 .LUT_INIT=16'b0001001000110101;
    LogicCell40 \uu2.bitmap_296_LC_8_4_7  (
            .in0(N__13963),
            .in1(N__13935),
            .in2(N__14149),
            .in3(N__13897),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_215C_net ),
            .ce(),
            .sr(N__20622));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI1T0O5_1_LC_8_5_0  (
            .in0(N__17796),
            .in1(N__13872),
            .in2(_gnd_net_),
            .in3(N__14591),
            .lcout(\Lab_UT.sec1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_8_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_8_5_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI5PT66_1_LC_8_5_1  (
            .in0(N__14520),
            .in1(N__17025),
            .in2(_gnd_net_),
            .in3(N__17795),
            .lcout(\Lab_UT.min1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_8_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_8_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_esr_RNI3V0O5_2_LC_8_5_2  (
            .in0(N__17794),
            .in1(N__14451),
            .in2(_gnd_net_),
            .in3(N__14421),
            .lcout(\Lab_UT.sec1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_8_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_8_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_2_LC_8_5_3  (
            .in0(_gnd_net_),
            .in1(N__14356),
            .in2(_gnd_net_),
            .in3(N__17892),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_5_4 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_5_4  (
            .in0(N__14301),
            .in1(N__20932),
            .in2(N__14262),
            .in3(N__16983),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_5_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_8_5_5  (
            .in0(N__16984),
            .in1(N__14242),
            .in2(N__14217),
            .in3(N__14214),
            .lcout(\Lab_UT.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22241),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_5_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_8_5_7  (
            .in0(N__16880),
            .in1(N__17300),
            .in2(N__16706),
            .in3(N__16748),
            .lcout(\Lab_UT.didp.countrce3.ce_12_0_a6_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_8_6_0 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_3_0_LC_8_6_0  (
            .in0(N__16878),
            .in1(N__14681),
            .in2(N__17611),
            .in3(N__14602),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxa_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_RNI3BF76_1_LC_8_6_1  (
            .in0(N__14603),
            .in1(N__17786),
            .in2(_gnd_net_),
            .in3(N__16879),
            .lcout(\Lab_UT.min2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_8_6_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI7RT66_2_LC_8_6_2  (
            .in0(N__17603),
            .in1(_gnd_net_),
            .in2(N__17802),
            .in3(N__14682),
            .lcout(\Lab_UT.min1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_esr_1_LC_8_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_esr_1_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21389),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22233),
            .ce(N__14628),
            .sr(N__20672));
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_1_LC_8_6_4 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_1_LC_8_6_4  (
            .in0(N__18206),
            .in1(N__18092),
            .in2(N__17998),
            .in3(N__14604),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_8_6_5 .LUT_INIT=16'b1111101111110000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_8_6_5  (
            .in0(N__14592),
            .in1(N__18093),
            .in2(N__14562),
            .in3(N__14533),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_8_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_8_6_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIH15E_0_2_LC_8_6_6  (
            .in0(N__17976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18202),
            .lcout(\Lab_UT.dispString.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNI5MKI1_LC_8_7_0  (
            .in0(N__19507),
            .in1(N__19883),
            .in2(N__18468),
            .in3(N__18330),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_ctle_LC_8_7_1  (
            .in0(N__14997),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20750),
            .lcout(\Lab_UT.bu_rx_data_rdy_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_8_7_2 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_8_7_2  (
            .in0(N__15074),
            .in1(N__15027),
            .in2(N__14826),
            .in3(N__14998),
            .lcout(\Lab_UT.dictrl.dicLdAMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22227),
            .ce(),
            .sr(N__20670));
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_LC_8_7_3 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_LC_8_7_3  (
            .in0(N__14999),
            .in1(N__15075),
            .in2(N__18363),
            .in3(N__18592),
            .lcout(\Lab_UT.dictrl.dicRun_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22227),
            .ce(),
            .sr(N__20670));
    defparam \Lab_UT.dictrl.state_ret_9_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_LC_8_7_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_9_LC_8_7_4 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_LC_8_7_4  (
            .in0(N__18591),
            .in1(N__15028),
            .in2(N__19133),
            .in3(N__15000),
            .lcout(\Lab_UT.dicLdSones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22227),
            .ce(),
            .sr(N__20670));
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_RNI9F571_LC_8_7_6  (
            .in0(N__18445),
            .in1(N__19882),
            .in2(_gnd_net_),
            .in3(N__14822),
            .lcout(\Lab_UT.LdAMones ),
            .ltout(\Lab_UT.LdAMones_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI14AG5_LC_8_7_7  (
            .in0(N__14843),
            .in1(N__18239),
            .in2(N__14799),
            .in3(N__14850),
            .lcout(\Lab_UT.loadalarm_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_8_8_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNI3FJ7D_LC_8_8_0  (
            .in0(N__14690),
            .in1(N__15308),
            .in2(_gnd_net_),
            .in3(N__14796),
            .lcout(\Lab_UT.next_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNI81O17_2_LC_8_8_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNI81O17_2_LC_8_8_1  (
            .in0(N__19282),
            .in1(N__15773),
            .in2(N__14720),
            .in3(N__18421),
            .lcout(\Lab_UT.dictrl.g0_1_mb_rn_0 ),
            .ltout(\Lab_UT.dictrl.g0_1_mb_rn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_2 .LUT_INIT=16'b0101000011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_2_LC_8_8_2  (
            .in0(N__14691),
            .in1(_gnd_net_),
            .in2(N__14790),
            .in3(N__15309),
            .lcout(\Lab_UT.state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22220),
            .ce(N__18507),
            .sr(N__20663));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_8_8_3 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNIFIQ9B_LC_8_8_3  (
            .in0(N__18299),
            .in1(N__14783),
            .in2(N__14753),
            .in3(N__18423),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_4 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__14716),
            .in2(N__14694),
            .in3(N__19286),
            .lcout(\Lab_UT.dictrl.state_i_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22220),
            .ce(N__18507),
            .sr(N__20663));
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_8_8_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_RNIR14R_LC_8_8_5  (
            .in0(N__18298),
            .in1(_gnd_net_),
            .in2(N__19293),
            .in3(N__18422),
            .lcout(\Lab_UT.dictrl.g0_1_mb_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_8_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_8_8_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_ess_RNINDRJ_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__18700),
            .in2(_gnd_net_),
            .in3(N__18297),
            .lcout(),
            .ltout(\Lab_UT.dictrl.un15_loadalarm_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_8_8_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_8_8_7 .LUT_INIT=16'b0011011111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI5S0R1_LC_8_8_7  (
            .in0(N__19103),
            .in1(N__18420),
            .in2(N__14853),
            .in3(N__19459),
            .lcout(\Lab_UT.dictrl.loadalarm_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUPT821_0_LC_8_9_0  (
            .in0(N__18930),
            .in1(N__17907),
            .in2(N__18824),
            .in3(N__15195),
            .lcout(\Lab_UT.next_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_0_LC_8_9_1  (
            .in0(N__15198),
            .in1(N__18823),
            .in2(N__18939),
            .in3(N__17910),
            .lcout(\Lab_UT.dictrl.state_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_LC_8_9_2  (
            .in0(N__18931),
            .in1(N__17908),
            .in2(N__18825),
            .in3(N__15196),
            .lcout(\Lab_UT.dictrl.state_0_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_0_LC_8_9_3  (
            .in0(N__15197),
            .in1(N__18822),
            .in2(N__18938),
            .in3(N__17909),
            .lcout(\Lab_UT.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNI78U61_LC_8_9_4  (
            .in0(N__18419),
            .in1(N__19458),
            .in2(N__15111),
            .in3(N__19831),
            .lcout(\Lab_UT.LdAStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_LC_8_9_5  (
            .in0(N__18671),
            .in1(_gnd_net_),
            .in2(N__18654),
            .in3(N__19254),
            .lcout(\Lab_UT.state_i_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6  (
            .in0(N__19253),
            .in1(N__18650),
            .in2(_gnd_net_),
            .in3(N__18670),
            .lcout(\Lab_UT.dictrl.stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_1_LC_8_9_7  (
            .in0(N__17164),
            .in1(N__17141),
            .in2(N__19628),
            .in3(N__19255),
            .lcout(Lab_UT_dictrl_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22214),
            .ce(N__18515),
            .sr(N__20671));
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNILQB86_1_LC_8_10_0  (
            .in0(N__19247),
            .in1(N__15152),
            .in2(N__15138),
            .in3(N__15112),
            .lcout(\Lab_UT.dictrl.next_state_RNILQB86Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_1_LC_8_10_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_LC_8_10_1  (
            .in0(N__15114),
            .in1(N__19595),
            .in2(N__17168),
            .in3(N__15153),
            .lcout(\Lab_UT.dictrl.next_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22206),
            .ce(N__18748),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_0_m2_0_LC_8_10_2  (
            .in0(N__14870),
            .in1(N__15164),
            .in2(N__15126),
            .in3(N__19471),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_20_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__g0_1_LC_8_10_3  (
            .in0(N__15113),
            .in1(N__19593),
            .in2(N__15090),
            .in3(N__15087),
            .lcout(),
            .ltout(\Lab_UT.next_state_1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_LC_8_10_4 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \Lab_UT.didp.g0_0_LC_8_10_4  (
            .in0(N__15063),
            .in1(N__14877),
            .in2(N__15036),
            .in3(N__15033),
            .lcout(\Lab_UT.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.g0_0_2_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.g0_0_2_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.g0_0_2_LC_8_10_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \Lab_UT.didp.g0_0_2_LC_8_10_5  (
            .in0(N__14980),
            .in1(N__14925),
            .in2(N__14915),
            .in3(N__19248),
            .lcout(\Lab_UT.didp.g0_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_LC_8_10_6  (
            .in0(N__14871),
            .in1(N__15165),
            .in2(N__19508),
            .in3(N__18684),
            .lcout(\Lab_UT.dictrl.N_20 ),
            .ltout(\Lab_UT.dictrl.N_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNITNH9H_3_LC_8_10_7  (
            .in0(N__19252),
            .in1(N__19594),
            .in2(N__14856),
            .in3(N__17140),
            .lcout(\Lab_UT.next_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_8_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m34_0_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__18455),
            .in2(_gnd_net_),
            .in3(N__19888),
            .lcout(\Lab_UT.dictrl.m34_0 ),
            .ltout(\Lab_UT.dictrl.m34_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m35_LC_8_11_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m35_LC_8_11_2  (
            .in0(N__15281),
            .in1(N__15490),
            .in2(N__15231),
            .in3(N__18336),
            .lcout(\Lab_UT.dictrl.next_state_1_3 ),
            .ltout(\Lab_UT.dictrl.next_state_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_8_11_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNINVFJ7_3_LC_8_11_3  (
            .in0(N__18629),
            .in1(_gnd_net_),
            .in2(N__15228),
            .in3(N__19231),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_8_11_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKOLT_0_2_LC_8_11_4  (
            .in0(N__19229),
            .in1(N__19601),
            .in2(_gnd_net_),
            .in3(N__18334),
            .lcout(\Lab_UT.dictrl.N_33_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_8_11_5 .LUT_INIT=16'b0000001000000010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIKOLT_2_LC_8_11_5  (
            .in0(N__18335),
            .in1(N__19230),
            .in2(N__19622),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_14_0_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_8_11_6 .LUT_INIT=16'b0010000001110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIN2PIH_1_LC_8_11_6  (
            .in0(N__19887),
            .in1(N__15171),
            .in2(N__15201),
            .in3(N__15288),
            .lcout(\Lab_UT.dictrl.N_26_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_3_LC_8_11_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Lab_UT.dictrl.next_state_3_LC_8_11_7  (
            .in0(N__18337),
            .in1(N__15180),
            .in2(N__15495),
            .in3(N__15282),
            .lcout(\Lab_UT.dictrl.next_state_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22200),
            .ce(N__18764),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_12_0 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_0_LC_8_12_0  (
            .in0(N__21466),
            .in1(N__15456),
            .in2(N__20140),
            .in3(N__18901),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIO0F67_LC_8_12_1  (
            .in0(N__19027),
            .in1(N__15273),
            .in2(N__15174),
            .in3(N__18902),
            .lcout(\Lab_UT.dictrl.N_60_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_8_12_2 .LUT_INIT=16'b0000101001100110;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_1_LC_8_12_2  (
            .in0(N__19920),
            .in1(N__20058),
            .in2(N__15486),
            .in3(N__18345),
            .lcout(\Lab_UT.dictrl.m19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \buart.Z_rx.shifter_RNIR1VT2_3_LC_8_12_3  (
            .in0(N__15457),
            .in1(N__21095),
            .in2(_gnd_net_),
            .in3(N__21467),
            .lcout(),
            .ltout(N_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4 .LUT_INIT=16'b0101000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNI27M74_LC_8_12_4  (
            .in0(N__19605),
            .in1(N__19134),
            .in2(N__15294),
            .in3(N__19496),
            .lcout(\Lab_UT.dictrl.G_6_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_8_12_5 .LUT_INIT=16'b1111101101010001;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNICD344_LC_8_12_5  (
            .in0(N__20128),
            .in1(N__21465),
            .in2(N__18913),
            .in3(N__18981),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNICDZ0Z344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_8_12_6 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIKMA19_LC_8_12_6  (
            .in0(N__15237),
            .in1(N__19028),
            .in2(N__15291),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_59_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_7 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m32_LC_8_12_7  (
            .in0(N__18557),
            .in1(N__19606),
            .in2(N__17253),
            .in3(N__18982),
            .lcout(\Lab_UT.dictrl.i8_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_13_0 .LUT_INIT=16'b1010101011111101;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_LC_8_13_0  (
            .in0(N__21437),
            .in1(N__15458),
            .in2(N__18905),
            .in3(N__20127),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNID8OZ0Z13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_x1_LC_8_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m22_x1_LC_8_13_1  (
            .in0(N__19338),
            .in1(N__21214),
            .in2(N__19775),
            .in3(N__19687),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m22_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m22_ns_LC_8_13_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.m22_ns_LC_8_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15267),
            .in3(N__15258),
            .lcout(\Lab_UT.dictrl.N_72_mux ),
            .ltout(\Lab_UT.dictrl.N_72_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_3 .LUT_INIT=16'b1100000011110011;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36V3_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__20125),
            .in2(N__15240),
            .in3(N__21436),
            .lcout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIB36VZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m7_a0_LC_8_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m7_a0_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m7_a0_LC_8_13_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.m7_a0_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(N__20196),
            .in2(_gnd_net_),
            .in3(N__19391),
            .lcout(m7_a0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_8_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_8_13_5 .LUT_INIT=16'b0011011100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4B1_LC_8_13_5  (
            .in0(N__19392),
            .in1(N__18887),
            .in2(N__20204),
            .in3(N__20126),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIIE4BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_8_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_8_13_6 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNID8O13_1_LC_8_13_6  (
            .in0(N__21435),
            .in1(_gnd_net_),
            .in2(N__15498),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m7_0_LC_8_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m7_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m7_0_LC_8_13_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dictrl.m7_0_LC_8_13_7  (
            .in0(N__15459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21438),
            .lcout(\Lab_UT.dictrl.N_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_5_4_LC_8_14_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.g0_5_4_LC_8_14_0  (
            .in0(N__15643),
            .in1(N__15668),
            .in2(N__18904),
            .in3(N__15377),
            .lcout(\Lab_UT.dictrl.g0_5Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_LC_8_14_1 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \Lab_UT.dictrl.g2_LC_8_14_1  (
            .in0(N__18886),
            .in1(N__19756),
            .in2(_gnd_net_),
            .in3(N__19345),
            .lcout(\Lab_UT.dictrl.gZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIT5E31_0_LC_8_14_2  (
            .in0(N__15642),
            .in1(N__15667),
            .in2(N__15441),
            .in3(N__15408),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_fast_esr_RNIT5E31Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_8_14_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_8_14_3 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNI0QVC1_0_LC_8_14_3  (
            .in0(N__15378),
            .in1(_gnd_net_),
            .in2(N__15354),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.g0_6_3 ),
            .ltout(\Lab_UT.dictrl.g0_6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_8_14_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_8_14_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI0CNA5_1_LC_8_14_4  (
            .in0(N__19885),
            .in1(N__15341),
            .in2(N__15327),
            .in3(N__15324),
            .lcout(\Lab_UT.dictrl.N_57_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_8_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_RNIS7QM1_LC_8_14_5  (
            .in0(N__17184),
            .in1(N__15831),
            .in2(N__15816),
            .in3(N__20205),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_RNITJ214_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15798),
            .in3(N__15795),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI7TE56_1_LC_8_14_7  (
            .in0(N__15789),
            .in1(N__15783),
            .in2(N__15777),
            .in3(N__19884),
            .lcout(\Lab_UT.dictrl.N_55_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_15_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_15_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_12_LC_8_15_3  (
            .in0(N__19773),
            .in1(N__19698),
            .in2(N__18903),
            .in3(N__15611),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_8_15_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_10_LC_8_15_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_10_LC_8_15_4  (
            .in0(N__15618),
            .in1(N__19346),
            .in2(N__15750),
            .in3(N__15740),
            .lcout(\Lab_UT.dictrl.N_72_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_8_15_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNO_11_LC_8_15_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNO_11_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__15669),
            .in2(_gnd_net_),
            .in3(N__15644),
            .lcout(\Lab_UT.dictrl.g0_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_rep1_LC_8_15_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_8_15_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_8_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15612),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22194),
            .ce(N__20791),
            .sr(N__20697));
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI43G8_3_LC_9_1_0  (
            .in0(N__16134),
            .in1(N__20333),
            .in2(N__15528),
            .in3(N__16232),
            .lcout(\uu2.un3_w_addr_user_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_9_1_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_9_1_1  (
            .in0(N__16234),
            .in1(N__16139),
            .in2(N__20342),
            .in3(N__21839),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15960),
            .sr(N__15948));
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI2OE4_8_LC_9_1_2  (
            .in0(N__15973),
            .in1(N__16153),
            .in2(_gnd_net_),
            .in3(N__21837),
            .lcout(),
            .ltout(\uu2.un3_w_addr_user_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_RNIINVH_4_LC_9_1_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uu2.w_addr_user_RNIINVH_4_LC_9_1_3  (
            .in0(N__16192),
            .in1(N__16299),
            .in2(N__16269),
            .in3(N__16266),
            .lcout(\uu2.un3_w_addr_user ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_4 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_w_addr_user.counter_gen_label_4__un404_ci_LC_9_1_4  (
            .in0(N__20340),
            .in1(N__21838),
            .in2(N__16140),
            .in3(N__16233),
            .lcout(\uu2.un404_ci ),
            .ltout(\uu2.un404_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_7_LC_9_1_5 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu2.w_addr_user_nesr_7_LC_9_1_5  (
            .in0(N__16154),
            .in1(N__16040),
            .in2(N__16197),
            .in3(N__16194),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15960),
            .sr(N__15948));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_9_1_6  (
            .in0(N__16135),
            .in1(N__21786),
            .in2(_gnd_net_),
            .in3(N__16122),
            .lcout(\uu2.mem0.w_addr_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_9_1_7 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_9_1_7  (
            .in0(N__16041),
            .in1(N__16001),
            .in2(N__15990),
            .in3(N__15974),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_3C_net ),
            .ce(N__15960),
            .sr(N__15948));
    defparam \uu2.w_addr_displaying_7_LC_9_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_7_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_7_LC_9_2_0 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uu2.w_addr_displaying_7_LC_9_2_0  (
            .in0(N__15867),
            .in1(N__15918),
            .in2(_gnd_net_),
            .in3(N__16616),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20628));
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_rep1_LC_9_2_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_rep1_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(N__15866),
            .in2(_gnd_net_),
            .in3(N__16529),
            .lcout(\uu2.w_addr_displaying_0_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20628));
    defparam \uu2.bitmap_111_LC_9_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_9_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_9_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_9_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17547),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_7C_net ),
            .ce(),
            .sr(N__20628));
    defparam \uu2.bitmap_314_LC_9_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_9_3_0 .LUT_INIT=16'b0000011000011101;
    LogicCell40 \uu2.bitmap_314_LC_9_3_0  (
            .in0(N__16911),
            .in1(N__17708),
            .in2(N__16446),
            .in3(N__16473),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20626));
    defparam \uu2.bitmap_218_LC_9_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_9_3_1 .LUT_INIT=16'b0001000000010101;
    LogicCell40 \uu2.bitmap_218_LC_9_3_1  (
            .in0(N__16472),
            .in1(N__16432),
            .in2(N__17718),
            .in3(N__16910),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20626));
    defparam \uu2.bitmap_90_LC_9_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_9_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_9_3_2 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \uu2.bitmap_90_LC_9_3_2  (
            .in0(N__16913),
            .in1(N__17712),
            .in2(N__16447),
            .in3(N__16475),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20626));
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIJ4K41_90_LC_9_3_3 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \uu2.bitmap_RNIJ4K41_90_LC_9_3_3  (
            .in0(N__16601),
            .in1(N__16563),
            .in2(N__16540),
            .in3(N__16497),
            .lcout(\uu2.bitmap_pmux_19_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_9_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_9_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_9_3_4 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_186_LC_9_3_4  (
            .in0(N__16909),
            .in1(N__17704),
            .in2(N__16445),
            .in3(N__16471),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20626));
    defparam \uu2.bitmap_58_LC_9_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_9_3_5 .LUT_INIT=16'b1111011001111101;
    LogicCell40 \uu2.bitmap_58_LC_9_3_5  (
            .in0(N__16474),
            .in1(N__16436),
            .in2(N__17719),
            .in3(N__16912),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__20626));
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIKGSI_58_LC_9_3_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIKGSI_58_LC_9_3_6  (
            .in0(N__16403),
            .in1(N__16383),
            .in2(_gnd_net_),
            .in3(N__16377),
            .lcout(),
            .ltout(\uu2.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIM5E21_314_LC_9_3_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uu2.bitmap_RNIM5E21_314_LC_9_3_7  (
            .in0(_gnd_net_),
            .in1(N__16370),
            .in2(N__16356),
            .in3(N__16347),
            .lcout(\uu2.bitmap_RNIM5E21Z0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_9_4_7  (
            .in0(N__16662),
            .in1(N__16668),
            .in2(N__17370),
            .in3(N__16702),
            .lcout(\Lab_UT.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22257),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_5_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__16882),
            .in2(_gnd_net_),
            .in3(N__17299),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_5_1 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_5_1  (
            .in0(N__17329),
            .in1(N__20933),
            .in2(N__16764),
            .in3(N__16742),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_5_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_9_5_2  (
            .in0(N__16743),
            .in1(N__17359),
            .in2(N__16761),
            .in3(N__16661),
            .lcout(\Lab_UT.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22249),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_9_5_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__17028),
            .in2(_gnd_net_),
            .in3(N__17102),
            .lcout(\Lab_UT.didp.reset_12_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_3_LC_9_5_4  (
            .in0(N__16741),
            .in1(N__16881),
            .in2(_gnd_net_),
            .in3(N__17298),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_9_5_5  (
            .in0(N__17328),
            .in1(N__21134),
            .in2(N__16710),
            .in3(N__16701),
            .lcout(\Lab_UT.didp.countrce3.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIBN0Q1_2_LC_9_5_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNIBN0Q1_2_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__17399),
            .in2(_gnd_net_),
            .in3(N__17330),
            .lcout(\Lab_UT.didp.un1_dicLdMones_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_5_7 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_9_5_7  (
            .in0(N__16883),
            .in1(N__16851),
            .in2(N__16650),
            .in3(N__17358),
            .lcout(\Lab_UT.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22249),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_9_6_0 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_9_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.sec_clkD_LC_9_6_0  (
            .in0(N__17546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uu0_sec_clkD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_9_6_2 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_9_6_2  (
            .in0(N__17316),
            .in1(N__20051),
            .in2(_gnd_net_),
            .in3(N__17292),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_9_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_9_6_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dispString.cnt_RNIFV4E_1_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__18112),
            .in2(_gnd_net_),
            .in3(N__18207),
            .lcout(\Lab_UT.dispString.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_6_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_6_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_9_6_4  (
            .in0(N__21395),
            .in1(N__17026),
            .in2(N__17676),
            .in3(N__17103),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_9_6_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_9_6_5  (
            .in0(N__17027),
            .in1(N__16838),
            .in2(N__17040),
            .in3(N__16781),
            .lcout(\Lab_UT.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22242),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_9_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_9_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNI1HI86_2_LC_9_6_6  (
            .in0(N__16978),
            .in1(N__17773),
            .in2(_gnd_net_),
            .in3(N__16947),
            .lcout(\Lab_UT.sec2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_7 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_1_LC_9_6_7  (
            .in0(N__17293),
            .in1(N__16884),
            .in2(N__21396),
            .in3(N__17317),
            .lcout(\Lab_UT.didp.countrce3.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_9_7_0 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_9_7_0  (
            .in0(N__16780),
            .in1(N__17610),
            .in2(N__17580),
            .in3(N__16842),
            .lcout(\Lab_UT.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22234),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIHGGI1_3_LC_9_7_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNIHGGI1_3_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__16809),
            .in2(_gnd_net_),
            .in3(N__17675),
            .lcout(\Lab_UT.didp.un1_dicLdMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_9_7_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIVEI86_1_LC_9_7_3  (
            .in0(N__17882),
            .in1(N__17832),
            .in2(_gnd_net_),
            .in3(N__17774),
            .lcout(\Lab_UT.sec2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_7_4 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_9_7_4  (
            .in0(N__17674),
            .in1(N__20926),
            .in2(N__17631),
            .in3(N__17609),
            .lcout(\Lab_UT.didp.countrce4.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_9_7_5 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_9_7_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__17558),
            .in2(_gnd_net_),
            .in3(N__17535),
            .lcout(oneSecStrb),
            .ltout(oneSecStrb_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIKUO21_2_LC_9_7_6 .LUT_INIT=16'b0001000110001001;
    LogicCell40 \Lab_UT.dispString.cnt_RNIKUO21_2_LC_9_7_6  (
            .in0(N__18117),
            .in1(N__17980),
            .in2(N__17433),
            .in3(N__18222),
            .lcout(\Lab_UT.dispString.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_7_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_7_7 .LUT_INIT=16'b0000110000001001;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_9_7_7  (
            .in0(N__17403),
            .in1(N__17376),
            .in2(N__17369),
            .in3(N__17331),
            .lcout(\Lab_UT.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22234),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_8_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_9_8_0 .LUT_INIT=16'b0011001000110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_LC_9_8_0  (
            .in0(N__19287),
            .in1(N__19148),
            .in2(N__18804),
            .in3(N__19055),
            .lcout(\Lab_UT.dictrl.state_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22228),
            .ce(N__18519),
            .sr(N__20667));
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_9_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_9_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_fast_ess_LC_9_8_1 .LUT_INIT=16'b0000111100011101;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_fast_ess_LC_9_8_1  (
            .in0(N__19056),
            .in1(N__18803),
            .in2(N__19152),
            .in3(N__19288),
            .lcout(\Lab_UT.dictrl.state_ret_2_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22228),
            .ce(N__18519),
            .sr(N__20667));
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_9_8_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_6_ess_LC_9_8_3 .LUT_INIT=16'b0000000111111101;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_ess_LC_9_8_3  (
            .in0(N__17172),
            .in1(N__19289),
            .in2(N__19629),
            .in3(N__17145),
            .lcout(\Lab_UT.dictrl.state_i_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22228),
            .ce(N__18519),
            .sr(N__20667));
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_9_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_9_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.next_state_1_3_0__m19_1_0_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__18704),
            .in2(_gnd_net_),
            .in3(N__18301),
            .lcout(\Lab_UT.dictrl.m19_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_esr_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_esr_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_esr_LC_9_8_5 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_esr_LC_9_8_5  (
            .in0(N__19290),
            .in1(N__18672),
            .in2(N__18649),
            .in3(N__18602),
            .lcout(\Lab_UT.dictrl.next_state66_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22228),
            .ce(N__18519),
            .sr(N__20667));
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_RNICG571_LC_9_8_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_RNICG571_LC_9_8_6  (
            .in0(N__18418),
            .in1(N__18359),
            .in2(_gnd_net_),
            .in3(N__18300),
            .lcout(\Lab_UT.LdASones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_9_9_2 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_9_9_2  (
            .in0(N__17975),
            .in1(N__18221),
            .in2(_gnd_net_),
            .in3(N__18118),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22221),
            .ce(),
            .sr(N__20673));
    defparam \Lab_UT.dictrl.g1_8_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_8_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_8_LC_9_10_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.g1_8_LC_9_10_0  (
            .in0(N__19776),
            .in1(N__19361),
            .in2(N__18914),
            .in3(N__19697),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_9_10_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIVDGG2_LC_9_10_1  (
            .in0(N__20095),
            .in1(N__17928),
            .in2(N__17916),
            .in3(N__19864),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_14_0_a2_4_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_9_10_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIIANV3_0_LC_9_10_2  (
            .in0(N__19304),
            .in1(N__19257),
            .in2(N__17913),
            .in3(N__18950),
            .lcout(\Lab_UT.dictrl.G_14_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_9_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_9_10_3 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_RNI0FPF_LC_9_10_3  (
            .in0(N__19360),
            .in1(N__18906),
            .in2(_gnd_net_),
            .in3(N__19777),
            .lcout(),
            .ltout(shifter_1_rep1_RNI0FPF_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_9_10_4 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSR2_LC_9_10_4  (
            .in0(N__19863),
            .in1(N__20094),
            .in2(N__18954),
            .in3(N__21494),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNI6QSRZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_9_10_5 .LUT_INIT=16'b1000101000001010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIG91L6_0_LC_9_10_5  (
            .in0(N__18951),
            .in1(N__21152),
            .in2(N__18942),
            .in3(N__19460),
            .lcout(\Lab_UT.dictrl.G_14_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_9_10_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_9_10_6 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_RNIR8D62_LC_9_10_6  (
            .in0(N__19778),
            .in1(N__21495),
            .in2(N__18915),
            .in3(N__19362),
            .lcout(),
            .ltout(N_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_9_10_7 .LUT_INIT=16'b1010000000100010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI53C16_0_LC_9_10_7  (
            .in0(N__18837),
            .in1(N__21153),
            .in2(N__18828),
            .in3(N__19461),
            .lcout(\Lab_UT.dictrl.N_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_11_0 .LUT_INIT=16'b0001101100010001;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_0_0_LC_9_11_0  (
            .in0(N__19618),
            .in1(N__20214),
            .in2(N__19164),
            .in3(N__19136),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_0Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.next_state_0_LC_9_11_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.dictrl.next_state_0_LC_9_11_1  (
            .in0(N__18799),
            .in1(_gnd_net_),
            .in2(N__18774),
            .in3(N__18714),
            .lcout(\Lab_UT.dictrl.next_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22207),
            .ce(N__18763),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m14_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m14_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m14_LC_9_11_2 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \Lab_UT.dictrl.m14_LC_9_11_2  (
            .in0(N__21091),
            .in1(N__21492),
            .in2(_gnd_net_),
            .in3(N__19041),
            .lcout(\Lab_UT.dictrl.N_15_0 ),
            .ltout(\Lab_UT.dictrl.N_15_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_11_3 .LUT_INIT=16'b1111000010111011;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNICL796_0_LC_9_11_3  (
            .in0(N__21093),
            .in1(N__20229),
            .in2(N__18720),
            .in3(N__19506),
            .lcout(\Lab_UT.dictrl.N_60 ),
            .ltout(\Lab_UT.dictrl.N_60_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_4 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_1_0_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(N__18962),
            .in2(N__18717),
            .in3(N__19917),
            .lcout(\Lab_UT.dictrl.next_state_RNO_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \Lab_UT.dictrl.next_state_RNIMMQU_0_LC_9_11_6  (
            .in0(N__19305),
            .in1(N__19291),
            .in2(_gnd_net_),
            .in3(N__19916),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_latmux_d_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_13_RNIIQPMC_LC_9_11_7  (
            .in0(N__18963),
            .in1(N__19292),
            .in2(N__19167),
            .in3(N__19163),
            .lcout(\Lab_UT.dictrl.state_ret_13_RNIIQPMCZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_0 .LUT_INIT=16'b0111010101110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_9_RNIUN0N1_LC_9_12_0  (
            .in0(N__19500),
            .in1(N__19135),
            .in2(N__19627),
            .in3(N__19910),
            .lcout(\Lab_UT.dictrl.G_6_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_12_2 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_RNI055E2_0_LC_9_12_2  (
            .in0(N__21237),
            .in1(N__20874),
            .in2(N__21379),
            .in3(N__21486),
            .lcout(),
            .ltout(G_6_0_a6_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3 .LUT_INIT=16'b0011000001000100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIIJEG7_3_LC_9_12_3  (
            .in0(N__18999),
            .in1(N__19617),
            .in2(N__19077),
            .in3(N__19074),
            .lcout(),
            .ltout(\Lab_UT.dictrl.G_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_9_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_9_12_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIBLGFF_0_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__19407),
            .in2(N__19068),
            .in3(N__19065),
            .lcout(\Lab_UT.dictrl.state_0_esr_RNIBLGFFZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_9_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_5_0_LC_9_12_5 .LUT_INIT=16'b0001101110011011;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_5_0_LC_9_12_5  (
            .in0(N__19909),
            .in1(N__21236),
            .in2(N__21493),
            .in3(N__19040),
            .lcout(\Lab_UT.dictrl.next_state_RNO_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIDUKB5_0_LC_9_12_6  (
            .in0(N__19501),
            .in1(N__18998),
            .in2(_gnd_net_),
            .in3(N__18986),
            .lcout(\Lab_UT.dictrl.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_7 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_2_0_LC_9_12_7  (
            .in0(N__19935),
            .in1(N__20228),
            .in2(N__21135),
            .in3(N__19502),
            .lcout(\Lab_UT.dictrl.i8_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_9_13_1 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4B1_LC_9_13_1  (
            .in0(N__21234),
            .in1(N__20203),
            .in2(N__20156),
            .in3(N__19393),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_0_rep1_esr_RNIJE4BZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_9_13_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \Lab_UT.dictrl.state_0_0_rep1_esr_RNIE8O13_0_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20061),
            .in3(N__21482),
            .lcout(\Lab_UT.dictrl.N_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_9_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_4_0_LC_9_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_4_0_LC_9_13_3  (
            .in0(N__20861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20007),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_state_RNO_4Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_9_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.next_state_RNO_3_0_LC_9_13_4 .LUT_INIT=16'b1011111101010101;
    LogicCell40 \Lab_UT.dictrl.next_state_RNO_3_0_LC_9_13_4  (
            .in0(N__19928),
            .in1(N__19640),
            .in2(N__19944),
            .in3(N__19941),
            .lcout(\Lab_UT.dictrl.i9_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_9_13_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_9_13_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \buart.Z_rx.shifter_0_rep1_RNINSO21_LC_9_13_6  (
            .in0(N__19927),
            .in1(N__21235),
            .in2(N__19779),
            .in3(N__19691),
            .lcout(),
            .ltout(G_6_0_a6_3_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_9_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_9_13_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNINQBN3_0_LC_9_13_7  (
            .in0(N__19641),
            .in1(N__19626),
            .in2(N__19515),
            .in3(N__19512),
            .lcout(\Lab_UT.dictrl.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20848),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__20796),
            .sr(N__20698));
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_14_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_14_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_9_14_2  (
            .in0(N__20847),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__20796),
            .sr(N__20698));
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_9_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_9_14_4 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_RNI055E2_LC_9_14_4  (
            .in0(N__20846),
            .in1(N__21480),
            .in2(N__21335),
            .in3(N__21233),
            .lcout(N_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_9_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21115),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22195),
            .ce(N__20796),
            .sr(N__20698));
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_11_1_0 .LUT_INIT=16'b1111100111111100;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_11_1_0  (
            .in0(N__21522),
            .in1(N__21558),
            .in2(N__20463),
            .in3(N__21583),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(),
            .sr(N__20699));
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_11_1_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_11_1_1  (
            .in0(N__21581),
            .in1(N__20461),
            .in2(_gnd_net_),
            .in3(N__21521),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(),
            .sr(N__20699));
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_11_1_2 .LUT_INIT=16'b1111111110010110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_11_1_2  (
            .in0(N__21603),
            .in1(N__21501),
            .in2(N__21588),
            .in3(N__20457),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(),
            .sr(N__20699));
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_11_1_3 .LUT_INIT=16'b0000100100000110;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_11_1_3  (
            .in0(N__21582),
            .in1(N__21609),
            .in2(N__20462),
            .in3(N__21540),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22273),
            .ce(),
            .sr(N__20699));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_1_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_11_1_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_11_1_4  (
            .in0(_gnd_net_),
            .in1(N__20453),
            .in2(_gnd_net_),
            .in3(N__21580),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_11_1_5  (
            .in0(N__20343),
            .in1(N__21805),
            .in2(_gnd_net_),
            .in3(N__20301),
            .lcout(\uu2.mem0.w_addr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_11_1_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_11_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_11_1_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_11_1_6  (
            .in0(N__21807),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21879),
            .lcout(\uu2.mem0.w_data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_11_1_7  (
            .in0(N__21840),
            .in1(N__21806),
            .in2(_gnd_net_),
            .in3(N__21693),
            .lcout(\uu2.mem0.w_addr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_11_2_0  (
            .in0(N__21519),
            .in1(N__21556),
            .in2(_gnd_net_),
            .in3(N__21584),
            .lcout(\buart.Z_tx.un1_bitcount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(N__21954),
            .in2(_gnd_net_),
            .in3(N__21938),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22271),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21937),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22271),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__21602),
            .in2(_gnd_net_),
            .in3(N__21518),
            .lcout(),
            .ltout(\buart.Z_tx.uart_busy_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6 .LUT_INIT=16'b1110111100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_11_2_6  (
            .in0(N__21538),
            .in1(N__21555),
            .in2(N__21591),
            .in3(N__21894),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_11_2_7  (
            .in0(N__21557),
            .in1(N__21539),
            .in2(N__21525),
            .in3(N__21520),
            .lcout(\buart.Z_tx.un1_bitcount_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_12_2_0  (
            .in0(_gnd_net_),
            .in1(N__21953),
            .in2(N__21939),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_2_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_12_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21918),
            .in3(N__22296),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__22274),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_12_2_2  (
            .in0(N__21896),
            .in1(N__21963),
            .in2(_gnd_net_),
            .in3(N__22293),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__22274),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_12_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21990),
            .in3(N__22290),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__22274),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_12_2_4  (
            .in0(N__21897),
            .in1(_gnd_net_),
            .in2(N__22002),
            .in3(N__22287),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__22274),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_12_2_5  (
            .in0(N__21977),
            .in1(N__21895),
            .in2(_gnd_net_),
            .in3(N__22284),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22274),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_12_2_6  (
            .in0(N__21998),
            .in1(N__21986),
            .in2(N__21978),
            .in3(N__21962),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_12_2_7  (
            .in0(N__21952),
            .in1(N__21933),
            .in2(N__21917),
            .in3(N__21903),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
