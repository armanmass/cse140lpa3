// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     May 20 2019 23:49:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "latticehx1k" view "INTERFACE"

module latticehx1k (
    led,
    o_serial_data,
    to_ir,
    sd,
    from_pc,
    clk_in);

    output [4:0] led;
    output o_serial_data;
    output to_ir;
    output sd;
    input from_pc;
    input clk_in;

    wire N__21862;
    wire N__21861;
    wire N__21860;
    wire N__21853;
    wire N__21852;
    wire N__21851;
    wire N__21844;
    wire N__21843;
    wire N__21842;
    wire N__21835;
    wire N__21834;
    wire N__21833;
    wire N__21826;
    wire N__21825;
    wire N__21824;
    wire N__21817;
    wire N__21816;
    wire N__21815;
    wire N__21808;
    wire N__21807;
    wire N__21806;
    wire N__21799;
    wire N__21798;
    wire N__21797;
    wire N__21790;
    wire N__21789;
    wire N__21788;
    wire N__21781;
    wire N__21780;
    wire N__21779;
    wire N__21762;
    wire N__21759;
    wire N__21758;
    wire N__21757;
    wire N__21756;
    wire N__21755;
    wire N__21752;
    wire N__21743;
    wire N__21738;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21730;
    wire N__21729;
    wire N__21720;
    wire N__21717;
    wire N__21714;
    wire N__21713;
    wire N__21712;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21689;
    wire N__21684;
    wire N__21681;
    wire N__21680;
    wire N__21675;
    wire N__21672;
    wire N__21671;
    wire N__21670;
    wire N__21669;
    wire N__21668;
    wire N__21667;
    wire N__21666;
    wire N__21665;
    wire N__21664;
    wire N__21663;
    wire N__21662;
    wire N__21661;
    wire N__21660;
    wire N__21659;
    wire N__21658;
    wire N__21657;
    wire N__21656;
    wire N__21655;
    wire N__21654;
    wire N__21653;
    wire N__21652;
    wire N__21651;
    wire N__21650;
    wire N__21649;
    wire N__21648;
    wire N__21647;
    wire N__21646;
    wire N__21645;
    wire N__21644;
    wire N__21643;
    wire N__21642;
    wire N__21641;
    wire N__21640;
    wire N__21639;
    wire N__21638;
    wire N__21637;
    wire N__21636;
    wire N__21635;
    wire N__21634;
    wire N__21633;
    wire N__21632;
    wire N__21631;
    wire N__21630;
    wire N__21629;
    wire N__21628;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21624;
    wire N__21623;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21615;
    wire N__21614;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21610;
    wire N__21609;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21601;
    wire N__21600;
    wire N__21599;
    wire N__21598;
    wire N__21597;
    wire N__21596;
    wire N__21595;
    wire N__21594;
    wire N__21593;
    wire N__21592;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21420;
    wire N__21419;
    wire N__21418;
    wire N__21417;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21397;
    wire N__21396;
    wire N__21393;
    wire N__21392;
    wire N__21391;
    wire N__21388;
    wire N__21383;
    wire N__21380;
    wire N__21375;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21334;
    wire N__21333;
    wire N__21332;
    wire N__21329;
    wire N__21328;
    wire N__21327;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21313;
    wire N__21310;
    wire N__21305;
    wire N__21302;
    wire N__21297;
    wire N__21292;
    wire N__21289;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21260;
    wire N__21259;
    wire N__21256;
    wire N__21255;
    wire N__21252;
    wire N__21251;
    wire N__21250;
    wire N__21247;
    wire N__21244;
    wire N__21243;
    wire N__21240;
    wire N__21239;
    wire N__21238;
    wire N__21237;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21217;
    wire N__21216;
    wire N__21213;
    wire N__21212;
    wire N__21211;
    wire N__21208;
    wire N__21205;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21180;
    wire N__21177;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21165;
    wire N__21160;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21141;
    wire N__21134;
    wire N__21129;
    wire N__21122;
    wire N__21105;
    wire N__21104;
    wire N__21103;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21099;
    wire N__21098;
    wire N__21097;
    wire N__21096;
    wire N__21093;
    wire N__21092;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21084;
    wire N__21083;
    wire N__21080;
    wire N__21079;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21053;
    wire N__21050;
    wire N__21049;
    wire N__21048;
    wire N__21045;
    wire N__21044;
    wire N__21041;
    wire N__21032;
    wire N__21029;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21021;
    wire N__21020;
    wire N__21013;
    wire N__21002;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20981;
    wire N__20978;
    wire N__20975;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20959;
    wire N__20956;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20931;
    wire N__20930;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20914;
    wire N__20911;
    wire N__20908;
    wire N__20907;
    wire N__20906;
    wire N__20903;
    wire N__20894;
    wire N__20893;
    wire N__20888;
    wire N__20887;
    wire N__20886;
    wire N__20885;
    wire N__20884;
    wire N__20883;
    wire N__20882;
    wire N__20881;
    wire N__20880;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20866;
    wire N__20863;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20831;
    wire N__20828;
    wire N__20823;
    wire N__20818;
    wire N__20815;
    wire N__20810;
    wire N__20803;
    wire N__20796;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20765;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20757;
    wire N__20756;
    wire N__20755;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20744;
    wire N__20743;
    wire N__20742;
    wire N__20741;
    wire N__20740;
    wire N__20739;
    wire N__20734;
    wire N__20733;
    wire N__20732;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20708;
    wire N__20705;
    wire N__20702;
    wire N__20699;
    wire N__20698;
    wire N__20697;
    wire N__20694;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20667;
    wire N__20662;
    wire N__20657;
    wire N__20654;
    wire N__20651;
    wire N__20648;
    wire N__20641;
    wire N__20634;
    wire N__20629;
    wire N__20610;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20604;
    wire N__20603;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20595;
    wire N__20594;
    wire N__20591;
    wire N__20588;
    wire N__20585;
    wire N__20582;
    wire N__20579;
    wire N__20578;
    wire N__20577;
    wire N__20574;
    wire N__20573;
    wire N__20572;
    wire N__20571;
    wire N__20570;
    wire N__20565;
    wire N__20558;
    wire N__20553;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20508;
    wire N__20507;
    wire N__20506;
    wire N__20503;
    wire N__20500;
    wire N__20499;
    wire N__20498;
    wire N__20497;
    wire N__20496;
    wire N__20493;
    wire N__20492;
    wire N__20491;
    wire N__20490;
    wire N__20489;
    wire N__20488;
    wire N__20483;
    wire N__20478;
    wire N__20473;
    wire N__20472;
    wire N__20471;
    wire N__20468;
    wire N__20465;
    wire N__20462;
    wire N__20459;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20440;
    wire N__20437;
    wire N__20432;
    wire N__20429;
    wire N__20428;
    wire N__20427;
    wire N__20426;
    wire N__20423;
    wire N__20418;
    wire N__20411;
    wire N__20406;
    wire N__20399;
    wire N__20388;
    wire N__20387;
    wire N__20386;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20376;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20363;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20336;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20320;
    wire N__20317;
    wire N__20304;
    wire N__20303;
    wire N__20302;
    wire N__20299;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20273;
    wire N__20270;
    wire N__20265;
    wire N__20264;
    wire N__20263;
    wire N__20258;
    wire N__20255;
    wire N__20254;
    wire N__20251;
    wire N__20250;
    wire N__20247;
    wire N__20246;
    wire N__20241;
    wire N__20234;
    wire N__20229;
    wire N__20224;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20184;
    wire N__20169;
    wire N__20168;
    wire N__20167;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20161;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20156;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20125;
    wire N__20122;
    wire N__20119;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20098;
    wire N__20091;
    wire N__20084;
    wire N__20079;
    wire N__20074;
    wire N__20065;
    wire N__20058;
    wire N__20057;
    wire N__20056;
    wire N__20053;
    wire N__20052;
    wire N__20049;
    wire N__20048;
    wire N__20045;
    wire N__20042;
    wire N__20039;
    wire N__20038;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20013;
    wire N__20012;
    wire N__20007;
    wire N__20004;
    wire N__20003;
    wire N__20000;
    wire N__19993;
    wire N__19988;
    wire N__19983;
    wire N__19978;
    wire N__19975;
    wire N__19970;
    wire N__19967;
    wire N__19956;
    wire N__19955;
    wire N__19952;
    wire N__19951;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19937;
    wire N__19934;
    wire N__19933;
    wire N__19930;
    wire N__19929;
    wire N__19928;
    wire N__19927;
    wire N__19926;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19897;
    wire N__19892;
    wire N__19889;
    wire N__19888;
    wire N__19885;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19873;
    wire N__19872;
    wire N__19869;
    wire N__19864;
    wire N__19861;
    wire N__19858;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19839;
    wire N__19832;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19811;
    wire N__19810;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19795;
    wire N__19794;
    wire N__19793;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19781;
    wire N__19780;
    wire N__19779;
    wire N__19778;
    wire N__19775;
    wire N__19774;
    wire N__19771;
    wire N__19766;
    wire N__19763;
    wire N__19758;
    wire N__19757;
    wire N__19756;
    wire N__19755;
    wire N__19750;
    wire N__19745;
    wire N__19744;
    wire N__19743;
    wire N__19740;
    wire N__19739;
    wire N__19736;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19713;
    wire N__19708;
    wire N__19705;
    wire N__19702;
    wire N__19695;
    wire N__19680;
    wire N__19677;
    wire N__19676;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19666;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19655;
    wire N__19654;
    wire N__19651;
    wire N__19650;
    wire N__19649;
    wire N__19648;
    wire N__19647;
    wire N__19646;
    wire N__19645;
    wire N__19642;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19590;
    wire N__19585;
    wire N__19578;
    wire N__19569;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19499;
    wire N__19498;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19421;
    wire N__19420;
    wire N__19419;
    wire N__19418;
    wire N__19417;
    wire N__19414;
    wire N__19409;
    wire N__19408;
    wire N__19407;
    wire N__19404;
    wire N__19403;
    wire N__19402;
    wire N__19397;
    wire N__19396;
    wire N__19395;
    wire N__19390;
    wire N__19385;
    wire N__19382;
    wire N__19377;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19362;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19319;
    wire N__19318;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19314;
    wire N__19313;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19289;
    wire N__19288;
    wire N__19287;
    wire N__19286;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19282;
    wire N__19279;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19241;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19236;
    wire N__19235;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19231;
    wire N__19230;
    wire N__19229;
    wire N__19228;
    wire N__19227;
    wire N__19226;
    wire N__19225;
    wire N__19224;
    wire N__19223;
    wire N__19222;
    wire N__19221;
    wire N__19220;
    wire N__19219;
    wire N__19218;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19214;
    wire N__19213;
    wire N__19212;
    wire N__19211;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19207;
    wire N__19206;
    wire N__19205;
    wire N__19204;
    wire N__19203;
    wire N__19202;
    wire N__19201;
    wire N__19200;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19178;
    wire N__19177;
    wire N__19176;
    wire N__19175;
    wire N__19174;
    wire N__19173;
    wire N__19172;
    wire N__19171;
    wire N__19170;
    wire N__19169;
    wire N__19168;
    wire N__19167;
    wire N__19166;
    wire N__19163;
    wire N__19160;
    wire N__19023;
    wire N__19020;
    wire N__19017;
    wire N__19014;
    wire N__19011;
    wire N__19010;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18999;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18987;
    wire N__18986;
    wire N__18983;
    wire N__18980;
    wire N__18977;
    wire N__18972;
    wire N__18969;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18945;
    wire N__18944;
    wire N__18943;
    wire N__18942;
    wire N__18941;
    wire N__18940;
    wire N__18937;
    wire N__18932;
    wire N__18927;
    wire N__18924;
    wire N__18917;
    wire N__18912;
    wire N__18911;
    wire N__18910;
    wire N__18905;
    wire N__18902;
    wire N__18901;
    wire N__18900;
    wire N__18899;
    wire N__18896;
    wire N__18893;
    wire N__18886;
    wire N__18879;
    wire N__18876;
    wire N__18875;
    wire N__18874;
    wire N__18869;
    wire N__18868;
    wire N__18867;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18855;
    wire N__18854;
    wire N__18853;
    wire N__18852;
    wire N__18851;
    wire N__18850;
    wire N__18847;
    wire N__18846;
    wire N__18843;
    wire N__18838;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18791;
    wire N__18790;
    wire N__18789;
    wire N__18788;
    wire N__18787;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18772;
    wire N__18767;
    wire N__18756;
    wire N__18753;
    wire N__18752;
    wire N__18751;
    wire N__18750;
    wire N__18749;
    wire N__18748;
    wire N__18747;
    wire N__18744;
    wire N__18739;
    wire N__18738;
    wire N__18735;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18720;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18710;
    wire N__18703;
    wire N__18698;
    wire N__18695;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18650;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18633;
    wire N__18632;
    wire N__18629;
    wire N__18628;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18542;
    wire N__18539;
    wire N__18536;
    wire N__18533;
    wire N__18530;
    wire N__18527;
    wire N__18522;
    wire N__18521;
    wire N__18516;
    wire N__18515;
    wire N__18512;
    wire N__18509;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18494;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18477;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18461;
    wire N__18458;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18428;
    wire N__18425;
    wire N__18424;
    wire N__18423;
    wire N__18420;
    wire N__18419;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18391;
    wire N__18384;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18380;
    wire N__18379;
    wire N__18376;
    wire N__18375;
    wire N__18370;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18354;
    wire N__18353;
    wire N__18348;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18315;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18303;
    wire N__18302;
    wire N__18299;
    wire N__18298;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18287;
    wire N__18286;
    wire N__18283;
    wire N__18278;
    wire N__18271;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18257;
    wire N__18254;
    wire N__18253;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18238;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18212;
    wire N__18209;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18176;
    wire N__18175;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18158;
    wire N__18155;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18134;
    wire N__18133;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18119;
    wire N__18116;
    wire N__18113;
    wire N__18108;
    wire N__18105;
    wire N__18104;
    wire N__18103;
    wire N__18098;
    wire N__18095;
    wire N__18090;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18078;
    wire N__18077;
    wire N__18072;
    wire N__18069;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18041;
    wire N__18036;
    wire N__18035;
    wire N__18034;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18006;
    wire N__18003;
    wire N__18002;
    wire N__17999;
    wire N__17998;
    wire N__17995;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17964;
    wire N__17961;
    wire N__17960;
    wire N__17957;
    wire N__17956;
    wire N__17953;
    wire N__17952;
    wire N__17951;
    wire N__17950;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17940;
    wire N__17937;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17898;
    wire N__17897;
    wire N__17896;
    wire N__17895;
    wire N__17892;
    wire N__17885;
    wire N__17882;
    wire N__17877;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17859;
    wire N__17856;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17827;
    wire N__17826;
    wire N__17825;
    wire N__17824;
    wire N__17821;
    wire N__17820;
    wire N__17819;
    wire N__17816;
    wire N__17815;
    wire N__17814;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17802;
    wire N__17799;
    wire N__17794;
    wire N__17791;
    wire N__17784;
    wire N__17769;
    wire N__17768;
    wire N__17767;
    wire N__17764;
    wire N__17763;
    wire N__17762;
    wire N__17761;
    wire N__17758;
    wire N__17757;
    wire N__17756;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17742;
    wire N__17739;
    wire N__17738;
    wire N__17737;
    wire N__17736;
    wire N__17731;
    wire N__17728;
    wire N__17719;
    wire N__17712;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17669;
    wire N__17666;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17651;
    wire N__17650;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17633;
    wire N__17632;
    wire N__17631;
    wire N__17630;
    wire N__17629;
    wire N__17628;
    wire N__17625;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17566;
    wire N__17561;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17544;
    wire N__17543;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17512;
    wire N__17505;
    wire N__17504;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17493;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17476;
    wire N__17473;
    wire N__17466;
    wire N__17465;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17436;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17421;
    wire N__17418;
    wire N__17413;
    wire N__17410;
    wire N__17403;
    wire N__17402;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17396;
    wire N__17395;
    wire N__17392;
    wire N__17391;
    wire N__17388;
    wire N__17387;
    wire N__17384;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17357;
    wire N__17354;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17337;
    wire N__17334;
    wire N__17329;
    wire N__17326;
    wire N__17319;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17308;
    wire N__17303;
    wire N__17300;
    wire N__17295;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17284;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17265;
    wire N__17264;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17237;
    wire N__17232;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17207;
    wire N__17206;
    wire N__17205;
    wire N__17204;
    wire N__17203;
    wire N__17198;
    wire N__17197;
    wire N__17192;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17172;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17129;
    wire N__17128;
    wire N__17127;
    wire N__17124;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17096;
    wire N__17091;
    wire N__17088;
    wire N__17087;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17076;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17061;
    wire N__17052;
    wire N__17051;
    wire N__17050;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17039;
    wire N__17036;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17013;
    wire N__17004;
    wire N__17003;
    wire N__17002;
    wire N__16997;
    wire N__16996;
    wire N__16993;
    wire N__16992;
    wire N__16991;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16978;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16956;
    wire N__16955;
    wire N__16954;
    wire N__16953;
    wire N__16946;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16908;
    wire N__16905;
    wire N__16904;
    wire N__16901;
    wire N__16900;
    wire N__16899;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16879;
    wire N__16876;
    wire N__16867;
    wire N__16864;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16844;
    wire N__16843;
    wire N__16842;
    wire N__16835;
    wire N__16832;
    wire N__16829;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16792;
    wire N__16785;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16774;
    wire N__16769;
    wire N__16766;
    wire N__16761;
    wire N__16752;
    wire N__16751;
    wire N__16750;
    wire N__16747;
    wire N__16746;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16732;
    wire N__16731;
    wire N__16726;
    wire N__16721;
    wire N__16720;
    wire N__16717;
    wire N__16714;
    wire N__16711;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16696;
    wire N__16691;
    wire N__16680;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16652;
    wire N__16651;
    wire N__16646;
    wire N__16643;
    wire N__16638;
    wire N__16635;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16627;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16613;
    wire N__16610;
    wire N__16605;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16535;
    wire N__16534;
    wire N__16533;
    wire N__16532;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16520;
    wire N__16519;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16485;
    wire N__16484;
    wire N__16481;
    wire N__16480;
    wire N__16479;
    wire N__16470;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16448;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16433;
    wire N__16432;
    wire N__16429;
    wire N__16424;
    wire N__16423;
    wire N__16422;
    wire N__16417;
    wire N__16412;
    wire N__16407;
    wire N__16406;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16379;
    wire N__16378;
    wire N__16377;
    wire N__16376;
    wire N__16373;
    wire N__16368;
    wire N__16367;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16339;
    wire N__16332;
    wire N__16325;
    wire N__16322;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16301;
    wire N__16298;
    wire N__16295;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16283;
    wire N__16280;
    wire N__16277;
    wire N__16272;
    wire N__16271;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16260;
    wire N__16259;
    wire N__16258;
    wire N__16253;
    wire N__16250;
    wire N__16247;
    wire N__16242;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16223;
    wire N__16220;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16178;
    wire N__16177;
    wire N__16176;
    wire N__16173;
    wire N__16166;
    wire N__16161;
    wire N__16160;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16145;
    wire N__16142;
    wire N__16139;
    wire N__16136;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16115;
    wire N__16114;
    wire N__16107;
    wire N__16106;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16091;
    wire N__16088;
    wire N__16083;
    wire N__16082;
    wire N__16081;
    wire N__16074;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16044;
    wire N__16043;
    wire N__16040;
    wire N__16039;
    wire N__16036;
    wire N__16035;
    wire N__16034;
    wire N__16031;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__15999;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15993;
    wire N__15990;
    wire N__15987;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15977;
    wire N__15974;
    wire N__15971;
    wire N__15960;
    wire N__15959;
    wire N__15958;
    wire N__15957;
    wire N__15956;
    wire N__15955;
    wire N__15942;
    wire N__15941;
    wire N__15938;
    wire N__15935;
    wire N__15932;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15903;
    wire N__15902;
    wire N__15901;
    wire N__15898;
    wire N__15897;
    wire N__15894;
    wire N__15887;
    wire N__15884;
    wire N__15881;
    wire N__15878;
    wire N__15873;
    wire N__15872;
    wire N__15871;
    wire N__15870;
    wire N__15869;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15832;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15820;
    wire N__15817;
    wire N__15810;
    wire N__15807;
    wire N__15806;
    wire N__15803;
    wire N__15802;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15779;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15752;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15744;
    wire N__15741;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15729;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15708;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15653;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15627;
    wire N__15622;
    wire N__15619;
    wire N__15618;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15603;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15584;
    wire N__15583;
    wire N__15582;
    wire N__15579;
    wire N__15578;
    wire N__15575;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15538;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15516;
    wire N__15513;
    wire N__15512;
    wire N__15509;
    wire N__15506;
    wire N__15501;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15493;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15477;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15469;
    wire N__15468;
    wire N__15467;
    wire N__15462;
    wire N__15455;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15434;
    wire N__15433;
    wire N__15432;
    wire N__15431;
    wire N__15430;
    wire N__15427;
    wire N__15426;
    wire N__15423;
    wire N__15414;
    wire N__15413;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15387;
    wire N__15386;
    wire N__15385;
    wire N__15382;
    wire N__15381;
    wire N__15380;
    wire N__15379;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15364;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15342;
    wire N__15341;
    wire N__15340;
    wire N__15339;
    wire N__15338;
    wire N__15335;
    wire N__15332;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15287;
    wire N__15286;
    wire N__15283;
    wire N__15282;
    wire N__15277;
    wire N__15272;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15260;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15252;
    wire N__15247;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15228;
    wire N__15227;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15219;
    wire N__15218;
    wire N__15215;
    wire N__15208;
    wire N__15203;
    wire N__15198;
    wire N__15197;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15189;
    wire N__15188;
    wire N__15185;
    wire N__15184;
    wire N__15179;
    wire N__15176;
    wire N__15171;
    wire N__15168;
    wire N__15163;
    wire N__15158;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15137;
    wire N__15136;
    wire N__15133;
    wire N__15130;
    wire N__15127;
    wire N__15124;
    wire N__15119;
    wire N__15118;
    wire N__15113;
    wire N__15110;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15098;
    wire N__15097;
    wire N__15094;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15062;
    wire N__15061;
    wire N__15060;
    wire N__15057;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15036;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15006;
    wire N__15005;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14965;
    wire N__14960;
    wire N__14957;
    wire N__14952;
    wire N__14949;
    wire N__14944;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14913;
    wire N__14910;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14891;
    wire N__14888;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14801;
    wire N__14800;
    wire N__14799;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14783;
    wire N__14782;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14764;
    wire N__14759;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14738;
    wire N__14735;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14717;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14691;
    wire N__14688;
    wire N__14681;
    wire N__14678;
    wire N__14673;
    wire N__14670;
    wire N__14667;
    wire N__14664;
    wire N__14661;
    wire N__14660;
    wire N__14655;
    wire N__14654;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14615;
    wire N__14614;
    wire N__14611;
    wire N__14606;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14582;
    wire N__14581;
    wire N__14580;
    wire N__14573;
    wire N__14572;
    wire N__14571;
    wire N__14570;
    wire N__14569;
    wire N__14568;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14562;
    wire N__14561;
    wire N__14558;
    wire N__14555;
    wire N__14548;
    wire N__14539;
    wire N__14536;
    wire N__14531;
    wire N__14526;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14489;
    wire N__14488;
    wire N__14487;
    wire N__14484;
    wire N__14483;
    wire N__14482;
    wire N__14481;
    wire N__14480;
    wire N__14477;
    wire N__14476;
    wire N__14473;
    wire N__14472;
    wire N__14471;
    wire N__14466;
    wire N__14459;
    wire N__14458;
    wire N__14457;
    wire N__14456;
    wire N__14455;
    wire N__14454;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14442;
    wire N__14441;
    wire N__14436;
    wire N__14433;
    wire N__14430;
    wire N__14425;
    wire N__14422;
    wire N__14415;
    wire N__14408;
    wire N__14407;
    wire N__14404;
    wire N__14399;
    wire N__14394;
    wire N__14391;
    wire N__14386;
    wire N__14383;
    wire N__14376;
    wire N__14367;
    wire N__14366;
    wire N__14365;
    wire N__14364;
    wire N__14363;
    wire N__14362;
    wire N__14361;
    wire N__14358;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14340;
    wire N__14337;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14324;
    wire N__14321;
    wire N__14316;
    wire N__14313;
    wire N__14312;
    wire N__14311;
    wire N__14310;
    wire N__14303;
    wire N__14298;
    wire N__14297;
    wire N__14292;
    wire N__14287;
    wire N__14284;
    wire N__14277;
    wire N__14272;
    wire N__14269;
    wire N__14264;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14234;
    wire N__14233;
    wire N__14232;
    wire N__14231;
    wire N__14230;
    wire N__14229;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14199;
    wire N__14196;
    wire N__14191;
    wire N__14184;
    wire N__14181;
    wire N__14180;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14163;
    wire N__14160;
    wire N__14159;
    wire N__14156;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14139;
    wire N__14136;
    wire N__14135;
    wire N__14134;
    wire N__14133;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14125;
    wire N__14124;
    wire N__14121;
    wire N__14116;
    wire N__14111;
    wire N__14108;
    wire N__14103;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14077;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14063;
    wire N__14062;
    wire N__14061;
    wire N__14060;
    wire N__14059;
    wire N__14052;
    wire N__14049;
    wire N__14038;
    wire N__14031;
    wire N__14030;
    wire N__14027;
    wire N__14024;
    wire N__14023;
    wire N__14020;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__13998;
    wire N__13997;
    wire N__13994;
    wire N__13991;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13980;
    wire N__13977;
    wire N__13972;
    wire N__13969;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13955;
    wire N__13954;
    wire N__13953;
    wire N__13950;
    wire N__13945;
    wire N__13942;
    wire N__13937;
    wire N__13932;
    wire N__13929;
    wire N__13928;
    wire N__13925;
    wire N__13922;
    wire N__13919;
    wire N__13918;
    wire N__13917;
    wire N__13916;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13906;
    wire N__13901;
    wire N__13898;
    wire N__13893;
    wire N__13888;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13861;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13849;
    wire N__13846;
    wire N__13839;
    wire N__13836;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13797;
    wire N__13794;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13779;
    wire N__13778;
    wire N__13777;
    wire N__13776;
    wire N__13775;
    wire N__13774;
    wire N__13773;
    wire N__13766;
    wire N__13757;
    wire N__13752;
    wire N__13751;
    wire N__13750;
    wire N__13749;
    wire N__13748;
    wire N__13747;
    wire N__13746;
    wire N__13743;
    wire N__13738;
    wire N__13729;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13718;
    wire N__13717;
    wire N__13716;
    wire N__13709;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13679;
    wire N__13678;
    wire N__13675;
    wire N__13672;
    wire N__13671;
    wire N__13670;
    wire N__13659;
    wire N__13658;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13643;
    wire N__13638;
    wire N__13637;
    wire N__13636;
    wire N__13635;
    wire N__13634;
    wire N__13623;
    wire N__13622;
    wire N__13621;
    wire N__13618;
    wire N__13613;
    wire N__13608;
    wire N__13607;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13601;
    wire N__13600;
    wire N__13599;
    wire N__13592;
    wire N__13583;
    wire N__13578;
    wire N__13577;
    wire N__13576;
    wire N__13575;
    wire N__13574;
    wire N__13573;
    wire N__13572;
    wire N__13565;
    wire N__13556;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13538;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13530;
    wire N__13521;
    wire N__13514;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13497;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13449;
    wire N__13440;
    wire N__13439;
    wire N__13438;
    wire N__13437;
    wire N__13434;
    wire N__13427;
    wire N__13422;
    wire N__13421;
    wire N__13420;
    wire N__13419;
    wire N__13416;
    wire N__13415;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13405;
    wire N__13404;
    wire N__13393;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13353;
    wire N__13350;
    wire N__13347;
    wire N__13344;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13338;
    wire N__13331;
    wire N__13328;
    wire N__13323;
    wire N__13320;
    wire N__13317;
    wire N__13316;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13304;
    wire N__13299;
    wire N__13296;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13281;
    wire N__13280;
    wire N__13275;
    wire N__13272;
    wire N__13269;
    wire N__13266;
    wire N__13263;
    wire N__13260;
    wire N__13257;
    wire N__13256;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13212;
    wire N__13207;
    wire N__13202;
    wire N__13201;
    wire N__13200;
    wire N__13199;
    wire N__13194;
    wire N__13189;
    wire N__13188;
    wire N__13187;
    wire N__13186;
    wire N__13185;
    wire N__13184;
    wire N__13183;
    wire N__13182;
    wire N__13181;
    wire N__13180;
    wire N__13177;
    wire N__13172;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13141;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13086;
    wire N__13085;
    wire N__13084;
    wire N__13081;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13075;
    wire N__13070;
    wire N__13069;
    wire N__13068;
    wire N__13065;
    wire N__13056;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13039;
    wire N__13036;
    wire N__13031;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13011;
    wire N__13010;
    wire N__13009;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12995;
    wire N__12990;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12982;
    wire N__12977;
    wire N__12972;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12963;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12927;
    wire N__12926;
    wire N__12925;
    wire N__12922;
    wire N__12921;
    wire N__12916;
    wire N__12913;
    wire N__12912;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12897;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12881;
    wire N__12878;
    wire N__12877;
    wire N__12874;
    wire N__12873;
    wire N__12870;
    wire N__12865;
    wire N__12862;
    wire N__12857;
    wire N__12852;
    wire N__12851;
    wire N__12850;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12842;
    wire N__12839;
    wire N__12834;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12816;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12766;
    wire N__12761;
    wire N__12758;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12725;
    wire N__12722;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12702;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12668;
    wire N__12667;
    wire N__12666;
    wire N__12657;
    wire N__12654;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12648;
    wire N__12641;
    wire N__12636;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12605;
    wire N__12604;
    wire N__12601;
    wire N__12596;
    wire N__12593;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12581;
    wire N__12580;
    wire N__12579;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12571;
    wire N__12568;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12560;
    wire N__12559;
    wire N__12558;
    wire N__12551;
    wire N__12548;
    wire N__12547;
    wire N__12544;
    wire N__12541;
    wire N__12538;
    wire N__12531;
    wire N__12528;
    wire N__12525;
    wire N__12520;
    wire N__12515;
    wire N__12504;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12479;
    wire N__12476;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12436;
    wire N__12435;
    wire N__12424;
    wire N__12419;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12377;
    wire N__12376;
    wire N__12375;
    wire N__12374;
    wire N__12373;
    wire N__12370;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12360;
    wire N__12359;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12347;
    wire N__12344;
    wire N__12341;
    wire N__12338;
    wire N__12333;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12263;
    wire N__12262;
    wire N__12259;
    wire N__12258;
    wire N__12257;
    wire N__12254;
    wire N__12253;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12234;
    wire N__12225;
    wire N__12222;
    wire N__12219;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12195;
    wire N__12194;
    wire N__12193;
    wire N__12192;
    wire N__12191;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12168;
    wire N__12165;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12095;
    wire N__12092;
    wire N__12091;
    wire N__12090;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12075;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12059;
    wire N__12058;
    wire N__12057;
    wire N__12054;
    wire N__12053;
    wire N__12048;
    wire N__12045;
    wire N__12040;
    wire N__12037;
    wire N__12030;
    wire N__12027;
    wire N__12026;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11970;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11958;
    wire N__11957;
    wire N__11954;
    wire N__11951;
    wire N__11948;
    wire N__11945;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11935;
    wire N__11930;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11915;
    wire N__11912;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11887;
    wire N__11884;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11865;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11851;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11828;
    wire N__11827;
    wire N__11826;
    wire N__11825;
    wire N__11824;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11820;
    wire N__11819;
    wire N__11814;
    wire N__11811;
    wire N__11804;
    wire N__11797;
    wire N__11796;
    wire N__11791;
    wire N__11782;
    wire N__11779;
    wire N__11772;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11764;
    wire N__11763;
    wire N__11760;
    wire N__11753;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11734;
    wire N__11731;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11711;
    wire N__11708;
    wire N__11707;
    wire N__11706;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11692;
    wire N__11685;
    wire N__11682;
    wire N__11681;
    wire N__11680;
    wire N__11679;
    wire N__11678;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11664;
    wire N__11655;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11638;
    wire N__11631;
    wire N__11628;
    wire N__11627;
    wire N__11626;
    wire N__11625;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11611;
    wire N__11604;
    wire N__11601;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11544;
    wire N__11543;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11533;
    wire N__11528;
    wire N__11523;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11517;
    wire N__11516;
    wire N__11511;
    wire N__11504;
    wire N__11499;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11491;
    wire N__11484;
    wire N__11481;
    wire N__11480;
    wire N__11479;
    wire N__11476;
    wire N__11475;
    wire N__11472;
    wire N__11467;
    wire N__11464;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11436;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11321;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11304;
    wire N__11303;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11276;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11259;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11255;
    wire N__11254;
    wire N__11253;
    wire N__11252;
    wire N__11251;
    wire N__11250;
    wire N__11241;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11225;
    wire N__11220;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11207;
    wire N__11206;
    wire N__11205;
    wire N__11204;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11186;
    wire N__11179;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11132;
    wire N__11131;
    wire N__11130;
    wire N__11121;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11115;
    wire N__11108;
    wire N__11103;
    wire N__11102;
    wire N__11101;
    wire N__11100;
    wire N__11091;
    wire N__11090;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11079;
    wire N__11076;
    wire N__11069;
    wire N__11064;
    wire N__11063;
    wire N__11062;
    wire N__11061;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11050;
    wire N__11049;
    wire N__11046;
    wire N__11037;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10979;
    wire N__10978;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10970;
    wire N__10965;
    wire N__10960;
    wire N__10957;
    wire N__10950;
    wire N__10947;
    wire N__10944;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10925;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10887;
    wire N__10884;
    wire N__10881;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10857;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10844;
    wire N__10843;
    wire N__10832;
    wire N__10831;
    wire N__10830;
    wire N__10829;
    wire N__10828;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10809;
    wire N__10800;
    wire N__10799;
    wire N__10798;
    wire N__10797;
    wire N__10794;
    wire N__10793;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10787;
    wire N__10784;
    wire N__10783;
    wire N__10780;
    wire N__10771;
    wire N__10764;
    wire N__10761;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10706;
    wire N__10701;
    wire N__10700;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10692;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10662;
    wire N__10653;
    wire N__10650;
    wire N__10649;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10638;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10612;
    wire N__10605;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10592;
    wire N__10587;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10579;
    wire N__10574;
    wire N__10573;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10552;
    wire N__10539;
    wire N__10536;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10526;
    wire N__10525;
    wire N__10524;
    wire N__10521;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10513;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10485;
    wire N__10484;
    wire N__10483;
    wire N__10482;
    wire N__10481;
    wire N__10480;
    wire N__10479;
    wire N__10478;
    wire N__10477;
    wire N__10476;
    wire N__10473;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10437;
    wire N__10436;
    wire N__10435;
    wire N__10428;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10422;
    wire N__10417;
    wire N__10414;
    wire N__10409;
    wire N__10404;
    wire N__10403;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10392;
    wire N__10391;
    wire N__10384;
    wire N__10381;
    wire N__10380;
    wire N__10379;
    wire N__10378;
    wire N__10377;
    wire N__10376;
    wire N__10375;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10357;
    wire N__10348;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10330;
    wire N__10329;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10317;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10303;
    wire N__10298;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10273;
    wire N__10270;
    wire N__10265;
    wire N__10258;
    wire N__10255;
    wire N__10250;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10218;
    wire N__10215;
    wire N__10212;
    wire N__10209;
    wire N__10206;
    wire N__10203;
    wire N__10200;
    wire N__10197;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10122;
    wire N__10121;
    wire N__10118;
    wire N__10117;
    wire N__10116;
    wire N__10115;
    wire N__10114;
    wire N__10111;
    wire N__10108;
    wire N__10103;
    wire N__10098;
    wire N__10095;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10077;
    wire N__10074;
    wire N__10071;
    wire N__10062;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10036;
    wire N__10029;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10005;
    wire N__10004;
    wire N__10003;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9846;
    wire N__9845;
    wire N__9840;
    wire N__9837;
    wire N__9832;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9798;
    wire N__9797;
    wire N__9796;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9784;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9759;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9741;
    wire N__9738;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9701;
    wire N__9694;
    wire N__9691;
    wire N__9686;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9668;
    wire N__9663;
    wire N__9662;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9650;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9638;
    wire N__9637;
    wire N__9636;
    wire N__9633;
    wire N__9632;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9585;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9575;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9561;
    wire N__9556;
    wire N__9547;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9489;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9476;
    wire N__9475;
    wire N__9474;
    wire N__9471;
    wire N__9470;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9405;
    wire N__9402;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9389;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9381;
    wire N__9380;
    wire N__9377;
    wire N__9376;
    wire N__9375;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9359;
    wire N__9354;
    wire N__9345;
    wire N__9342;
    wire N__9341;
    wire N__9340;
    wire N__9339;
    wire N__9338;
    wire N__9335;
    wire N__9328;
    wire N__9325;
    wire N__9318;
    wire N__9317;
    wire N__9316;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9304;
    wire N__9299;
    wire N__9294;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9270;
    wire N__9269;
    wire N__9268;
    wire N__9267;
    wire N__9264;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9243;
    wire N__9242;
    wire N__9241;
    wire N__9236;
    wire N__9233;
    wire N__9228;
    wire N__9225;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9216;
    wire N__9211;
    wire N__9208;
    wire N__9203;
    wire N__9198;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9186;
    wire N__9185;
    wire N__9184;
    wire N__9181;
    wire N__9180;
    wire N__9179;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9156;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9144;
    wire N__9143;
    wire N__9140;
    wire N__9139;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9123;
    wire N__9122;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9095;
    wire N__9090;
    wire N__9087;
    wire N__9086;
    wire N__9085;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9067;
    wire N__9064;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9041;
    wire N__9040;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9034;
    wire N__9023;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9005;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8995;
    wire N__8992;
    wire N__8987;
    wire N__8984;
    wire N__8979;
    wire N__8978;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8905;
    wire N__8900;
    wire N__8899;
    wire N__8898;
    wire N__8893;
    wire N__8890;
    wire N__8889;
    wire N__8886;
    wire N__8885;
    wire N__8884;
    wire N__8883;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8871;
    wire N__8862;
    wire N__8853;
    wire N__8852;
    wire N__8851;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8834;
    wire N__8833;
    wire N__8832;
    wire N__8825;
    wire N__8822;
    wire N__8817;
    wire N__8816;
    wire N__8815;
    wire N__8814;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8806;
    wire N__8805;
    wire N__8804;
    wire N__8803;
    wire N__8802;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8763;
    wire N__8758;
    wire N__8745;
    wire N__8742;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8730;
    wire N__8729;
    wire N__8728;
    wire N__8727;
    wire N__8726;
    wire N__8725;
    wire N__8724;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8693;
    wire N__8684;
    wire N__8681;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8658;
    wire N__8657;
    wire N__8654;
    wire N__8653;
    wire N__8650;
    wire N__8643;
    wire N__8640;
    wire N__8639;
    wire N__8638;
    wire N__8633;
    wire N__8630;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8612;
    wire N__8611;
    wire N__8608;
    wire N__8607;
    wire N__8606;
    wire N__8605;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8589;
    wire N__8586;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8566;
    wire N__8565;
    wire N__8564;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8538;
    wire N__8535;
    wire N__8534;
    wire N__8533;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8525;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8499;
    wire N__8498;
    wire N__8497;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8485;
    wire N__8480;
    wire N__8475;
    wire N__8472;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8460;
    wire N__8455;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8391;
    wire N__8388;
    wire N__8385;
    wire N__8382;
    wire N__8381;
    wire N__8380;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8368;
    wire N__8361;
    wire N__8358;
    wire N__8357;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8339;
    wire N__8334;
    wire N__8331;
    wire N__8328;
    wire N__8325;
    wire N__8324;
    wire N__8323;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8295;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8252;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8235;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8218;
    wire N__8217;
    wire N__8208;
    wire N__8205;
    wire N__8204;
    wire N__8203;
    wire N__8200;
    wire N__8195;
    wire N__8192;
    wire N__8187;
    wire N__8184;
    wire N__8183;
    wire N__8182;
    wire N__8181;
    wire N__8178;
    wire N__8175;
    wire N__8170;
    wire N__8167;
    wire N__8160;
    wire N__8159;
    wire N__8158;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8140;
    wire N__8133;
    wire N__8132;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8090;
    wire N__8089;
    wire N__8088;
    wire N__8085;
    wire N__8078;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8064;
    wire N__8063;
    wire N__8062;
    wire N__8061;
    wire N__8060;
    wire N__8059;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8030;
    wire N__8025;
    wire N__8022;
    wire N__8021;
    wire N__8020;
    wire N__8013;
    wire N__8010;
    wire N__8009;
    wire N__8008;
    wire N__8005;
    wire N__8000;
    wire N__7995;
    wire N__7992;
    wire N__7991;
    wire N__7990;
    wire N__7989;
    wire N__7988;
    wire N__7985;
    wire N__7984;
    wire N__7971;
    wire N__7968;
    wire N__7967;
    wire N__7966;
    wire N__7965;
    wire N__7964;
    wire N__7955;
    wire N__7952;
    wire N__7947;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7939;
    wire N__7938;
    wire N__7931;
    wire N__7928;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7918;
    wire N__7917;
    wire N__7916;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7897;
    wire N__7894;
    wire N__7887;
    wire N__7884;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7874;
    wire N__7873;
    wire N__7870;
    wire N__7865;
    wire N__7860;
    wire N__7857;
    wire N__7856;
    wire N__7855;
    wire N__7854;
    wire N__7853;
    wire N__7846;
    wire N__7841;
    wire N__7836;
    wire N__7835;
    wire N__7834;
    wire N__7831;
    wire N__7828;
    wire N__7823;
    wire N__7818;
    wire N__7815;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7768;
    wire N__7765;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire clk_in_c;
    wire VCCG0;
    wire GNDG0;
    wire \uu2.mem0.N_137 ;
    wire \uu2.mem0.N_141 ;
    wire \uu2.bitmap_pmux_u_0_a2_0_cascade_ ;
    wire \uu2.mem0.N_140 ;
    wire \uu2.mem0.N_139 ;
    wire \INVuu2.w_addr_user_1C_net ;
    wire uart_RXD;
    wire \uu0.l_precountZ0Z_1 ;
    wire \uu0.l_precountZ0Z_3 ;
    wire \uu0.un4_l_count_11_cascade_ ;
    wire \uu0.un4_l_count_16_cascade_ ;
    wire \uu0.delay_lineZ0Z_1 ;
    wire \uu0.un4_l_count_0_cascade_ ;
    wire \uu0.delay_lineZ0Z_0 ;
    wire \uu0.un11_l_count_i ;
    wire \uu0.l_precountZ0Z_2 ;
    wire \uu0.un4_l_count_13 ;
    wire \uu0.un55_ci_cascade_ ;
    wire \uu0.l_countZ0Z_0 ;
    wire \uu0.l_countZ0Z_1 ;
    wire \uu0.l_countZ0Z_2 ;
    wire \uu0.l_precountZ0Z_0 ;
    wire \uu0.un4_l_count_14_cascade_ ;
    wire \uu0.un4_l_count_18 ;
    wire \uu0.l_countZ0Z_11 ;
    wire \uu0.un154_ci_9_cascade_ ;
    wire \uu0.l_countZ0Z_10 ;
    wire \uu0.un143_ci_0 ;
    wire \uu0.l_countZ0Z_8 ;
    wire \uu0.un187_ci_1_cascade_ ;
    wire \uu0.un165_ci_0 ;
    wire \uu0.l_countZ0Z_13 ;
    wire \uu0.l_countZ0Z_12 ;
    wire \uu0.un4_l_count_0_8 ;
    wire \uu0.un154_ci_9 ;
    wire \uu0.l_countZ0Z_15 ;
    wire \uu0.un4_l_count_0_8_cascade_ ;
    wire \uu0.l_countZ0Z_14 ;
    wire \uu0.l_countZ0Z_4 ;
    wire \uu0.l_countZ0Z_5 ;
    wire \uu2.N_34_cascade_ ;
    wire \uu2.N_114 ;
    wire \uu2.mem0.w_data_6 ;
    wire \uu2.mem0.N_31_i ;
    wire \uu2.mem0.N_61_cascade_ ;
    wire \uu2.mem0.w_data_1 ;
    wire \uu2.mem0.w_data_4 ;
    wire \uu2.N_922_tz_tz ;
    wire \uu2.bitmap_pmux ;
    wire \uu2.bitmap_pmux_cascade_ ;
    wire \uu2.mem0.w_data_3 ;
    wire \uu2.N_37 ;
    wire \uu2.mem0.N_59 ;
    wire \uu2.mem0.w_data_0 ;
    wire \uu2.un404_ci_cascade_ ;
    wire \uu2.r_addrZ0Z_8 ;
    wire \uu2.vbuf_raddr.un426_ci_3 ;
    wire \uu2.vbuf_raddr.un426_ci_3_cascade_ ;
    wire \uu2.r_addrZ0Z_7 ;
    wire \uu2.vbuf_raddr.un448_ci_0 ;
    wire \uu2.r_addrZ0Z_6 ;
    wire \uu2.r_addrZ0Z_3 ;
    wire \uu2.trig_rd_is_det_0 ;
    wire \INVuu2.w_addr_user_4C_net ;
    wire \uu2.r_addrZ0Z_2 ;
    wire \uu2.r_addrZ0Z_0 ;
    wire \uu2.r_addrZ0Z_1 ;
    wire \uu2.r_addrZ0Z_4 ;
    wire \uu2.un404_ci ;
    wire \uu2.r_addrZ0Z_5 ;
    wire \uu0.un66_ci ;
    wire \uu0.un110_ci ;
    wire \uu0.un198_ci_2 ;
    wire \uu0.un110_ci_cascade_ ;
    wire \uu0.l_countZ0Z_16 ;
    wire \uu0.un4_l_count_0 ;
    wire \uu0.un220_ci_cascade_ ;
    wire \uu0.l_countZ0Z_18 ;
    wire \uu0.un11_l_count_i_g ;
    wire \uu0.l_countZ0Z_9 ;
    wire \uu0.l_countZ0Z_7 ;
    wire \uu0.l_countZ0Z_17 ;
    wire \uu0.l_countZ0Z_3 ;
    wire \uu0.un4_l_count_12 ;
    wire \uu2.un1_l_count_2_2_cascade_ ;
    wire \uu2.un1_l_count_2_0_cascade_ ;
    wire \uu2.un1_l_count_1_3 ;
    wire \uu2.un1_l_count_2_0 ;
    wire \uu2.l_countZ0Z_9 ;
    wire \uu2.un1_l_count_1_2_0 ;
    wire \uu2.l_countZ0Z_1 ;
    wire \uu2.l_countZ0Z_0 ;
    wire \uu2.l_countZ0Z_3 ;
    wire \uu2.un306_ci ;
    wire \uu2.l_countZ0Z_7 ;
    wire \uu2.un306_ci_cascade_ ;
    wire \uu2.l_countZ0Z_6 ;
    wire \uu2.un284_ci ;
    wire \uu2.l_countZ0Z_2 ;
    wire \uu2.un350_ci ;
    wire \uu2.l_countZ0Z_8 ;
    wire \uu0.un88_ci_3 ;
    wire \uu0.l_countZ0Z_6 ;
    wire \uu0.un99_ci_0 ;
    wire \uu2.w_data_0_a2_0_6_cascade_ ;
    wire \uu2.w_data_0_a2_2_6 ;
    wire \INVuu2.w_addr_displaying_nesr_4C_net ;
    wire \uu2.bitmap_pmux_u_0_a2_0_2_0 ;
    wire \uu2.w_addr_displayingZ0Z_4 ;
    wire \uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_ ;
    wire \INVuu2.w_addr_displaying_fast_2C_net ;
    wire \uu2.w_addr_displaying_fastZ0Z_2 ;
    wire \uu2.bitmapZ0Z_186 ;
    wire \uu2.bitmapZ0Z_58 ;
    wire \INVuu2.bitmap_186C_net ;
    wire \uu2.bitmapZ0Z_93 ;
    wire \uu2.bitmapZ0Z_221 ;
    wire \uu2.bitmap_RNIRETJ1Z0Z_93_cascade_ ;
    wire \uu2.bitmap_pmux_27_ns_1_cascade_ ;
    wire \uu2.N_404 ;
    wire \uu2.mem0.N_135 ;
    wire \uu2.mem0.N_134 ;
    wire \INVuu2.w_addr_displaying_nesr_7C_net ;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_ ;
    wire \uu2.N_32_0 ;
    wire \uu2.mem0.N_133 ;
    wire \uu2.w_addr_userZ0Z_8 ;
    wire \uu2.N_161_cascade_ ;
    wire \INVuu2.w_addr_user_nesr_8C_net ;
    wire \uu2.N_101_cascade_ ;
    wire \uu2.w_addr_userZ0Z_1 ;
    wire \uu2.w_addr_userZ0Z_0 ;
    wire \uu2.N_106_cascade_ ;
    wire \uu2.N_164 ;
    wire \uu2.w_addr_userZ0Z_2 ;
    wire \uu2.w_addr_user_3_i_a2_3_6 ;
    wire \uu2.w_addr_user_3_i_a2_2_6_cascade_ ;
    wire \uu2.N_230 ;
    wire \uu2.w_addr_userZ0Z_3 ;
    wire \uu2.mem0.N_138 ;
    wire oneSecStrb_cascade_;
    wire clk;
    wire \uu2.vram_wr_en_0_iZ0 ;
    wire \uu2.N_102 ;
    wire \uu2.mem0.N_54_i ;
    wire \uu2.r_data_wire_0 ;
    wire \uu2.r_data_wire_1 ;
    wire \uu2.r_data_wire_2 ;
    wire \uu2.r_data_wire_3 ;
    wire \uu2.r_data_wire_4 ;
    wire \uu2.r_data_wire_5 ;
    wire \uu2.r_data_wire_6 ;
    wire \uu2.r_data_wire_7 ;
    wire \INVuu2.r_data_reg_0C_net ;
    wire \uu2.trig_rd_detZ0Z_1 ;
    wire \uu2.trig_rd_detZ0Z_0 ;
    wire \uu2.trig_rd_is_det ;
    wire \uu2.l_countZ0Z_4 ;
    wire \uu2.l_countZ0Z_5 ;
    wire \uu2.vbuf_count.un328_ci_3 ;
    wire bfn_4_11_0_;
    wire \buart.Z_rx.bitcount_cry_0_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_0 ;
    wire \buart.Z_rx.bitcount_cry_1_THRU_CO ;
    wire \buart.Z_rx.bitcount_cry_1 ;
    wire \buart.Z_rx.bitcount_cry_2 ;
    wire \buart.Z_rx.bitcount_cry_3 ;
    wire bfn_4_12_0_;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_2 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_4 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ;
    wire \uu2.bitmapZ0Z_194 ;
    wire \uu2.bitmap_pmux_25_i_m2_am_1_cascade_ ;
    wire \uu2.bitmap_RNIG91I1Z0Z_66 ;
    wire \uu2.bitmapZ0Z_69 ;
    wire \uu2.bitmapZ0Z_66 ;
    wire \uu2.bitmapZ0Z_197 ;
    wire \INVuu2.bitmap_194C_net ;
    wire \uu2.w_addr_displayingZ0Z_2 ;
    wire \uu2.N_34 ;
    wire \uu2.w_addr_displayingZ0Z_3 ;
    wire \uu2.N_47 ;
    wire \uu2.N_38 ;
    wire \uu2.w_addr_displaying_RNI0ES07Z0Z_5 ;
    wire \uu2.N_33 ;
    wire \uu2.w_addr_displayingZ0Z_1 ;
    wire \INVuu2.w_addr_displaying_3_rep1C_net ;
    wire L3_tx_data_rdy;
    wire \uu2.mem0.N_136 ;
    wire \uu2.bitmap_RNIFJI02Z0Z_212 ;
    wire \uu2.N_65 ;
    wire \uu2.bitmap_pmux_u_0_83_0 ;
    wire \uu2.w_addr_displayingZ0Z_5 ;
    wire \uu2.w_addr_displayingZ0Z_6 ;
    wire \uu2.bitmap_pmux_sn_N_42 ;
    wire \uu2.N_112_i ;
    wire \uu2.N_100_cascade_ ;
    wire \uu2.N_921_tz_tz ;
    wire \uu2.bitmap_pmux_sn_N_20 ;
    wire \uu2.N_923_tz_cascade_ ;
    wire \uu2.w_addr_displaying_RNI8ND5GZ0Z_3 ;
    wire \INVuu2.bitmap_314C_net ;
    wire \uu2.bitmapZ0Z_218 ;
    wire \uu2.bitmapZ0Z_90 ;
    wire \uu2.bitmap_pmux_25_i_m2_bm_1 ;
    wire \uu2.w_addr_displaying_fastZ0Z_7 ;
    wire \uu2.bitmap_pmux_21_ns_1_cascade_ ;
    wire \uu2.bitmap_pmux_sn_N_11 ;
    wire \uu2.N_393_cascade_ ;
    wire \uu2.N_397 ;
    wire \uu2.bitmapZ0Z_314 ;
    wire \uu2.N_128 ;
    wire \uu2.N_131 ;
    wire \uu2.un1_l_count_1_0 ;
    wire \Lab_UT.didp.countrce1.q_5_0_cascade_ ;
    wire \Lab_UT.sec2_1 ;
    wire \Lab_UT.sec2_2 ;
    wire \Lab_UT.sec2_3 ;
    wire \uu2.un28_w_addr_user_i_0_a2_0Z0Z_4 ;
    wire \Lab_UT.dispString.un42_dOutP_cascade_ ;
    wire \uu2.un28_w_addr_user_i_0_a2_0Z0Z_0 ;
    wire \Lab_UT.dispString.N_211_cascade_ ;
    wire \Lab_UT.dispString.dOutP_0_iv_0_2 ;
    wire \Lab_UT.dispString.dOutP_0_iv_1_2 ;
    wire \uu2.vram_rd_clk_det_RNI95711Z0Z_1 ;
    wire L3_tx_data_4;
    wire L3_tx_data_2;
    wire \uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_ ;
    wire L3_tx_data_0;
    wire \uu2.un1_w_user_cr_0 ;
    wire L3_tx_data_5;
    wire vbuf_tx_data_0;
    wire \buart.Z_tx.shifterZ0Z_1 ;
    wire \buart.Z_tx.shifterZ0Z_0 ;
    wire o_serial_data_c;
    wire vbuf_tx_data_1;
    wire \buart.Z_tx.shifterZ0Z_2 ;
    wire vbuf_tx_data_2;
    wire \buart.Z_tx.shifterZ0Z_3 ;
    wire vbuf_tx_data_3;
    wire \buart.Z_tx.shifterZ0Z_4 ;
    wire vbuf_tx_data_4;
    wire \buart.Z_tx.shifterZ0Z_5 ;
    wire vbuf_tx_data_5;
    wire \buart.Z_tx.shifterZ0Z_6 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ;
    wire \Lab_UT.dispString.N_191 ;
    wire \buart.Z_tx.bitcount_RNO_0Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_3 ;
    wire \buart.Z_tx.uart_busy_0_0 ;
    wire \buart.Z_rx.hhZ0Z_0 ;
    wire \buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_0 ;
    wire \buart.Z_tx.bitcountZ0Z_2 ;
    wire \buart.Z_tx.bitcountZ0Z_1 ;
    wire \buart.Z_tx.un1_bitcount_c3 ;
    wire \buart.Z_rx.idle_0_cascade_ ;
    wire \buart.Z_rx.idle ;
    wire \buart.Z_rx.bitcount_cry_2_THRU_CO ;
    wire \buart.Z_rx.bitcountZ0Z_3 ;
    wire \buart.Z_rx.bitcountZ0Z_1 ;
    wire \buart.Z_rx.bitcountZ0Z_4 ;
    wire \buart.Z_rx.valid_1_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_2 ;
    wire \buart.Z_rx.N_27_0_i ;
    wire \buart.Z_rx.bitcounte_0_0 ;
    wire \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_1 ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ;
    wire \buart.Z_rx.ser_clk ;
    wire \buart.Z_rx.un1_sample_0 ;
    wire \buart.Z_rx.ser_clk_cascade_ ;
    wire \buart.Z_rx.bitcountZ0Z_0 ;
    wire \buart.Z_rx.sample ;
    wire \buart.Z_rx.startbit ;
    wire \buart.Z_rx.Z_baudgen.counterZ0Z_0 ;
    wire \uu2.bitmapZ0Z_168 ;
    wire \uu2.bitmapZ0Z_75 ;
    wire \uu2.bitmapZ0Z_203 ;
    wire \uu2.bitmapZ0Z_162 ;
    wire \INVuu2.bitmap_168C_net ;
    wire \uu2.bitmapZ0Z_34 ;
    wire \uu2.w_addr_displaying_fastZ0Z_3 ;
    wire \uu2.bitmapZ0Z_290 ;
    wire \uu2.bitmap_pmux_24_bm_1 ;
    wire \uu2.bitmapZ0Z_72 ;
    wire \uu2.bitmapZ0Z_200 ;
    wire \uu2.w_addr_displayingZ0Z_0 ;
    wire \uu2.bitmap_RNI5T9T1Z0Z_72 ;
    wire \INVuu2.bitmap_296C_net ;
    wire \uu2.bitmap_pmux_sn_N_54_mux ;
    wire \uu2.N_237 ;
    wire \uu2.bitmap_pmux_sn_N_15 ;
    wire \uu2.N_395_cascade_ ;
    wire \uu2.N_401 ;
    wire \uu2.bitmapZ0Z_296 ;
    wire \uu2.w_addr_displaying_3_repZ0Z1 ;
    wire \uu2.bitmapZ0Z_40 ;
    wire \uu2.bitmap_pmux_15_i_m2_ns_1 ;
    wire \uu2.N_123 ;
    wire \uu2.w_addr_displayingZ0Z_8 ;
    wire \uu2.bitmapZ0Z_308 ;
    wire \uu2.bitmap_RNIU2ISZ0Z_52 ;
    wire \uu2.bitmapZ0Z_52 ;
    wire \INVuu2.bitmap_308C_net ;
    wire \uu2.w_addr_displayingZ0Z_7 ;
    wire \uu2.bitmapZ0Z_84 ;
    wire \uu2.bitmapZ0Z_87 ;
    wire \uu2.w_addr_displaying_fastZ0Z_0 ;
    wire \uu2.bitmap_pmux_24_am_1 ;
    wire \Lab_UT.min1_1 ;
    wire \Lab_UT.dispString.un46_dOutP_2 ;
    wire \Lab_UT.sec2_0 ;
    wire G_190;
    wire G_190_cascade_;
    wire \Lab_UT.dispString.i21_mux ;
    wire \Lab_UT.dispString.m28_ns_1_cascade_ ;
    wire \Lab_UT.dispString.N_204 ;
    wire \Lab_UT.di_ASones_0 ;
    wire \uu2.w_addr_userZ0Z_6 ;
    wire \uu2.w_addr_userZ0Z_4 ;
    wire \uu2.N_106 ;
    wire \uu2.w_addr_userZ0Z_5 ;
    wire \INVuu2.w_addr_user_nesr_5C_net ;
    wire \uu2.un28_w_addr_user_i_0_0 ;
    wire G_193;
    wire G_193_cascade_;
    wire \Lab_UT.dispString.N_219 ;
    wire \Lab_UT.dispString.N_222_cascade_ ;
    wire L3_tx_data_3;
    wire G_189;
    wire G_189_cascade_;
    wire \Lab_UT.dispString.un42_dOutP ;
    wire L3_tx_data_6;
    wire uu0_sec_clkD;
    wire \Lab_UT.dispString.m44_ns_1 ;
    wire L3_tx_data_1;
    wire \Lab_UT.dispString.m42_ns_1 ;
    wire vbuf_tx_data_6;
    wire \buart.Z_tx.shifterZ0Z_7 ;
    wire vbuf_tx_data_rdy;
    wire vbuf_tx_data_7;
    wire \buart.Z_tx.shifterZ0Z_8 ;
    wire \buart.Z_tx.un1_uart_wr_i_0_i ;
    wire \Lab_UT.dispString.cntZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_0 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_1 ;
    wire bfn_6_10_0_;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_1 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_2 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_3 ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_4 ;
    wire \buart.Z_tx.ser_clk ;
    wire \buart.Z_tx.Z_baudgen.un2_counter_cry_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_5 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_4 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_6 ;
    wire \buart.Z_tx.Z_baudgen.counterZ0Z_3 ;
    wire \buart.Z_tx.Z_baudgen.ser_clk_4 ;
    wire \Lab_UT.dictrl.g1Z0Z_5 ;
    wire \Lab_UT.dictrl.g1_cascade_ ;
    wire \Lab_UT.dictrl.g0_2_3_cascade_ ;
    wire \Lab_UT.dictrl.g0_17_a6_1_7 ;
    wire \Lab_UT.dictrl.g0_17_a6_1Z0Z_6 ;
    wire \Lab_UT.dictrl.g0_17_a6_1_5_cascade_ ;
    wire \Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_ ;
    wire \Lab_UT.dictrl.g0_17_a6_2 ;
    wire \Lab_UT.dictrl.N_19 ;
    wire \Lab_UT.dictrl.g0_17_o6_1Z0Z_5 ;
    wire \Lab_UT.min2_3 ;
    wire \Lab_UT.min1_3 ;
    wire \Lab_UT.min1_2 ;
    wire \Lab_UT.min1_0 ;
    wire \Lab_UT.min2_1 ;
    wire \Lab_UT.min2_0 ;
    wire \Lab_UT.min2_2 ;
    wire \Lab_UT.dispString.N_18_0_cascade_ ;
    wire \Lab_UT.dispString.dOut_RNO_0Z0Z_1 ;
    wire \uu2.N_101 ;
    wire \uu2.N_111 ;
    wire \uu2.un28_w_addr_user_i_0 ;
    wire \uu2.w_addr_userZ0Z_7 ;
    wire o_One_Sec_Pulse;
    wire \uu2.bitmapZ0Z_111 ;
    wire \uu2.vram_rd_clkZ0 ;
    wire \uu2.vram_rd_clk_detZ0Z_0 ;
    wire \uu2.vram_rd_clk_detZ0Z_1 ;
    wire \uu2.bitmapZ0Z_180 ;
    wire \uu2.bitmapZ0Z_215 ;
    wire \Lab_UT.sec1_2 ;
    wire \Lab_UT.sec1_1 ;
    wire \Lab_UT.sec1_0 ;
    wire \uu2.bitmapZ0Z_212 ;
    wire \INVuu2.w_addr_user_7C_net ;
    wire \Lab_UT.sec1_3 ;
    wire \Lab_UT.di_AMtens_1 ;
    wire \Lab_UT.di_AMtens_2 ;
    wire \Lab_UT.didp.countrce4.q_5_1_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_1 ;
    wire \Lab_UT.didp.countrce4.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_5_2_cascade_ ;
    wire \Lab_UT.dictrl.N_95_cascade_ ;
    wire \Lab_UT.dictrl.N_21_0_cascade_ ;
    wire \Lab_UT.i16_mux ;
    wire \Lab_UT.dictrl.i18_mux ;
    wire \Lab_UT.dispString.dOut_RNO_1Z0Z_1 ;
    wire \Lab_UT.dispString.cntZ0Z_0 ;
    wire \Lab_UT.dispString.cntZ0Z_1 ;
    wire \Lab_UT.dispString.m49_ns_1 ;
    wire \Lab_UT.didp.countrce1.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce1.q_5_3_cascade_ ;
    wire \Lab_UT.un1_idle_1_0_iclkZ0 ;
    wire G_186_cascade_;
    wire G_191;
    wire \Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_ ;
    wire \Lab_UT.dictrl.G_10_1 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ;
    wire \Lab_UT.dicRun_2 ;
    wire \Lab_UT.didp.ceZ0Z_0 ;
    wire \Lab_UT.didp.ceZ0Z_1 ;
    wire \buart.Z_rx.hhZ0Z_1 ;
    wire \Lab_UT.dictrl.N_90_0 ;
    wire \Lab_UT.dictrl.N_95_0 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ;
    wire \Lab_UT.LdStens_i_3 ;
    wire \Lab_UT.dictrl.state_fast_1 ;
    wire \Lab_UT.dictrl.N_95_0_0_cascade_ ;
    wire \Lab_UT.dictrl.g0_3_0_cascade_ ;
    wire \Lab_UT.dictrl.g4_cascade_ ;
    wire \Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_ ;
    wire \Lab_UT.dictrl.g2_5 ;
    wire \Lab_UT.dictrl.g0_2Z0Z_5_cascade_ ;
    wire \Lab_UT.dictrl.g2_0 ;
    wire \Lab_UT.dictrl.g1_1 ;
    wire \Lab_UT.dictrl.g2_0_cascade_ ;
    wire \Lab_UT.dictrl.N_90_0_0_0 ;
    wire \Lab_UT.dictrl.m40_N_5_mux_0 ;
    wire \Lab_UT.dictrl.g2Z0Z_1_cascade_ ;
    wire \Lab_UT.dictrl.g1_0 ;
    wire \Lab_UT.dictrl.g0_17_a6_2_1 ;
    wire \Lab_UT.dictrl.g0_17_a6_3_6 ;
    wire \Lab_UT.dictrl.g0_17_a6_3_8 ;
    wire \Lab_UT.dictrl.N_22_cascade_ ;
    wire \Lab_UT.dictrl.g0_17_0_cascade_ ;
    wire \Lab_UT.dictrl.g2_0_0 ;
    wire bu_rx_data_fast_3;
    wire \Lab_UT.didp.reset_12_1_3 ;
    wire \Lab_UT.didp.di_Mtens_2 ;
    wire \Lab_UT.didp.ce_12_3_cascade_ ;
    wire oneSecStrb;
    wire \Lab_UT.didp.countrce2.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.countrce4.q_5_0 ;
    wire \Lab_UT.didp.ceZ0Z_3 ;
    wire \Lab_UT.didp.un24_ce_2 ;
    wire \Lab_UT.LdMtens ;
    wire \Lab_UT.didp.countrce4.un20_qPone ;
    wire \Lab_UT.didp.resetZ0Z_3 ;
    wire \Lab_UT.didp.countrce4.q_5_3_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdMtens_0 ;
    wire \Lab_UT.didp.countrce2.q_5_1 ;
    wire \Lab_UT.didp.countrce3.un20_qPone_cascade_ ;
    wire \Lab_UT.didp.di_Mtens_3 ;
    wire \Lab_UT.didp.countrce2.q_5_3 ;
    wire \Lab_UT.didp.countrce2.q_5_0 ;
    wire \Lab_UT.didp.di_Stens_0 ;
    wire \Lab_UT.didp.di_Stens_1 ;
    wire \Lab_UT.didp.di_Stens_3 ;
    wire \Lab_UT.didp.regrce3.did_alarmMatch_3 ;
    wire \Lab_UT.didp.did_alarmMatch_0 ;
    wire \Lab_UT.didp.did_alarmMatch_1_cascade_ ;
    wire \Lab_UT.didp.did_alarmMatch_2 ;
    wire \Lab_UT.didp.un1_dicLdStens_0 ;
    wire \Lab_UT.didp.resetZ0Z_1 ;
    wire \Lab_UT.didp.did_alarmMatch_7 ;
    wire \Lab_UT.didp.did_alarmMatch_4_cascade_ ;
    wire \Lab_UT.didp.did_alarmMatch_5 ;
    wire \Lab_UT.did_alarmMatch_13_cascade_ ;
    wire \Lab_UT.dictrl.alarmstate_1_0_cascade_ ;
    wire \Lab_UT.did_alarmMatch_13 ;
    wire G_183_cascade_;
    wire \Lab_UT.did_alarmMatch_12 ;
    wire \Lab_UT.didp.countrce2.un13_qPone ;
    wire \Lab_UT.didp.di_Stens_2 ;
    wire \Lab_UT.didp.countrce2.q_5_2 ;
    wire rst;
    wire \Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ;
    wire G_184;
    wire \Lab_UT.alarmstate_0_sqmuxa_1 ;
    wire \Lab_UT.didp.countrce1.un13_qPone ;
    wire \Lab_UT.didp.countrce1.q_5_2_cascade_ ;
    wire \Lab_UT.didp.un1_dicLdSones_0 ;
    wire \Lab_UT.didp.resetZ0Z_0 ;
    wire \Lab_UT.un1_armed_2_0_iso_iZ0 ;
    wire \Lab_UT.un1_idle_5_0_iclkZ0 ;
    wire CONSTANT_ONE_NET;
    wire \Lab_UT.un1_armed_2_0_iso_iZ0_cascade_ ;
    wire G_192;
    wire \Lab_UT.dictrl.N_113_cascade_ ;
    wire \Lab_UT.dictrl.state_fast_2 ;
    wire \Lab_UT.dictrl.g0_17_0 ;
    wire \Lab_UT.dictrl.g0_17_1 ;
    wire \Lab_UT.didp.di_Sones_2 ;
    wire \Lab_UT.didp.di_Sones_3 ;
    wire \Lab_UT.didp.un18_ce ;
    wire \Lab_UT.LdSones_i_3 ;
    wire \Lab_UT.dictrl.next_stateZ0Z_1 ;
    wire \Lab_UT.LdStens ;
    wire bu_rx_data_rdy_0_g;
    wire \Lab_UT.dictrl.m30_0Z0Z_0 ;
    wire \Lab_UT.dictrl.m25Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.m59_ns_1_xZ0Z1 ;
    wire \Lab_UT.dictrl.N_81_1_cascade_ ;
    wire \Lab_UT.dictrl.N_113_1 ;
    wire \Lab_UT.dictrl.N_113_1_cascade_ ;
    wire \Lab_UT.dictrl.next_stateZ0Z_0 ;
    wire \Lab_UT.dictrl.m59_ns_1 ;
    wire \Lab_UT.dictrl.N_81_0 ;
    wire \Lab_UT.dictrl.N_16_mux_0_cascade_ ;
    wire \Lab_UT.dictrl.N_113_0_0 ;
    wire \Lab_UT.dictrl.state_2_rep1 ;
    wire \Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_ ;
    wire \Lab_UT.dictrl.N_5_0 ;
    wire \Lab_UT.dictrl.g2_2_cascade_ ;
    wire \Lab_UT.dictrl.i9_mux_0 ;
    wire \Lab_UT.dictrl.N_77_0 ;
    wire \Lab_UT.dictrl.state_3_rep1 ;
    wire \Lab_UT.dictrl.g0_0Z0Z_1 ;
    wire \Lab_UT.dictrl.g0_2Z0Z_4 ;
    wire \Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.N_77_1_0 ;
    wire \Lab_UT.dictrl.N_77_1_0_cascade_ ;
    wire \Lab_UT.dictrl.N_2353_0_0 ;
    wire buart__rx_shifter_fast_6;
    wire bu_rx_data_fast_7;
    wire \Lab_UT.dictrl.state_fast_3 ;
    wire \Lab_UT.dictrl.g1_6 ;
    wire \Lab_UT.dictrl.m47_xZ0Z0_cascade_ ;
    wire bu_rx_data_fast_4;
    wire \Lab_UT.dictrl.m30Z0Z_1 ;
    wire bu_rx_data_fast_1;
    wire bu_rx_data_3_rep1;
    wire \Lab_UT.dictrl.g1_1Z0Z_1 ;
    wire \Lab_UT.dictrl.g2_1_0 ;
    wire \Lab_UT.dictrl.g2 ;
    wire \Lab_UT.didp.countrce3.ce_12_2_3 ;
    wire \Lab_UT.di_AMtens_3 ;
    wire \Lab_UT.didp.regrce4.LdAMtens_0 ;
    wire \Lab_UT.didp.un1_dicLdMones_0_cascade_ ;
    wire \Lab_UT.didp.countrce3.q_5_1 ;
    wire \Lab_UT.didp.ceZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_0 ;
    wire \Lab_UT.didp.di_Mtens_0 ;
    wire \Lab_UT.di_AMtens_0 ;
    wire \Lab_UT.didp.regrce4.did_alarmMatch_6 ;
    wire \Lab_UT.didp.resetZ0Z_2 ;
    wire \Lab_UT.didp.countrce3.q_5_3 ;
    wire \Lab_UT.didp.un1_dicLdMones_0 ;
    wire \Lab_UT.didp.di_Mones_3 ;
    wire \Lab_UT.didp.di_Mones_0 ;
    wire \Lab_UT.didp.di_Mones_1 ;
    wire \Lab_UT.LdMones ;
    wire \Lab_UT.didp.countrce3.un13_qPone_cascade_ ;
    wire \Lab_UT.didp.di_Mones_2 ;
    wire \Lab_UT.didp.countrce3.q_5_2 ;
    wire \Lab_UT.di_AStens_0 ;
    wire \Lab_UT.di_AStens_1 ;
    wire \Lab_UT.di_AStens_2 ;
    wire \Lab_UT.di_AStens_3 ;
    wire \Lab_UT.di_AMones_0 ;
    wire \Lab_UT.di_AMones_1 ;
    wire \Lab_UT.di_AMones_2 ;
    wire \Lab_UT.N_13_0 ;
    wire \Lab_UT.di_AMones_3 ;
    wire \Lab_UT.di_ASones_1 ;
    wire \Lab_UT.di_ASones_2 ;
    wire \Lab_UT.di_ASones_3 ;
    wire G_183;
    wire G_185;
    wire \Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.m3_0 ;
    wire \Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_ ;
    wire G_188;
    wire \Lab_UT.dictrl.alarmstate8Z0Z_3 ;
    wire G_188_cascade_;
    wire G_187;
    wire G_186;
    wire G_187_cascade_;
    wire \Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ;
    wire \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ;
    wire \Lab_UT.state_i_3_0 ;
    wire \Lab_UT.dictrl.g0_2Z0Z_2_cascade_ ;
    wire \Lab_UT.dictrl.m40_N_5_mux_1 ;
    wire \Lab_UT.dictrl.alarmstate8Z0Z_4 ;
    wire \Lab_UT.didp.di_Sones_0 ;
    wire \Lab_UT.LdSones ;
    wire \Lab_UT.didp.di_Sones_1 ;
    wire \Lab_UT.didp.countrce1.q_5_1 ;
    wire \Lab_UT.dictrl.N_4_cascade_ ;
    wire \Lab_UT.dictrl.N_12 ;
    wire \Lab_UT.dictrl.N_81 ;
    wire \Lab_UT.dictrl.next_state_i_1_2 ;
    wire \Lab_UT.dictrl.P8_mux ;
    wire \Lab_UT.dictrl.next_state_1_3 ;
    wire \Lab_UT.dictrl.P6_mux_0 ;
    wire \Lab_UT.dictrl.state_i_3_2 ;
    wire \Lab_UT.dictrl.N_114_mux ;
    wire \Lab_UT.dictrl.N_69 ;
    wire \Lab_UT.dictrl.i10_mux ;
    wire \Lab_UT.dictrl.N_69_cascade_ ;
    wire \Lab_UT.dictrl.next_state_1_0_3 ;
    wire \Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1 ;
    wire \Lab_UT.dictrl.g0_17_a6_0_1 ;
    wire \Lab_UT.dictrl.P6_mux ;
    wire \Lab_UT.dictrl.N_189 ;
    wire \Lab_UT.dictrl.m40_N_5_mux ;
    wire \Lab_UT.dictrl.N_77 ;
    wire \Lab_UT.dictrl.N_77_cascade_ ;
    wire \Lab_UT.dictrl.m73Z0Z_1 ;
    wire \Lab_UT.dictrl.m77_ns_1 ;
    wire \Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_ ;
    wire \Lab_UT.dictrl.i9_mux_0_0 ;
    wire \Lab_UT.dictrl.N_106_mux ;
    wire \Lab_UT.dictrl.m51_0 ;
    wire \Lab_UT.dictrl.state_i_3_1 ;
    wire \Lab_UT.dictrl.N_118_mux_cascade_ ;
    wire \Lab_UT.dictrl.next_state_latmux_3_1_1 ;
    wire \Lab_UT.dictrl.g0_17_a6_3Z0Z_7 ;
    wire buart__rx_shifter_fast_0;
    wire bu_rx_data_1_rep1;
    wire bu_rx_data_fast_2;
    wire buart__rx_shifter_fast_5;
    wire bu_rx_data_2_rep1;
    wire \Lab_UT.dictrl.N_103_mux ;
    wire \Lab_UT.dictrl.N_4_0_cascade_ ;
    wire \Lab_UT.dictrl.state_1_rep1 ;
    wire \Lab_UT.dictrl.N_12_0 ;
    wire \Lab_UT.LdASones ;
    wire \Lab_UT.didp.regrce1.LdASones_0 ;
    wire bu_rx_data_7_rep1;
    wire shifter_7_rep1_RNIG7Q01;
    wire \buart.Z_rx.P7_mux ;
    wire N_16_mux;
    wire shifter_7_rep1_RNIG7Q01_cascade_;
    wire N_97;
    wire bu_rx_data_4_rep1;
    wire bu_rx_data_rdy_0;
    wire Lab_UT_dictrl_state_3_rep2;
    wire \Lab_UT.dictrl.g0_5_a4_1_5_cascade_ ;
    wire \Lab_UT.dictrl.N_13_cascade_ ;
    wire \Lab_UT.dictrl.N_90 ;
    wire \buart.Z_rx.sample_g ;
    wire rst_g;
    wire bu_rx_data_rdy;
    wire \Lab_UT.dictrl.m25Z0Z_0 ;
    wire N_119_mux_cascade_;
    wire bu_rx_data_3_rep2;
    wire \Lab_UT.dictrl.g0_5_a4_1_4 ;
    wire \Lab_UT.dictrl.m86Z0Z_0_cascade_ ;
    wire \Lab_UT.dictrl.m86Z0Z_2 ;
    wire \Lab_UT.state_3 ;
    wire \Lab_UT.dictrl.un1_next_state66_0 ;
    wire \Lab_UT.state_0 ;
    wire \Lab_UT.dictrl.next_state_latmux_1_a0_0_0 ;
    wire bu_rx_data_2;
    wire bu_rx_data_5;
    wire bu_rx_data_3;
    wire bu_rx_data_7;
    wire bu_rx_data_1;
    wire bu_rx_data_6;
    wire bu_rx_data_4;
    wire bu_rx_data_0;
    wire \Lab_UT.dictrl.g0_5_o4_3 ;
    wire \Lab_UT.dictrl.stateZ0Z_2 ;
    wire \Lab_UT.dictrl.g0_5_o4_4_cascade_ ;
    wire \Lab_UT.dictrl.stateZ0Z_1 ;
    wire \Lab_UT.dictrl.N_11 ;
    wire N_117_cascade_;
    wire resetGen_reset_count_0;
    wire resetGen_reset_count_1;
    wire resetGen_reset_count_2_2_cascade_;
    wire resetGen_reset_count_2;
    wire \resetGen.reset_countZ0Z_3 ;
    wire N_91_i;
    wire clk_g;
    wire N_119_mux;
    wire resetGen_reset_count_4;
    wire m87;
    wire _gnd_net_;

    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .TEST_MODE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .PLLOUT_SELECT="GENCLK";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FILTER_RANGE=3'b001;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .ENABLE_ICEGATE=1'b0;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVR=4'b0000;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVQ=3'b110;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DIVF=7'b0111111;
    defparam \latticehx1k_pll_inst.latticehx1k_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \latticehx1k_pll_inst.latticehx1k_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .SCLK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(clk),
            .REFERENCECLK(N__7686),
            .RESETB(N__15729),
            .BYPASS(GNDG0),
            .SDI(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_0=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .WRITE_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .READ_MODE=1;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_F=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_E=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_D=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_C=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_B=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_A=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_9=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_8=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_7=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_6=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_5=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_4=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_3=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_2=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    defparam \uu2.mem0.ram512X8_inst_physical .INIT_1=256'b0000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000;
    SB_RAM40_4K \uu2.mem0.ram512X8_inst_physical  (
            .RDATA({dangling_wire_0,\uu2.r_data_wire_7 ,dangling_wire_1,\uu2.r_data_wire_6 ,dangling_wire_2,\uu2.r_data_wire_5 ,dangling_wire_3,\uu2.r_data_wire_4 ,dangling_wire_4,\uu2.r_data_wire_3 ,dangling_wire_5,\uu2.r_data_wire_2 ,dangling_wire_6,\uu2.r_data_wire_1 ,dangling_wire_7,\uu2.r_data_wire_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__8436,N__8412,N__8385,N__8475,N__8538,N__8361,N__8328,N__8577,N__8619}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__9489,N__9528,N__9540,N__10239,N__7725,N__9777,N__7752,N__7698,N__7713}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__8103,dangling_wire_31,N__8295,dangling_wire_32,N__8280,dangling_wire_33,N__8259,dangling_wire_34,N__9981,dangling_wire_35,N__8286,dangling_wire_36,N__8229}),
            .RCLKE(),
            .RCLK(N__21667),
            .RE(N__15744),
            .WCLKE(N__9737),
            .WCLK(N__21666),
            .WE(N__9738));
    IO_PAD led_obuft_3_iopad (
            .OE(N__21862),
            .DIN(N__21861),
            .DOUT(N__21860),
            .PACKAGEPIN(led[3]));
    defparam led_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_3_preio (
            .PADOEN(N__21862),
            .PADOUT(N__21861),
            .PADIN(N__21860),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_0_iopad (
            .OE(N__21853),
            .DIN(N__21852),
            .DOUT(N__21851),
            .PACKAGEPIN(led[0]));
    defparam led_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_0_preio (
            .PADOEN(N__21853),
            .PADOUT(N__21852),
            .PADIN(N__21851),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_4_iopad (
            .OE(N__21844),
            .DIN(N__21843),
            .DOUT(N__21842),
            .PACKAGEPIN(led[4]));
    defparam led_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_4_preio (
            .PADOEN(N__21844),
            .PADOUT(N__21843),
            .PADIN(N__21842),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD \Z_rcxd.Z_io_iopad  (
            .OE(N__21835),
            .DIN(N__21834),
            .DOUT(N__21833),
            .PACKAGEPIN(from_pc));
    defparam \Z_rcxd.Z_io_preio .PIN_TYPE=6'b000000;
    PRE_IO \Z_rcxd.Z_io_preio  (
            .PADOEN(N__21835),
            .PADOUT(N__21834),
            .PADIN(N__21833),
            .CLOCKENABLE(),
            .DOUT1(GNDG0),
            .OUTPUTENABLE(),
            .DIN0(uart_RXD),
            .DOUT0(GNDG0),
            .INPUTCLK(N__21630),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clk_in_ibuf_iopad (
            .OE(N__21826),
            .DIN(N__21825),
            .DOUT(N__21824),
            .PACKAGEPIN(clk_in));
    defparam clk_in_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_in_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_in_ibuf_preio (
            .PADOEN(N__21826),
            .PADOUT(N__21825),
            .PADIN(N__21824),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_in_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_1_iopad (
            .OE(N__21817),
            .DIN(N__21816),
            .DOUT(N__21815),
            .PACKAGEPIN(led[1]));
    defparam led_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_1_preio (
            .PADOEN(N__21817),
            .PADOUT(N__21816),
            .PADIN(N__21815),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD led_obuft_2_iopad (
            .OE(N__21808),
            .DIN(N__21807),
            .DOUT(N__21806),
            .PACKAGEPIN(led[2]));
    defparam led_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam led_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO led_obuft_2_preio (
            .PADOEN(N__21808),
            .PADOUT(N__21807),
            .PADIN(N__21806),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD to_ir_obuf_iopad (
            .OE(N__21799),
            .DIN(N__21798),
            .DOUT(N__21797),
            .PACKAGEPIN(to_ir));
    defparam to_ir_obuf_preio.NEG_TRIGGER=1'b0;
    defparam to_ir_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO to_ir_obuf_preio (
            .PADOEN(N__21799),
            .PADOUT(N__21798),
            .PADIN(N__21797),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_serial_data_obuf_iopad (
            .OE(N__21790),
            .DIN(N__21789),
            .DOUT(N__21788),
            .PACKAGEPIN(o_serial_data));
    defparam o_serial_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam o_serial_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO o_serial_data_obuf_preio (
            .PADOEN(N__21790),
            .PADOUT(N__21789),
            .PADIN(N__21788),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11433),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sd_obuf_iopad (
            .OE(N__21781),
            .DIN(N__21780),
            .DOUT(N__21779),
            .PACKAGEPIN(sd));
    defparam sd_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sd_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sd_obuf_preio (
            .PADOEN(N__21781),
            .PADOUT(N__21780),
            .PADIN(N__21779),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__5345 (
            .O(N__21762),
            .I(N_117_cascade_));
    InMux I__5344 (
            .O(N__21759),
            .I(N__21752));
    InMux I__5343 (
            .O(N__21758),
            .I(N__21743));
    InMux I__5342 (
            .O(N__21757),
            .I(N__21743));
    InMux I__5341 (
            .O(N__21756),
            .I(N__21743));
    InMux I__5340 (
            .O(N__21755),
            .I(N__21743));
    LocalMux I__5339 (
            .O(N__21752),
            .I(resetGen_reset_count_0));
    LocalMux I__5338 (
            .O(N__21743),
            .I(resetGen_reset_count_0));
    CascadeMux I__5337 (
            .O(N__21738),
            .I(N__21734));
    CascadeMux I__5336 (
            .O(N__21737),
            .I(N__21731));
    InMux I__5335 (
            .O(N__21734),
            .I(N__21720));
    InMux I__5334 (
            .O(N__21731),
            .I(N__21720));
    InMux I__5333 (
            .O(N__21730),
            .I(N__21720));
    InMux I__5332 (
            .O(N__21729),
            .I(N__21720));
    LocalMux I__5331 (
            .O(N__21720),
            .I(resetGen_reset_count_1));
    CascadeMux I__5330 (
            .O(N__21717),
            .I(resetGen_reset_count_2_2_cascade_));
    CascadeMux I__5329 (
            .O(N__21714),
            .I(N__21708));
    CascadeMux I__5328 (
            .O(N__21713),
            .I(N__21705));
    InMux I__5327 (
            .O(N__21712),
            .I(N__21696));
    InMux I__5326 (
            .O(N__21711),
            .I(N__21696));
    InMux I__5325 (
            .O(N__21708),
            .I(N__21696));
    InMux I__5324 (
            .O(N__21705),
            .I(N__21696));
    LocalMux I__5323 (
            .O(N__21696),
            .I(resetGen_reset_count_2));
    CascadeMux I__5322 (
            .O(N__21693),
            .I(N__21690));
    InMux I__5321 (
            .O(N__21690),
            .I(N__21684));
    InMux I__5320 (
            .O(N__21689),
            .I(N__21684));
    LocalMux I__5319 (
            .O(N__21684),
            .I(\resetGen.reset_countZ0Z_3 ));
    InMux I__5318 (
            .O(N__21681),
            .I(N__21675));
    InMux I__5317 (
            .O(N__21680),
            .I(N__21675));
    LocalMux I__5316 (
            .O(N__21675),
            .I(N_91_i));
    ClkMux I__5315 (
            .O(N__21672),
            .I(N__21429));
    ClkMux I__5314 (
            .O(N__21671),
            .I(N__21429));
    ClkMux I__5313 (
            .O(N__21670),
            .I(N__21429));
    ClkMux I__5312 (
            .O(N__21669),
            .I(N__21429));
    ClkMux I__5311 (
            .O(N__21668),
            .I(N__21429));
    ClkMux I__5310 (
            .O(N__21667),
            .I(N__21429));
    ClkMux I__5309 (
            .O(N__21666),
            .I(N__21429));
    ClkMux I__5308 (
            .O(N__21665),
            .I(N__21429));
    ClkMux I__5307 (
            .O(N__21664),
            .I(N__21429));
    ClkMux I__5306 (
            .O(N__21663),
            .I(N__21429));
    ClkMux I__5305 (
            .O(N__21662),
            .I(N__21429));
    ClkMux I__5304 (
            .O(N__21661),
            .I(N__21429));
    ClkMux I__5303 (
            .O(N__21660),
            .I(N__21429));
    ClkMux I__5302 (
            .O(N__21659),
            .I(N__21429));
    ClkMux I__5301 (
            .O(N__21658),
            .I(N__21429));
    ClkMux I__5300 (
            .O(N__21657),
            .I(N__21429));
    ClkMux I__5299 (
            .O(N__21656),
            .I(N__21429));
    ClkMux I__5298 (
            .O(N__21655),
            .I(N__21429));
    ClkMux I__5297 (
            .O(N__21654),
            .I(N__21429));
    ClkMux I__5296 (
            .O(N__21653),
            .I(N__21429));
    ClkMux I__5295 (
            .O(N__21652),
            .I(N__21429));
    ClkMux I__5294 (
            .O(N__21651),
            .I(N__21429));
    ClkMux I__5293 (
            .O(N__21650),
            .I(N__21429));
    ClkMux I__5292 (
            .O(N__21649),
            .I(N__21429));
    ClkMux I__5291 (
            .O(N__21648),
            .I(N__21429));
    ClkMux I__5290 (
            .O(N__21647),
            .I(N__21429));
    ClkMux I__5289 (
            .O(N__21646),
            .I(N__21429));
    ClkMux I__5288 (
            .O(N__21645),
            .I(N__21429));
    ClkMux I__5287 (
            .O(N__21644),
            .I(N__21429));
    ClkMux I__5286 (
            .O(N__21643),
            .I(N__21429));
    ClkMux I__5285 (
            .O(N__21642),
            .I(N__21429));
    ClkMux I__5284 (
            .O(N__21641),
            .I(N__21429));
    ClkMux I__5283 (
            .O(N__21640),
            .I(N__21429));
    ClkMux I__5282 (
            .O(N__21639),
            .I(N__21429));
    ClkMux I__5281 (
            .O(N__21638),
            .I(N__21429));
    ClkMux I__5280 (
            .O(N__21637),
            .I(N__21429));
    ClkMux I__5279 (
            .O(N__21636),
            .I(N__21429));
    ClkMux I__5278 (
            .O(N__21635),
            .I(N__21429));
    ClkMux I__5277 (
            .O(N__21634),
            .I(N__21429));
    ClkMux I__5276 (
            .O(N__21633),
            .I(N__21429));
    ClkMux I__5275 (
            .O(N__21632),
            .I(N__21429));
    ClkMux I__5274 (
            .O(N__21631),
            .I(N__21429));
    ClkMux I__5273 (
            .O(N__21630),
            .I(N__21429));
    ClkMux I__5272 (
            .O(N__21629),
            .I(N__21429));
    ClkMux I__5271 (
            .O(N__21628),
            .I(N__21429));
    ClkMux I__5270 (
            .O(N__21627),
            .I(N__21429));
    ClkMux I__5269 (
            .O(N__21626),
            .I(N__21429));
    ClkMux I__5268 (
            .O(N__21625),
            .I(N__21429));
    ClkMux I__5267 (
            .O(N__21624),
            .I(N__21429));
    ClkMux I__5266 (
            .O(N__21623),
            .I(N__21429));
    ClkMux I__5265 (
            .O(N__21622),
            .I(N__21429));
    ClkMux I__5264 (
            .O(N__21621),
            .I(N__21429));
    ClkMux I__5263 (
            .O(N__21620),
            .I(N__21429));
    ClkMux I__5262 (
            .O(N__21619),
            .I(N__21429));
    ClkMux I__5261 (
            .O(N__21618),
            .I(N__21429));
    ClkMux I__5260 (
            .O(N__21617),
            .I(N__21429));
    ClkMux I__5259 (
            .O(N__21616),
            .I(N__21429));
    ClkMux I__5258 (
            .O(N__21615),
            .I(N__21429));
    ClkMux I__5257 (
            .O(N__21614),
            .I(N__21429));
    ClkMux I__5256 (
            .O(N__21613),
            .I(N__21429));
    ClkMux I__5255 (
            .O(N__21612),
            .I(N__21429));
    ClkMux I__5254 (
            .O(N__21611),
            .I(N__21429));
    ClkMux I__5253 (
            .O(N__21610),
            .I(N__21429));
    ClkMux I__5252 (
            .O(N__21609),
            .I(N__21429));
    ClkMux I__5251 (
            .O(N__21608),
            .I(N__21429));
    ClkMux I__5250 (
            .O(N__21607),
            .I(N__21429));
    ClkMux I__5249 (
            .O(N__21606),
            .I(N__21429));
    ClkMux I__5248 (
            .O(N__21605),
            .I(N__21429));
    ClkMux I__5247 (
            .O(N__21604),
            .I(N__21429));
    ClkMux I__5246 (
            .O(N__21603),
            .I(N__21429));
    ClkMux I__5245 (
            .O(N__21602),
            .I(N__21429));
    ClkMux I__5244 (
            .O(N__21601),
            .I(N__21429));
    ClkMux I__5243 (
            .O(N__21600),
            .I(N__21429));
    ClkMux I__5242 (
            .O(N__21599),
            .I(N__21429));
    ClkMux I__5241 (
            .O(N__21598),
            .I(N__21429));
    ClkMux I__5240 (
            .O(N__21597),
            .I(N__21429));
    ClkMux I__5239 (
            .O(N__21596),
            .I(N__21429));
    ClkMux I__5238 (
            .O(N__21595),
            .I(N__21429));
    ClkMux I__5237 (
            .O(N__21594),
            .I(N__21429));
    ClkMux I__5236 (
            .O(N__21593),
            .I(N__21429));
    ClkMux I__5235 (
            .O(N__21592),
            .I(N__21429));
    GlobalMux I__5234 (
            .O(N__21429),
            .I(N__21426));
    gio2CtrlBuf I__5233 (
            .O(N__21426),
            .I(clk_g));
    InMux I__5232 (
            .O(N__21423),
            .I(N__21402));
    InMux I__5231 (
            .O(N__21422),
            .I(N__21402));
    InMux I__5230 (
            .O(N__21421),
            .I(N__21402));
    InMux I__5229 (
            .O(N__21420),
            .I(N__21402));
    InMux I__5228 (
            .O(N__21419),
            .I(N__21402));
    InMux I__5227 (
            .O(N__21418),
            .I(N__21402));
    InMux I__5226 (
            .O(N__21417),
            .I(N__21402));
    LocalMux I__5225 (
            .O(N__21402),
            .I(N_119_mux));
    InMux I__5224 (
            .O(N__21399),
            .I(N__21393));
    InMux I__5223 (
            .O(N__21398),
            .I(N__21388));
    InMux I__5222 (
            .O(N__21397),
            .I(N__21383));
    InMux I__5221 (
            .O(N__21396),
            .I(N__21383));
    LocalMux I__5220 (
            .O(N__21393),
            .I(N__21380));
    InMux I__5219 (
            .O(N__21392),
            .I(N__21375));
    InMux I__5218 (
            .O(N__21391),
            .I(N__21375));
    LocalMux I__5217 (
            .O(N__21388),
            .I(resetGen_reset_count_4));
    LocalMux I__5216 (
            .O(N__21383),
            .I(resetGen_reset_count_4));
    Odrv12 I__5215 (
            .O(N__21380),
            .I(resetGen_reset_count_4));
    LocalMux I__5214 (
            .O(N__21375),
            .I(resetGen_reset_count_4));
    InMux I__5213 (
            .O(N__21366),
            .I(N__21363));
    LocalMux I__5212 (
            .O(N__21363),
            .I(m87));
    CascadeMux I__5211 (
            .O(N__21360),
            .I(N_119_mux_cascade_));
    CascadeMux I__5210 (
            .O(N__21357),
            .I(N__21352));
    CascadeMux I__5209 (
            .O(N__21356),
            .I(N__21349));
    CascadeMux I__5208 (
            .O(N__21355),
            .I(N__21345));
    InMux I__5207 (
            .O(N__21352),
            .I(N__21342));
    InMux I__5206 (
            .O(N__21349),
            .I(N__21339));
    InMux I__5205 (
            .O(N__21348),
            .I(N__21334));
    InMux I__5204 (
            .O(N__21345),
            .I(N__21334));
    LocalMux I__5203 (
            .O(N__21342),
            .I(N__21329));
    LocalMux I__5202 (
            .O(N__21339),
            .I(N__21321));
    LocalMux I__5201 (
            .O(N__21334),
            .I(N__21318));
    InMux I__5200 (
            .O(N__21333),
            .I(N__21313));
    InMux I__5199 (
            .O(N__21332),
            .I(N__21313));
    Span4Mux_s2_h I__5198 (
            .O(N__21329),
            .I(N__21310));
    InMux I__5197 (
            .O(N__21328),
            .I(N__21305));
    InMux I__5196 (
            .O(N__21327),
            .I(N__21305));
    InMux I__5195 (
            .O(N__21326),
            .I(N__21302));
    InMux I__5194 (
            .O(N__21325),
            .I(N__21297));
    InMux I__5193 (
            .O(N__21324),
            .I(N__21297));
    Span4Mux_h I__5192 (
            .O(N__21321),
            .I(N__21292));
    Span4Mux_h I__5191 (
            .O(N__21318),
            .I(N__21292));
    LocalMux I__5190 (
            .O(N__21313),
            .I(N__21289));
    Odrv4 I__5189 (
            .O(N__21310),
            .I(bu_rx_data_3_rep2));
    LocalMux I__5188 (
            .O(N__21305),
            .I(bu_rx_data_3_rep2));
    LocalMux I__5187 (
            .O(N__21302),
            .I(bu_rx_data_3_rep2));
    LocalMux I__5186 (
            .O(N__21297),
            .I(bu_rx_data_3_rep2));
    Odrv4 I__5185 (
            .O(N__21292),
            .I(bu_rx_data_3_rep2));
    Odrv12 I__5184 (
            .O(N__21289),
            .I(bu_rx_data_3_rep2));
    InMux I__5183 (
            .O(N__21276),
            .I(N__21273));
    LocalMux I__5182 (
            .O(N__21273),
            .I(\Lab_UT.dictrl.g0_5_a4_1_4 ));
    CascadeMux I__5181 (
            .O(N__21270),
            .I(\Lab_UT.dictrl.m86Z0Z_0_cascade_ ));
    InMux I__5180 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__5179 (
            .O(N__21264),
            .I(\Lab_UT.dictrl.m86Z0Z_2 ));
    CascadeMux I__5178 (
            .O(N__21261),
            .I(N__21256));
    InMux I__5177 (
            .O(N__21260),
            .I(N__21252));
    CascadeMux I__5176 (
            .O(N__21259),
            .I(N__21247));
    InMux I__5175 (
            .O(N__21256),
            .I(N__21244));
    CascadeMux I__5174 (
            .O(N__21255),
            .I(N__21240));
    LocalMux I__5173 (
            .O(N__21252),
            .I(N__21233));
    InMux I__5172 (
            .O(N__21251),
            .I(N__21230));
    InMux I__5171 (
            .O(N__21250),
            .I(N__21227));
    InMux I__5170 (
            .O(N__21247),
            .I(N__21224));
    LocalMux I__5169 (
            .O(N__21244),
            .I(N__21221));
    InMux I__5168 (
            .O(N__21243),
            .I(N__21218));
    InMux I__5167 (
            .O(N__21240),
            .I(N__21213));
    CascadeMux I__5166 (
            .O(N__21239),
            .I(N__21208));
    CascadeMux I__5165 (
            .O(N__21238),
            .I(N__21205));
    CascadeMux I__5164 (
            .O(N__21237),
            .I(N__21201));
    InMux I__5163 (
            .O(N__21236),
            .I(N__21198));
    Span4Mux_v I__5162 (
            .O(N__21233),
            .I(N__21191));
    LocalMux I__5161 (
            .O(N__21230),
            .I(N__21191));
    LocalMux I__5160 (
            .O(N__21227),
            .I(N__21188));
    LocalMux I__5159 (
            .O(N__21224),
            .I(N__21185));
    Span4Mux_h I__5158 (
            .O(N__21221),
            .I(N__21180));
    LocalMux I__5157 (
            .O(N__21218),
            .I(N__21180));
    InMux I__5156 (
            .O(N__21217),
            .I(N__21177));
    CascadeMux I__5155 (
            .O(N__21216),
            .I(N__21173));
    LocalMux I__5154 (
            .O(N__21213),
            .I(N__21170));
    InMux I__5153 (
            .O(N__21212),
            .I(N__21165));
    InMux I__5152 (
            .O(N__21211),
            .I(N__21165));
    InMux I__5151 (
            .O(N__21208),
            .I(N__21160));
    InMux I__5150 (
            .O(N__21205),
            .I(N__21160));
    InMux I__5149 (
            .O(N__21204),
            .I(N__21155));
    InMux I__5148 (
            .O(N__21201),
            .I(N__21155));
    LocalMux I__5147 (
            .O(N__21198),
            .I(N__21152));
    InMux I__5146 (
            .O(N__21197),
            .I(N__21149));
    InMux I__5145 (
            .O(N__21196),
            .I(N__21146));
    Span4Mux_h I__5144 (
            .O(N__21191),
            .I(N__21141));
    Span4Mux_h I__5143 (
            .O(N__21188),
            .I(N__21141));
    Span4Mux_h I__5142 (
            .O(N__21185),
            .I(N__21134));
    Span4Mux_h I__5141 (
            .O(N__21180),
            .I(N__21134));
    LocalMux I__5140 (
            .O(N__21177),
            .I(N__21134));
    InMux I__5139 (
            .O(N__21176),
            .I(N__21129));
    InMux I__5138 (
            .O(N__21173),
            .I(N__21129));
    Span4Mux_h I__5137 (
            .O(N__21170),
            .I(N__21122));
    LocalMux I__5136 (
            .O(N__21165),
            .I(N__21122));
    LocalMux I__5135 (
            .O(N__21160),
            .I(N__21122));
    LocalMux I__5134 (
            .O(N__21155),
            .I(\Lab_UT.state_3 ));
    Odrv12 I__5133 (
            .O(N__21152),
            .I(\Lab_UT.state_3 ));
    LocalMux I__5132 (
            .O(N__21149),
            .I(\Lab_UT.state_3 ));
    LocalMux I__5131 (
            .O(N__21146),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5130 (
            .O(N__21141),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5129 (
            .O(N__21134),
            .I(\Lab_UT.state_3 ));
    LocalMux I__5128 (
            .O(N__21129),
            .I(\Lab_UT.state_3 ));
    Odrv4 I__5127 (
            .O(N__21122),
            .I(\Lab_UT.state_3 ));
    InMux I__5126 (
            .O(N__21105),
            .I(N__21093));
    CascadeMux I__5125 (
            .O(N__21104),
            .I(N__21088));
    InMux I__5124 (
            .O(N__21103),
            .I(N__21085));
    CascadeMux I__5123 (
            .O(N__21102),
            .I(N__21080));
    InMux I__5122 (
            .O(N__21101),
            .I(N__21075));
    InMux I__5121 (
            .O(N__21100),
            .I(N__21072));
    InMux I__5120 (
            .O(N__21099),
            .I(N__21065));
    InMux I__5119 (
            .O(N__21098),
            .I(N__21065));
    InMux I__5118 (
            .O(N__21097),
            .I(N__21065));
    InMux I__5117 (
            .O(N__21096),
            .I(N__21062));
    LocalMux I__5116 (
            .O(N__21093),
            .I(N__21059));
    CascadeMux I__5115 (
            .O(N__21092),
            .I(N__21053));
    CascadeMux I__5114 (
            .O(N__21091),
            .I(N__21050));
    InMux I__5113 (
            .O(N__21088),
            .I(N__21045));
    LocalMux I__5112 (
            .O(N__21085),
            .I(N__21041));
    InMux I__5111 (
            .O(N__21084),
            .I(N__21032));
    InMux I__5110 (
            .O(N__21083),
            .I(N__21032));
    InMux I__5109 (
            .O(N__21080),
            .I(N__21032));
    InMux I__5108 (
            .O(N__21079),
            .I(N__21032));
    InMux I__5107 (
            .O(N__21078),
            .I(N__21029));
    LocalMux I__5106 (
            .O(N__21075),
            .I(N__21024));
    LocalMux I__5105 (
            .O(N__21072),
            .I(N__21024));
    LocalMux I__5104 (
            .O(N__21065),
            .I(N__21013));
    LocalMux I__5103 (
            .O(N__21062),
            .I(N__21013));
    Span4Mux_s1_h I__5102 (
            .O(N__21059),
            .I(N__21013));
    InMux I__5101 (
            .O(N__21058),
            .I(N__21002));
    InMux I__5100 (
            .O(N__21057),
            .I(N__21002));
    InMux I__5099 (
            .O(N__21056),
            .I(N__21002));
    InMux I__5098 (
            .O(N__21053),
            .I(N__21002));
    InMux I__5097 (
            .O(N__21050),
            .I(N__21002));
    InMux I__5096 (
            .O(N__21049),
            .I(N__20997));
    InMux I__5095 (
            .O(N__21048),
            .I(N__20997));
    LocalMux I__5094 (
            .O(N__21045),
            .I(N__20994));
    CascadeMux I__5093 (
            .O(N__21044),
            .I(N__20991));
    Span4Mux_v I__5092 (
            .O(N__21041),
            .I(N__20988));
    LocalMux I__5091 (
            .O(N__21032),
            .I(N__20981));
    LocalMux I__5090 (
            .O(N__21029),
            .I(N__20981));
    Span4Mux_v I__5089 (
            .O(N__21024),
            .I(N__20981));
    InMux I__5088 (
            .O(N__21023),
            .I(N__20978));
    InMux I__5087 (
            .O(N__21022),
            .I(N__20975));
    InMux I__5086 (
            .O(N__21021),
            .I(N__20970));
    InMux I__5085 (
            .O(N__21020),
            .I(N__20970));
    Span4Mux_h I__5084 (
            .O(N__21013),
            .I(N__20967));
    LocalMux I__5083 (
            .O(N__21002),
            .I(N__20964));
    LocalMux I__5082 (
            .O(N__20997),
            .I(N__20959));
    Span4Mux_v I__5081 (
            .O(N__20994),
            .I(N__20959));
    InMux I__5080 (
            .O(N__20991),
            .I(N__20956));
    Odrv4 I__5079 (
            .O(N__20988),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5078 (
            .O(N__20981),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__5077 (
            .O(N__20978),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__5076 (
            .O(N__20975),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__5075 (
            .O(N__20970),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5074 (
            .O(N__20967),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv12 I__5073 (
            .O(N__20964),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    Odrv4 I__5072 (
            .O(N__20959),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    LocalMux I__5071 (
            .O(N__20956),
            .I(\Lab_UT.dictrl.un1_next_state66_0 ));
    CascadeMux I__5070 (
            .O(N__20937),
            .I(N__20931));
    InMux I__5069 (
            .O(N__20936),
            .I(N__20920));
    InMux I__5068 (
            .O(N__20935),
            .I(N__20917));
    InMux I__5067 (
            .O(N__20934),
            .I(N__20914));
    InMux I__5066 (
            .O(N__20931),
            .I(N__20911));
    InMux I__5065 (
            .O(N__20930),
            .I(N__20908));
    InMux I__5064 (
            .O(N__20929),
            .I(N__20903));
    InMux I__5063 (
            .O(N__20928),
            .I(N__20894));
    InMux I__5062 (
            .O(N__20927),
            .I(N__20894));
    InMux I__5061 (
            .O(N__20926),
            .I(N__20894));
    InMux I__5060 (
            .O(N__20925),
            .I(N__20894));
    InMux I__5059 (
            .O(N__20924),
            .I(N__20888));
    InMux I__5058 (
            .O(N__20923),
            .I(N__20888));
    LocalMux I__5057 (
            .O(N__20920),
            .I(N__20874));
    LocalMux I__5056 (
            .O(N__20917),
            .I(N__20871));
    LocalMux I__5055 (
            .O(N__20914),
            .I(N__20866));
    LocalMux I__5054 (
            .O(N__20911),
            .I(N__20866));
    LocalMux I__5053 (
            .O(N__20908),
            .I(N__20863));
    InMux I__5052 (
            .O(N__20907),
            .I(N__20858));
    InMux I__5051 (
            .O(N__20906),
            .I(N__20858));
    LocalMux I__5050 (
            .O(N__20903),
            .I(N__20855));
    LocalMux I__5049 (
            .O(N__20894),
            .I(N__20852));
    InMux I__5048 (
            .O(N__20893),
            .I(N__20849));
    LocalMux I__5047 (
            .O(N__20888),
            .I(N__20846));
    InMux I__5046 (
            .O(N__20887),
            .I(N__20843));
    InMux I__5045 (
            .O(N__20886),
            .I(N__20840));
    InMux I__5044 (
            .O(N__20885),
            .I(N__20831));
    InMux I__5043 (
            .O(N__20884),
            .I(N__20831));
    InMux I__5042 (
            .O(N__20883),
            .I(N__20831));
    InMux I__5041 (
            .O(N__20882),
            .I(N__20831));
    InMux I__5040 (
            .O(N__20881),
            .I(N__20828));
    InMux I__5039 (
            .O(N__20880),
            .I(N__20823));
    InMux I__5038 (
            .O(N__20879),
            .I(N__20823));
    InMux I__5037 (
            .O(N__20878),
            .I(N__20818));
    InMux I__5036 (
            .O(N__20877),
            .I(N__20818));
    Span4Mux_v I__5035 (
            .O(N__20874),
            .I(N__20815));
    Span4Mux_v I__5034 (
            .O(N__20871),
            .I(N__20810));
    Span4Mux_v I__5033 (
            .O(N__20866),
            .I(N__20810));
    Span4Mux_v I__5032 (
            .O(N__20863),
            .I(N__20803));
    LocalMux I__5031 (
            .O(N__20858),
            .I(N__20803));
    Span4Mux_h I__5030 (
            .O(N__20855),
            .I(N__20803));
    Span4Mux_s3_h I__5029 (
            .O(N__20852),
            .I(N__20796));
    LocalMux I__5028 (
            .O(N__20849),
            .I(N__20796));
    Span4Mux_h I__5027 (
            .O(N__20846),
            .I(N__20796));
    LocalMux I__5026 (
            .O(N__20843),
            .I(\Lab_UT.state_0 ));
    LocalMux I__5025 (
            .O(N__20840),
            .I(\Lab_UT.state_0 ));
    LocalMux I__5024 (
            .O(N__20831),
            .I(\Lab_UT.state_0 ));
    LocalMux I__5023 (
            .O(N__20828),
            .I(\Lab_UT.state_0 ));
    LocalMux I__5022 (
            .O(N__20823),
            .I(\Lab_UT.state_0 ));
    LocalMux I__5021 (
            .O(N__20818),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5020 (
            .O(N__20815),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5019 (
            .O(N__20810),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5018 (
            .O(N__20803),
            .I(\Lab_UT.state_0 ));
    Odrv4 I__5017 (
            .O(N__20796),
            .I(\Lab_UT.state_0 ));
    InMux I__5016 (
            .O(N__20775),
            .I(N__20772));
    LocalMux I__5015 (
            .O(N__20772),
            .I(N__20769));
    Odrv12 I__5014 (
            .O(N__20769),
            .I(\Lab_UT.dictrl.next_state_latmux_1_a0_0_0 ));
    InMux I__5013 (
            .O(N__20766),
            .I(N__20761));
    InMux I__5012 (
            .O(N__20765),
            .I(N__20758));
    CascadeMux I__5011 (
            .O(N__20764),
            .I(N__20749));
    LocalMux I__5010 (
            .O(N__20761),
            .I(N__20744));
    LocalMux I__5009 (
            .O(N__20758),
            .I(N__20744));
    InMux I__5008 (
            .O(N__20757),
            .I(N__20734));
    InMux I__5007 (
            .O(N__20756),
            .I(N__20734));
    CascadeMux I__5006 (
            .O(N__20755),
            .I(N__20728));
    InMux I__5005 (
            .O(N__20754),
            .I(N__20725));
    InMux I__5004 (
            .O(N__20753),
            .I(N__20722));
    InMux I__5003 (
            .O(N__20752),
            .I(N__20719));
    InMux I__5002 (
            .O(N__20749),
            .I(N__20716));
    Span4Mux_v I__5001 (
            .O(N__20744),
            .I(N__20713));
    InMux I__5000 (
            .O(N__20743),
            .I(N__20708));
    InMux I__4999 (
            .O(N__20742),
            .I(N__20708));
    InMux I__4998 (
            .O(N__20741),
            .I(N__20705));
    InMux I__4997 (
            .O(N__20740),
            .I(N__20702));
    InMux I__4996 (
            .O(N__20739),
            .I(N__20699));
    LocalMux I__4995 (
            .O(N__20734),
            .I(N__20694));
    InMux I__4994 (
            .O(N__20733),
            .I(N__20689));
    InMux I__4993 (
            .O(N__20732),
            .I(N__20689));
    InMux I__4992 (
            .O(N__20731),
            .I(N__20686));
    InMux I__4991 (
            .O(N__20728),
            .I(N__20683));
    LocalMux I__4990 (
            .O(N__20725),
            .I(N__20680));
    LocalMux I__4989 (
            .O(N__20722),
            .I(N__20677));
    LocalMux I__4988 (
            .O(N__20719),
            .I(N__20672));
    LocalMux I__4987 (
            .O(N__20716),
            .I(N__20672));
    Span4Mux_v I__4986 (
            .O(N__20713),
            .I(N__20667));
    LocalMux I__4985 (
            .O(N__20708),
            .I(N__20662));
    LocalMux I__4984 (
            .O(N__20705),
            .I(N__20662));
    LocalMux I__4983 (
            .O(N__20702),
            .I(N__20657));
    LocalMux I__4982 (
            .O(N__20699),
            .I(N__20657));
    InMux I__4981 (
            .O(N__20698),
            .I(N__20654));
    InMux I__4980 (
            .O(N__20697),
            .I(N__20651));
    Span4Mux_s2_h I__4979 (
            .O(N__20694),
            .I(N__20648));
    LocalMux I__4978 (
            .O(N__20689),
            .I(N__20641));
    LocalMux I__4977 (
            .O(N__20686),
            .I(N__20641));
    LocalMux I__4976 (
            .O(N__20683),
            .I(N__20641));
    Span4Mux_v I__4975 (
            .O(N__20680),
            .I(N__20634));
    Span4Mux_h I__4974 (
            .O(N__20677),
            .I(N__20634));
    Span4Mux_s3_h I__4973 (
            .O(N__20672),
            .I(N__20634));
    InMux I__4972 (
            .O(N__20671),
            .I(N__20629));
    InMux I__4971 (
            .O(N__20670),
            .I(N__20629));
    Odrv4 I__4970 (
            .O(N__20667),
            .I(bu_rx_data_2));
    Odrv12 I__4969 (
            .O(N__20662),
            .I(bu_rx_data_2));
    Odrv4 I__4968 (
            .O(N__20657),
            .I(bu_rx_data_2));
    LocalMux I__4967 (
            .O(N__20654),
            .I(bu_rx_data_2));
    LocalMux I__4966 (
            .O(N__20651),
            .I(bu_rx_data_2));
    Odrv4 I__4965 (
            .O(N__20648),
            .I(bu_rx_data_2));
    Odrv12 I__4964 (
            .O(N__20641),
            .I(bu_rx_data_2));
    Odrv4 I__4963 (
            .O(N__20634),
            .I(bu_rx_data_2));
    LocalMux I__4962 (
            .O(N__20629),
            .I(bu_rx_data_2));
    InMux I__4961 (
            .O(N__20610),
            .I(N__20605));
    CascadeMux I__4960 (
            .O(N__20609),
            .I(N__20599));
    InMux I__4959 (
            .O(N__20608),
            .I(N__20596));
    LocalMux I__4958 (
            .O(N__20605),
            .I(N__20591));
    InMux I__4957 (
            .O(N__20604),
            .I(N__20588));
    InMux I__4956 (
            .O(N__20603),
            .I(N__20585));
    InMux I__4955 (
            .O(N__20602),
            .I(N__20582));
    InMux I__4954 (
            .O(N__20599),
            .I(N__20579));
    LocalMux I__4953 (
            .O(N__20596),
            .I(N__20574));
    InMux I__4952 (
            .O(N__20595),
            .I(N__20565));
    InMux I__4951 (
            .O(N__20594),
            .I(N__20565));
    Span4Mux_v I__4950 (
            .O(N__20591),
            .I(N__20558));
    LocalMux I__4949 (
            .O(N__20588),
            .I(N__20558));
    LocalMux I__4948 (
            .O(N__20585),
            .I(N__20558));
    LocalMux I__4947 (
            .O(N__20582),
            .I(N__20553));
    LocalMux I__4946 (
            .O(N__20579),
            .I(N__20553));
    InMux I__4945 (
            .O(N__20578),
            .I(N__20548));
    InMux I__4944 (
            .O(N__20577),
            .I(N__20548));
    Span4Mux_v I__4943 (
            .O(N__20574),
            .I(N__20545));
    InMux I__4942 (
            .O(N__20573),
            .I(N__20542));
    InMux I__4941 (
            .O(N__20572),
            .I(N__20537));
    InMux I__4940 (
            .O(N__20571),
            .I(N__20537));
    InMux I__4939 (
            .O(N__20570),
            .I(N__20534));
    LocalMux I__4938 (
            .O(N__20565),
            .I(N__20531));
    Span4Mux_h I__4937 (
            .O(N__20558),
            .I(N__20528));
    Span4Mux_v I__4936 (
            .O(N__20553),
            .I(N__20525));
    LocalMux I__4935 (
            .O(N__20548),
            .I(bu_rx_data_5));
    Odrv4 I__4934 (
            .O(N__20545),
            .I(bu_rx_data_5));
    LocalMux I__4933 (
            .O(N__20542),
            .I(bu_rx_data_5));
    LocalMux I__4932 (
            .O(N__20537),
            .I(bu_rx_data_5));
    LocalMux I__4931 (
            .O(N__20534),
            .I(bu_rx_data_5));
    Odrv4 I__4930 (
            .O(N__20531),
            .I(bu_rx_data_5));
    Odrv4 I__4929 (
            .O(N__20528),
            .I(bu_rx_data_5));
    Odrv4 I__4928 (
            .O(N__20525),
            .I(bu_rx_data_5));
    InMux I__4927 (
            .O(N__20508),
            .I(N__20503));
    InMux I__4926 (
            .O(N__20507),
            .I(N__20500));
    CascadeMux I__4925 (
            .O(N__20506),
            .I(N__20493));
    LocalMux I__4924 (
            .O(N__20503),
            .I(N__20483));
    LocalMux I__4923 (
            .O(N__20500),
            .I(N__20483));
    InMux I__4922 (
            .O(N__20499),
            .I(N__20478));
    InMux I__4921 (
            .O(N__20498),
            .I(N__20478));
    InMux I__4920 (
            .O(N__20497),
            .I(N__20473));
    InMux I__4919 (
            .O(N__20496),
            .I(N__20473));
    InMux I__4918 (
            .O(N__20493),
            .I(N__20468));
    InMux I__4917 (
            .O(N__20492),
            .I(N__20465));
    InMux I__4916 (
            .O(N__20491),
            .I(N__20462));
    InMux I__4915 (
            .O(N__20490),
            .I(N__20459));
    InMux I__4914 (
            .O(N__20489),
            .I(N__20454));
    InMux I__4913 (
            .O(N__20488),
            .I(N__20454));
    Span4Mux_s2_v I__4912 (
            .O(N__20483),
            .I(N__20451));
    LocalMux I__4911 (
            .O(N__20478),
            .I(N__20448));
    LocalMux I__4910 (
            .O(N__20473),
            .I(N__20445));
    InMux I__4909 (
            .O(N__20472),
            .I(N__20440));
    InMux I__4908 (
            .O(N__20471),
            .I(N__20440));
    LocalMux I__4907 (
            .O(N__20468),
            .I(N__20437));
    LocalMux I__4906 (
            .O(N__20465),
            .I(N__20432));
    LocalMux I__4905 (
            .O(N__20462),
            .I(N__20432));
    LocalMux I__4904 (
            .O(N__20459),
            .I(N__20429));
    LocalMux I__4903 (
            .O(N__20454),
            .I(N__20423));
    Span4Mux_v I__4902 (
            .O(N__20451),
            .I(N__20418));
    Span4Mux_v I__4901 (
            .O(N__20448),
            .I(N__20418));
    Span4Mux_v I__4900 (
            .O(N__20445),
            .I(N__20411));
    LocalMux I__4899 (
            .O(N__20440),
            .I(N__20411));
    Span4Mux_s2_h I__4898 (
            .O(N__20437),
            .I(N__20411));
    Span4Mux_h I__4897 (
            .O(N__20432),
            .I(N__20406));
    Span4Mux_s2_h I__4896 (
            .O(N__20429),
            .I(N__20406));
    InMux I__4895 (
            .O(N__20428),
            .I(N__20399));
    InMux I__4894 (
            .O(N__20427),
            .I(N__20399));
    InMux I__4893 (
            .O(N__20426),
            .I(N__20399));
    Odrv4 I__4892 (
            .O(N__20423),
            .I(bu_rx_data_3));
    Odrv4 I__4891 (
            .O(N__20418),
            .I(bu_rx_data_3));
    Odrv4 I__4890 (
            .O(N__20411),
            .I(bu_rx_data_3));
    Odrv4 I__4889 (
            .O(N__20406),
            .I(bu_rx_data_3));
    LocalMux I__4888 (
            .O(N__20399),
            .I(bu_rx_data_3));
    InMux I__4887 (
            .O(N__20388),
            .I(N__20381));
    InMux I__4886 (
            .O(N__20387),
            .I(N__20381));
    InMux I__4885 (
            .O(N__20386),
            .I(N__20376));
    LocalMux I__4884 (
            .O(N__20381),
            .I(N__20370));
    InMux I__4883 (
            .O(N__20380),
            .I(N__20367));
    InMux I__4882 (
            .O(N__20379),
            .I(N__20364));
    LocalMux I__4881 (
            .O(N__20376),
            .I(N__20359));
    InMux I__4880 (
            .O(N__20375),
            .I(N__20356));
    InMux I__4879 (
            .O(N__20374),
            .I(N__20353));
    InMux I__4878 (
            .O(N__20373),
            .I(N__20350));
    Span4Mux_v I__4877 (
            .O(N__20370),
            .I(N__20347));
    LocalMux I__4876 (
            .O(N__20367),
            .I(N__20344));
    LocalMux I__4875 (
            .O(N__20364),
            .I(N__20341));
    InMux I__4874 (
            .O(N__20363),
            .I(N__20336));
    InMux I__4873 (
            .O(N__20362),
            .I(N__20336));
    Span4Mux_v I__4872 (
            .O(N__20359),
            .I(N__20331));
    LocalMux I__4871 (
            .O(N__20356),
            .I(N__20331));
    LocalMux I__4870 (
            .O(N__20353),
            .I(N__20328));
    LocalMux I__4869 (
            .O(N__20350),
            .I(N__20325));
    Span4Mux_h I__4868 (
            .O(N__20347),
            .I(N__20320));
    Span4Mux_v I__4867 (
            .O(N__20344),
            .I(N__20320));
    Span4Mux_h I__4866 (
            .O(N__20341),
            .I(N__20317));
    LocalMux I__4865 (
            .O(N__20336),
            .I(bu_rx_data_7));
    Odrv4 I__4864 (
            .O(N__20331),
            .I(bu_rx_data_7));
    Odrv4 I__4863 (
            .O(N__20328),
            .I(bu_rx_data_7));
    Odrv12 I__4862 (
            .O(N__20325),
            .I(bu_rx_data_7));
    Odrv4 I__4861 (
            .O(N__20320),
            .I(bu_rx_data_7));
    Odrv4 I__4860 (
            .O(N__20317),
            .I(bu_rx_data_7));
    InMux I__4859 (
            .O(N__20304),
            .I(N__20299));
    InMux I__4858 (
            .O(N__20303),
            .I(N__20292));
    InMux I__4857 (
            .O(N__20302),
            .I(N__20289));
    LocalMux I__4856 (
            .O(N__20299),
            .I(N__20281));
    InMux I__4855 (
            .O(N__20298),
            .I(N__20278));
    InMux I__4854 (
            .O(N__20297),
            .I(N__20273));
    InMux I__4853 (
            .O(N__20296),
            .I(N__20273));
    InMux I__4852 (
            .O(N__20295),
            .I(N__20270));
    LocalMux I__4851 (
            .O(N__20292),
            .I(N__20265));
    LocalMux I__4850 (
            .O(N__20289),
            .I(N__20265));
    InMux I__4849 (
            .O(N__20288),
            .I(N__20258));
    InMux I__4848 (
            .O(N__20287),
            .I(N__20258));
    InMux I__4847 (
            .O(N__20286),
            .I(N__20255));
    InMux I__4846 (
            .O(N__20285),
            .I(N__20251));
    InMux I__4845 (
            .O(N__20284),
            .I(N__20247));
    Span4Mux_h I__4844 (
            .O(N__20281),
            .I(N__20241));
    LocalMux I__4843 (
            .O(N__20278),
            .I(N__20241));
    LocalMux I__4842 (
            .O(N__20273),
            .I(N__20234));
    LocalMux I__4841 (
            .O(N__20270),
            .I(N__20234));
    Span4Mux_h I__4840 (
            .O(N__20265),
            .I(N__20234));
    InMux I__4839 (
            .O(N__20264),
            .I(N__20229));
    InMux I__4838 (
            .O(N__20263),
            .I(N__20229));
    LocalMux I__4837 (
            .O(N__20258),
            .I(N__20224));
    LocalMux I__4836 (
            .O(N__20255),
            .I(N__20224));
    CascadeMux I__4835 (
            .O(N__20254),
            .I(N__20220));
    LocalMux I__4834 (
            .O(N__20251),
            .I(N__20217));
    InMux I__4833 (
            .O(N__20250),
            .I(N__20214));
    LocalMux I__4832 (
            .O(N__20247),
            .I(N__20211));
    InMux I__4831 (
            .O(N__20246),
            .I(N__20208));
    Sp12to4 I__4830 (
            .O(N__20241),
            .I(N__20205));
    Span4Mux_v I__4829 (
            .O(N__20234),
            .I(N__20200));
    LocalMux I__4828 (
            .O(N__20229),
            .I(N__20200));
    Span4Mux_v I__4827 (
            .O(N__20224),
            .I(N__20197));
    InMux I__4826 (
            .O(N__20223),
            .I(N__20194));
    InMux I__4825 (
            .O(N__20220),
            .I(N__20191));
    Span4Mux_v I__4824 (
            .O(N__20217),
            .I(N__20184));
    LocalMux I__4823 (
            .O(N__20214),
            .I(N__20184));
    Span4Mux_s2_h I__4822 (
            .O(N__20211),
            .I(N__20184));
    LocalMux I__4821 (
            .O(N__20208),
            .I(bu_rx_data_1));
    Odrv12 I__4820 (
            .O(N__20205),
            .I(bu_rx_data_1));
    Odrv4 I__4819 (
            .O(N__20200),
            .I(bu_rx_data_1));
    Odrv4 I__4818 (
            .O(N__20197),
            .I(bu_rx_data_1));
    LocalMux I__4817 (
            .O(N__20194),
            .I(bu_rx_data_1));
    LocalMux I__4816 (
            .O(N__20191),
            .I(bu_rx_data_1));
    Odrv4 I__4815 (
            .O(N__20184),
            .I(bu_rx_data_1));
    InMux I__4814 (
            .O(N__20169),
            .I(N__20164));
    InMux I__4813 (
            .O(N__20168),
            .I(N__20152));
    InMux I__4812 (
            .O(N__20167),
            .I(N__20149));
    LocalMux I__4811 (
            .O(N__20164),
            .I(N__20146));
    CascadeMux I__4810 (
            .O(N__20163),
            .I(N__20143));
    InMux I__4809 (
            .O(N__20162),
            .I(N__20139));
    InMux I__4808 (
            .O(N__20161),
            .I(N__20136));
    InMux I__4807 (
            .O(N__20160),
            .I(N__20133));
    InMux I__4806 (
            .O(N__20159),
            .I(N__20130));
    InMux I__4805 (
            .O(N__20158),
            .I(N__20125));
    InMux I__4804 (
            .O(N__20157),
            .I(N__20125));
    InMux I__4803 (
            .O(N__20156),
            .I(N__20122));
    InMux I__4802 (
            .O(N__20155),
            .I(N__20119));
    LocalMux I__4801 (
            .O(N__20152),
            .I(N__20116));
    LocalMux I__4800 (
            .O(N__20149),
            .I(N__20113));
    Span4Mux_s1_h I__4799 (
            .O(N__20146),
            .I(N__20110));
    InMux I__4798 (
            .O(N__20143),
            .I(N__20107));
    InMux I__4797 (
            .O(N__20142),
            .I(N__20104));
    LocalMux I__4796 (
            .O(N__20139),
            .I(N__20101));
    LocalMux I__4795 (
            .O(N__20136),
            .I(N__20098));
    LocalMux I__4794 (
            .O(N__20133),
            .I(N__20091));
    LocalMux I__4793 (
            .O(N__20130),
            .I(N__20091));
    LocalMux I__4792 (
            .O(N__20125),
            .I(N__20091));
    LocalMux I__4791 (
            .O(N__20122),
            .I(N__20084));
    LocalMux I__4790 (
            .O(N__20119),
            .I(N__20084));
    Span4Mux_s3_h I__4789 (
            .O(N__20116),
            .I(N__20084));
    Span4Mux_v I__4788 (
            .O(N__20113),
            .I(N__20079));
    Span4Mux_h I__4787 (
            .O(N__20110),
            .I(N__20079));
    LocalMux I__4786 (
            .O(N__20107),
            .I(N__20074));
    LocalMux I__4785 (
            .O(N__20104),
            .I(N__20074));
    Span4Mux_s3_h I__4784 (
            .O(N__20101),
            .I(N__20065));
    Span4Mux_v I__4783 (
            .O(N__20098),
            .I(N__20065));
    Span4Mux_v I__4782 (
            .O(N__20091),
            .I(N__20065));
    Span4Mux_v I__4781 (
            .O(N__20084),
            .I(N__20065));
    Odrv4 I__4780 (
            .O(N__20079),
            .I(bu_rx_data_6));
    Odrv4 I__4779 (
            .O(N__20074),
            .I(bu_rx_data_6));
    Odrv4 I__4778 (
            .O(N__20065),
            .I(bu_rx_data_6));
    CascadeMux I__4777 (
            .O(N__20058),
            .I(N__20053));
    InMux I__4776 (
            .O(N__20057),
            .I(N__20049));
    InMux I__4775 (
            .O(N__20056),
            .I(N__20045));
    InMux I__4774 (
            .O(N__20053),
            .I(N__20042));
    CascadeMux I__4773 (
            .O(N__20052),
            .I(N__20039));
    LocalMux I__4772 (
            .O(N__20049),
            .I(N__20034));
    InMux I__4771 (
            .O(N__20048),
            .I(N__20031));
    LocalMux I__4770 (
            .O(N__20045),
            .I(N__20026));
    LocalMux I__4769 (
            .O(N__20042),
            .I(N__20023));
    InMux I__4768 (
            .O(N__20039),
            .I(N__20020));
    InMux I__4767 (
            .O(N__20038),
            .I(N__20017));
    InMux I__4766 (
            .O(N__20037),
            .I(N__20014));
    Span4Mux_v I__4765 (
            .O(N__20034),
            .I(N__20007));
    LocalMux I__4764 (
            .O(N__20031),
            .I(N__20007));
    InMux I__4763 (
            .O(N__20030),
            .I(N__20004));
    InMux I__4762 (
            .O(N__20029),
            .I(N__20000));
    Span4Mux_v I__4761 (
            .O(N__20026),
            .I(N__19993));
    Span4Mux_s1_h I__4760 (
            .O(N__20023),
            .I(N__19993));
    LocalMux I__4759 (
            .O(N__20020),
            .I(N__19993));
    LocalMux I__4758 (
            .O(N__20017),
            .I(N__19988));
    LocalMux I__4757 (
            .O(N__20014),
            .I(N__19988));
    InMux I__4756 (
            .O(N__20013),
            .I(N__19983));
    InMux I__4755 (
            .O(N__20012),
            .I(N__19983));
    Span4Mux_v I__4754 (
            .O(N__20007),
            .I(N__19978));
    LocalMux I__4753 (
            .O(N__20004),
            .I(N__19978));
    InMux I__4752 (
            .O(N__20003),
            .I(N__19975));
    LocalMux I__4751 (
            .O(N__20000),
            .I(N__19970));
    Span4Mux_h I__4750 (
            .O(N__19993),
            .I(N__19970));
    Span4Mux_h I__4749 (
            .O(N__19988),
            .I(N__19967));
    LocalMux I__4748 (
            .O(N__19983),
            .I(bu_rx_data_4));
    Odrv4 I__4747 (
            .O(N__19978),
            .I(bu_rx_data_4));
    LocalMux I__4746 (
            .O(N__19975),
            .I(bu_rx_data_4));
    Odrv4 I__4745 (
            .O(N__19970),
            .I(bu_rx_data_4));
    Odrv4 I__4744 (
            .O(N__19967),
            .I(bu_rx_data_4));
    InMux I__4743 (
            .O(N__19956),
            .I(N__19952));
    InMux I__4742 (
            .O(N__19955),
            .I(N__19945));
    LocalMux I__4741 (
            .O(N__19952),
            .I(N__19942));
    InMux I__4740 (
            .O(N__19951),
            .I(N__19937));
    InMux I__4739 (
            .O(N__19950),
            .I(N__19937));
    InMux I__4738 (
            .O(N__19949),
            .I(N__19934));
    InMux I__4737 (
            .O(N__19948),
            .I(N__19930));
    LocalMux I__4736 (
            .O(N__19945),
            .I(N__19919));
    Span4Mux_v I__4735 (
            .O(N__19942),
            .I(N__19919));
    LocalMux I__4734 (
            .O(N__19937),
            .I(N__19919));
    LocalMux I__4733 (
            .O(N__19934),
            .I(N__19916));
    InMux I__4732 (
            .O(N__19933),
            .I(N__19913));
    LocalMux I__4731 (
            .O(N__19930),
            .I(N__19909));
    InMux I__4730 (
            .O(N__19929),
            .I(N__19906));
    InMux I__4729 (
            .O(N__19928),
            .I(N__19902));
    InMux I__4728 (
            .O(N__19927),
            .I(N__19897));
    InMux I__4727 (
            .O(N__19926),
            .I(N__19897));
    Span4Mux_h I__4726 (
            .O(N__19919),
            .I(N__19892));
    Span4Mux_h I__4725 (
            .O(N__19916),
            .I(N__19892));
    LocalMux I__4724 (
            .O(N__19913),
            .I(N__19889));
    InMux I__4723 (
            .O(N__19912),
            .I(N__19885));
    Span4Mux_s2_v I__4722 (
            .O(N__19909),
            .I(N__19880));
    LocalMux I__4721 (
            .O(N__19906),
            .I(N__19880));
    InMux I__4720 (
            .O(N__19905),
            .I(N__19877));
    LocalMux I__4719 (
            .O(N__19902),
            .I(N__19874));
    LocalMux I__4718 (
            .O(N__19897),
            .I(N__19869));
    Span4Mux_v I__4717 (
            .O(N__19892),
            .I(N__19864));
    Span4Mux_v I__4716 (
            .O(N__19889),
            .I(N__19864));
    InMux I__4715 (
            .O(N__19888),
            .I(N__19861));
    LocalMux I__4714 (
            .O(N__19885),
            .I(N__19858));
    Span4Mux_v I__4713 (
            .O(N__19880),
            .I(N__19853));
    LocalMux I__4712 (
            .O(N__19877),
            .I(N__19853));
    Span12Mux_s8_v I__4711 (
            .O(N__19874),
            .I(N__19850));
    InMux I__4710 (
            .O(N__19873),
            .I(N__19847));
    InMux I__4709 (
            .O(N__19872),
            .I(N__19844));
    Span4Mux_v I__4708 (
            .O(N__19869),
            .I(N__19839));
    Span4Mux_h I__4707 (
            .O(N__19864),
            .I(N__19839));
    LocalMux I__4706 (
            .O(N__19861),
            .I(N__19832));
    Span4Mux_h I__4705 (
            .O(N__19858),
            .I(N__19832));
    Span4Mux_h I__4704 (
            .O(N__19853),
            .I(N__19832));
    Odrv12 I__4703 (
            .O(N__19850),
            .I(bu_rx_data_0));
    LocalMux I__4702 (
            .O(N__19847),
            .I(bu_rx_data_0));
    LocalMux I__4701 (
            .O(N__19844),
            .I(bu_rx_data_0));
    Odrv4 I__4700 (
            .O(N__19839),
            .I(bu_rx_data_0));
    Odrv4 I__4699 (
            .O(N__19832),
            .I(bu_rx_data_0));
    InMux I__4698 (
            .O(N__19821),
            .I(N__19818));
    LocalMux I__4697 (
            .O(N__19818),
            .I(N__19815));
    Odrv4 I__4696 (
            .O(N__19815),
            .I(\Lab_UT.dictrl.g0_5_o4_3 ));
    InMux I__4695 (
            .O(N__19812),
            .I(N__19806));
    InMux I__4694 (
            .O(N__19811),
            .I(N__19803));
    CascadeMux I__4693 (
            .O(N__19810),
            .I(N__19799));
    CascadeMux I__4692 (
            .O(N__19809),
            .I(N__19796));
    LocalMux I__4691 (
            .O(N__19806),
            .I(N__19788));
    LocalMux I__4690 (
            .O(N__19803),
            .I(N__19788));
    InMux I__4689 (
            .O(N__19802),
            .I(N__19785));
    InMux I__4688 (
            .O(N__19799),
            .I(N__19782));
    InMux I__4687 (
            .O(N__19796),
            .I(N__19775));
    InMux I__4686 (
            .O(N__19795),
            .I(N__19771));
    InMux I__4685 (
            .O(N__19794),
            .I(N__19766));
    InMux I__4684 (
            .O(N__19793),
            .I(N__19766));
    Span4Mux_v I__4683 (
            .O(N__19788),
            .I(N__19763));
    LocalMux I__4682 (
            .O(N__19785),
            .I(N__19758));
    LocalMux I__4681 (
            .O(N__19782),
            .I(N__19758));
    InMux I__4680 (
            .O(N__19781),
            .I(N__19750));
    InMux I__4679 (
            .O(N__19780),
            .I(N__19750));
    InMux I__4678 (
            .O(N__19779),
            .I(N__19745));
    InMux I__4677 (
            .O(N__19778),
            .I(N__19745));
    LocalMux I__4676 (
            .O(N__19775),
            .I(N__19740));
    InMux I__4675 (
            .O(N__19774),
            .I(N__19736));
    LocalMux I__4674 (
            .O(N__19771),
            .I(N__19727));
    LocalMux I__4673 (
            .O(N__19766),
            .I(N__19727));
    Span4Mux_h I__4672 (
            .O(N__19763),
            .I(N__19727));
    Span4Mux_h I__4671 (
            .O(N__19758),
            .I(N__19727));
    InMux I__4670 (
            .O(N__19757),
            .I(N__19724));
    InMux I__4669 (
            .O(N__19756),
            .I(N__19721));
    InMux I__4668 (
            .O(N__19755),
            .I(N__19718));
    LocalMux I__4667 (
            .O(N__19750),
            .I(N__19713));
    LocalMux I__4666 (
            .O(N__19745),
            .I(N__19713));
    InMux I__4665 (
            .O(N__19744),
            .I(N__19708));
    InMux I__4664 (
            .O(N__19743),
            .I(N__19708));
    Span4Mux_v I__4663 (
            .O(N__19740),
            .I(N__19705));
    InMux I__4662 (
            .O(N__19739),
            .I(N__19702));
    LocalMux I__4661 (
            .O(N__19736),
            .I(N__19695));
    Span4Mux_v I__4660 (
            .O(N__19727),
            .I(N__19695));
    LocalMux I__4659 (
            .O(N__19724),
            .I(N__19695));
    LocalMux I__4658 (
            .O(N__19721),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4657 (
            .O(N__19718),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__4656 (
            .O(N__19713),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4655 (
            .O(N__19708),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__4654 (
            .O(N__19705),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    LocalMux I__4653 (
            .O(N__19702),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    Odrv4 I__4652 (
            .O(N__19695),
            .I(\Lab_UT.dictrl.stateZ0Z_2 ));
    CascadeMux I__4651 (
            .O(N__19680),
            .I(\Lab_UT.dictrl.g0_5_o4_4_cascade_ ));
    CascadeMux I__4650 (
            .O(N__19677),
            .I(N__19673));
    InMux I__4649 (
            .O(N__19676),
            .I(N__19666));
    InMux I__4648 (
            .O(N__19673),
            .I(N__19662));
    InMux I__4647 (
            .O(N__19672),
            .I(N__19659));
    InMux I__4646 (
            .O(N__19671),
            .I(N__19656));
    InMux I__4645 (
            .O(N__19670),
            .I(N__19651));
    InMux I__4644 (
            .O(N__19669),
            .I(N__19642));
    LocalMux I__4643 (
            .O(N__19666),
            .I(N__19638));
    InMux I__4642 (
            .O(N__19665),
            .I(N__19635));
    LocalMux I__4641 (
            .O(N__19662),
            .I(N__19632));
    LocalMux I__4640 (
            .O(N__19659),
            .I(N__19629));
    LocalMux I__4639 (
            .O(N__19656),
            .I(N__19626));
    InMux I__4638 (
            .O(N__19655),
            .I(N__19621));
    InMux I__4637 (
            .O(N__19654),
            .I(N__19621));
    LocalMux I__4636 (
            .O(N__19651),
            .I(N__19618));
    InMux I__4635 (
            .O(N__19650),
            .I(N__19615));
    InMux I__4634 (
            .O(N__19649),
            .I(N__19612));
    InMux I__4633 (
            .O(N__19648),
            .I(N__19609));
    InMux I__4632 (
            .O(N__19647),
            .I(N__19604));
    InMux I__4631 (
            .O(N__19646),
            .I(N__19604));
    InMux I__4630 (
            .O(N__19645),
            .I(N__19601));
    LocalMux I__4629 (
            .O(N__19642),
            .I(N__19598));
    InMux I__4628 (
            .O(N__19641),
            .I(N__19595));
    Span4Mux_h I__4627 (
            .O(N__19638),
            .I(N__19590));
    LocalMux I__4626 (
            .O(N__19635),
            .I(N__19590));
    Span4Mux_s3_h I__4625 (
            .O(N__19632),
            .I(N__19585));
    Span4Mux_v I__4624 (
            .O(N__19629),
            .I(N__19585));
    Span4Mux_v I__4623 (
            .O(N__19626),
            .I(N__19578));
    LocalMux I__4622 (
            .O(N__19621),
            .I(N__19578));
    Span4Mux_v I__4621 (
            .O(N__19618),
            .I(N__19578));
    LocalMux I__4620 (
            .O(N__19615),
            .I(N__19569));
    LocalMux I__4619 (
            .O(N__19612),
            .I(N__19569));
    LocalMux I__4618 (
            .O(N__19609),
            .I(N__19569));
    LocalMux I__4617 (
            .O(N__19604),
            .I(N__19569));
    LocalMux I__4616 (
            .O(N__19601),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__4615 (
            .O(N__19598),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    LocalMux I__4614 (
            .O(N__19595),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__4613 (
            .O(N__19590),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__4612 (
            .O(N__19585),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv4 I__4611 (
            .O(N__19578),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    Odrv12 I__4610 (
            .O(N__19569),
            .I(\Lab_UT.dictrl.stateZ0Z_1 ));
    InMux I__4609 (
            .O(N__19554),
            .I(N__19551));
    LocalMux I__4608 (
            .O(N__19551),
            .I(N__19548));
    Odrv4 I__4607 (
            .O(N__19548),
            .I(\Lab_UT.dictrl.N_11 ));
    InMux I__4606 (
            .O(N__19545),
            .I(N__19542));
    LocalMux I__4605 (
            .O(N__19542),
            .I(N__19539));
    Odrv4 I__4604 (
            .O(N__19539),
            .I(\buart.Z_rx.P7_mux ));
    InMux I__4603 (
            .O(N__19536),
            .I(N__19533));
    LocalMux I__4602 (
            .O(N__19533),
            .I(N_16_mux));
    CascadeMux I__4601 (
            .O(N__19530),
            .I(shifter_7_rep1_RNIG7Q01_cascade_));
    InMux I__4600 (
            .O(N__19527),
            .I(N__19524));
    LocalMux I__4599 (
            .O(N__19524),
            .I(N__19521));
    Span4Mux_h I__4598 (
            .O(N__19521),
            .I(N__19517));
    InMux I__4597 (
            .O(N__19520),
            .I(N__19514));
    Span4Mux_s3_h I__4596 (
            .O(N__19517),
            .I(N__19509));
    LocalMux I__4595 (
            .O(N__19514),
            .I(N__19509));
    Span4Mux_v I__4594 (
            .O(N__19509),
            .I(N__19506));
    Odrv4 I__4593 (
            .O(N__19506),
            .I(N_97));
    InMux I__4592 (
            .O(N__19503),
            .I(N__19500));
    LocalMux I__4591 (
            .O(N__19500),
            .I(N__19492));
    InMux I__4590 (
            .O(N__19499),
            .I(N__19489));
    InMux I__4589 (
            .O(N__19498),
            .I(N__19486));
    InMux I__4588 (
            .O(N__19497),
            .I(N__19483));
    InMux I__4587 (
            .O(N__19496),
            .I(N__19480));
    InMux I__4586 (
            .O(N__19495),
            .I(N__19477));
    Span4Mux_v I__4585 (
            .O(N__19492),
            .I(N__19472));
    LocalMux I__4584 (
            .O(N__19489),
            .I(N__19472));
    LocalMux I__4583 (
            .O(N__19486),
            .I(N__19469));
    LocalMux I__4582 (
            .O(N__19483),
            .I(N__19466));
    LocalMux I__4581 (
            .O(N__19480),
            .I(N__19461));
    LocalMux I__4580 (
            .O(N__19477),
            .I(N__19461));
    Span4Mux_h I__4579 (
            .O(N__19472),
            .I(N__19458));
    Sp12to4 I__4578 (
            .O(N__19469),
            .I(N__19455));
    Span4Mux_h I__4577 (
            .O(N__19466),
            .I(N__19452));
    Span4Mux_h I__4576 (
            .O(N__19461),
            .I(N__19449));
    Span4Mux_v I__4575 (
            .O(N__19458),
            .I(N__19446));
    Odrv12 I__4574 (
            .O(N__19455),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__4573 (
            .O(N__19452),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__4572 (
            .O(N__19449),
            .I(bu_rx_data_4_rep1));
    Odrv4 I__4571 (
            .O(N__19446),
            .I(bu_rx_data_4_rep1));
    IoInMux I__4570 (
            .O(N__19437),
            .I(N__19434));
    LocalMux I__4569 (
            .O(N__19434),
            .I(N__19431));
    Odrv4 I__4568 (
            .O(N__19431),
            .I(bu_rx_data_rdy_0));
    CascadeMux I__4567 (
            .O(N__19428),
            .I(N__19425));
    InMux I__4566 (
            .O(N__19425),
            .I(N__19422));
    LocalMux I__4565 (
            .O(N__19422),
            .I(N__19414));
    InMux I__4564 (
            .O(N__19421),
            .I(N__19409));
    InMux I__4563 (
            .O(N__19420),
            .I(N__19409));
    InMux I__4562 (
            .O(N__19419),
            .I(N__19404));
    InMux I__4561 (
            .O(N__19418),
            .I(N__19397));
    InMux I__4560 (
            .O(N__19417),
            .I(N__19397));
    Span4Mux_v I__4559 (
            .O(N__19414),
            .I(N__19390));
    LocalMux I__4558 (
            .O(N__19409),
            .I(N__19390));
    InMux I__4557 (
            .O(N__19408),
            .I(N__19385));
    InMux I__4556 (
            .O(N__19407),
            .I(N__19385));
    LocalMux I__4555 (
            .O(N__19404),
            .I(N__19382));
    InMux I__4554 (
            .O(N__19403),
            .I(N__19377));
    InMux I__4553 (
            .O(N__19402),
            .I(N__19377));
    LocalMux I__4552 (
            .O(N__19397),
            .I(N__19373));
    InMux I__4551 (
            .O(N__19396),
            .I(N__19370));
    InMux I__4550 (
            .O(N__19395),
            .I(N__19367));
    Span4Mux_h I__4549 (
            .O(N__19390),
            .I(N__19362));
    LocalMux I__4548 (
            .O(N__19385),
            .I(N__19362));
    Span4Mux_v I__4547 (
            .O(N__19382),
            .I(N__19357));
    LocalMux I__4546 (
            .O(N__19377),
            .I(N__19357));
    InMux I__4545 (
            .O(N__19376),
            .I(N__19354));
    Span12Mux_s6_v I__4544 (
            .O(N__19373),
            .I(N__19351));
    LocalMux I__4543 (
            .O(N__19370),
            .I(Lab_UT_dictrl_state_3_rep2));
    LocalMux I__4542 (
            .O(N__19367),
            .I(Lab_UT_dictrl_state_3_rep2));
    Odrv4 I__4541 (
            .O(N__19362),
            .I(Lab_UT_dictrl_state_3_rep2));
    Odrv4 I__4540 (
            .O(N__19357),
            .I(Lab_UT_dictrl_state_3_rep2));
    LocalMux I__4539 (
            .O(N__19354),
            .I(Lab_UT_dictrl_state_3_rep2));
    Odrv12 I__4538 (
            .O(N__19351),
            .I(Lab_UT_dictrl_state_3_rep2));
    CascadeMux I__4537 (
            .O(N__19338),
            .I(\Lab_UT.dictrl.g0_5_a4_1_5_cascade_ ));
    CascadeMux I__4536 (
            .O(N__19335),
            .I(\Lab_UT.dictrl.N_13_cascade_ ));
    InMux I__4535 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__4534 (
            .O(N__19329),
            .I(N__19326));
    Span4Mux_h I__4533 (
            .O(N__19326),
            .I(N__19323));
    Odrv4 I__4532 (
            .O(N__19323),
            .I(\Lab_UT.dictrl.N_90 ));
    CEMux I__4531 (
            .O(N__19320),
            .I(N__19296));
    CEMux I__4530 (
            .O(N__19319),
            .I(N__19296));
    CEMux I__4529 (
            .O(N__19318),
            .I(N__19296));
    CEMux I__4528 (
            .O(N__19317),
            .I(N__19296));
    CEMux I__4527 (
            .O(N__19316),
            .I(N__19296));
    CEMux I__4526 (
            .O(N__19315),
            .I(N__19296));
    CEMux I__4525 (
            .O(N__19314),
            .I(N__19296));
    CEMux I__4524 (
            .O(N__19313),
            .I(N__19296));
    GlobalMux I__4523 (
            .O(N__19296),
            .I(N__19293));
    gio2CtrlBuf I__4522 (
            .O(N__19293),
            .I(\buart.Z_rx.sample_g ));
    CascadeMux I__4521 (
            .O(N__19290),
            .I(N__19279));
    InMux I__4520 (
            .O(N__19289),
            .I(N__19275));
    InMux I__4519 (
            .O(N__19288),
            .I(N__19272));
    InMux I__4518 (
            .O(N__19287),
            .I(N__19269));
    InMux I__4517 (
            .O(N__19286),
            .I(N__19266));
    InMux I__4516 (
            .O(N__19285),
            .I(N__19263));
    InMux I__4515 (
            .O(N__19284),
            .I(N__19260));
    InMux I__4514 (
            .O(N__19283),
            .I(N__19257));
    InMux I__4513 (
            .O(N__19282),
            .I(N__19254));
    InMux I__4512 (
            .O(N__19279),
            .I(N__19251));
    InMux I__4511 (
            .O(N__19278),
            .I(N__19248));
    LocalMux I__4510 (
            .O(N__19275),
            .I(N__19245));
    LocalMux I__4509 (
            .O(N__19272),
            .I(N__19242));
    LocalMux I__4508 (
            .O(N__19269),
            .I(N__19196));
    LocalMux I__4507 (
            .O(N__19266),
            .I(N__19193));
    LocalMux I__4506 (
            .O(N__19263),
            .I(N__19190));
    LocalMux I__4505 (
            .O(N__19260),
            .I(N__19187));
    LocalMux I__4504 (
            .O(N__19257),
            .I(N__19184));
    LocalMux I__4503 (
            .O(N__19254),
            .I(N__19181));
    LocalMux I__4502 (
            .O(N__19251),
            .I(N__19163));
    LocalMux I__4501 (
            .O(N__19248),
            .I(N__19160));
    Glb2LocalMux I__4500 (
            .O(N__19245),
            .I(N__19023));
    Glb2LocalMux I__4499 (
            .O(N__19242),
            .I(N__19023));
    SRMux I__4498 (
            .O(N__19241),
            .I(N__19023));
    SRMux I__4497 (
            .O(N__19240),
            .I(N__19023));
    SRMux I__4496 (
            .O(N__19239),
            .I(N__19023));
    SRMux I__4495 (
            .O(N__19238),
            .I(N__19023));
    SRMux I__4494 (
            .O(N__19237),
            .I(N__19023));
    SRMux I__4493 (
            .O(N__19236),
            .I(N__19023));
    SRMux I__4492 (
            .O(N__19235),
            .I(N__19023));
    SRMux I__4491 (
            .O(N__19234),
            .I(N__19023));
    SRMux I__4490 (
            .O(N__19233),
            .I(N__19023));
    SRMux I__4489 (
            .O(N__19232),
            .I(N__19023));
    SRMux I__4488 (
            .O(N__19231),
            .I(N__19023));
    SRMux I__4487 (
            .O(N__19230),
            .I(N__19023));
    SRMux I__4486 (
            .O(N__19229),
            .I(N__19023));
    SRMux I__4485 (
            .O(N__19228),
            .I(N__19023));
    SRMux I__4484 (
            .O(N__19227),
            .I(N__19023));
    SRMux I__4483 (
            .O(N__19226),
            .I(N__19023));
    SRMux I__4482 (
            .O(N__19225),
            .I(N__19023));
    SRMux I__4481 (
            .O(N__19224),
            .I(N__19023));
    SRMux I__4480 (
            .O(N__19223),
            .I(N__19023));
    SRMux I__4479 (
            .O(N__19222),
            .I(N__19023));
    SRMux I__4478 (
            .O(N__19221),
            .I(N__19023));
    SRMux I__4477 (
            .O(N__19220),
            .I(N__19023));
    SRMux I__4476 (
            .O(N__19219),
            .I(N__19023));
    SRMux I__4475 (
            .O(N__19218),
            .I(N__19023));
    SRMux I__4474 (
            .O(N__19217),
            .I(N__19023));
    SRMux I__4473 (
            .O(N__19216),
            .I(N__19023));
    SRMux I__4472 (
            .O(N__19215),
            .I(N__19023));
    SRMux I__4471 (
            .O(N__19214),
            .I(N__19023));
    SRMux I__4470 (
            .O(N__19213),
            .I(N__19023));
    SRMux I__4469 (
            .O(N__19212),
            .I(N__19023));
    SRMux I__4468 (
            .O(N__19211),
            .I(N__19023));
    SRMux I__4467 (
            .O(N__19210),
            .I(N__19023));
    SRMux I__4466 (
            .O(N__19209),
            .I(N__19023));
    SRMux I__4465 (
            .O(N__19208),
            .I(N__19023));
    SRMux I__4464 (
            .O(N__19207),
            .I(N__19023));
    SRMux I__4463 (
            .O(N__19206),
            .I(N__19023));
    SRMux I__4462 (
            .O(N__19205),
            .I(N__19023));
    SRMux I__4461 (
            .O(N__19204),
            .I(N__19023));
    SRMux I__4460 (
            .O(N__19203),
            .I(N__19023));
    SRMux I__4459 (
            .O(N__19202),
            .I(N__19023));
    SRMux I__4458 (
            .O(N__19201),
            .I(N__19023));
    SRMux I__4457 (
            .O(N__19200),
            .I(N__19023));
    SRMux I__4456 (
            .O(N__19199),
            .I(N__19023));
    Glb2LocalMux I__4455 (
            .O(N__19196),
            .I(N__19023));
    Glb2LocalMux I__4454 (
            .O(N__19193),
            .I(N__19023));
    Glb2LocalMux I__4453 (
            .O(N__19190),
            .I(N__19023));
    Glb2LocalMux I__4452 (
            .O(N__19187),
            .I(N__19023));
    Glb2LocalMux I__4451 (
            .O(N__19184),
            .I(N__19023));
    Glb2LocalMux I__4450 (
            .O(N__19181),
            .I(N__19023));
    SRMux I__4449 (
            .O(N__19180),
            .I(N__19023));
    SRMux I__4448 (
            .O(N__19179),
            .I(N__19023));
    SRMux I__4447 (
            .O(N__19178),
            .I(N__19023));
    SRMux I__4446 (
            .O(N__19177),
            .I(N__19023));
    SRMux I__4445 (
            .O(N__19176),
            .I(N__19023));
    SRMux I__4444 (
            .O(N__19175),
            .I(N__19023));
    SRMux I__4443 (
            .O(N__19174),
            .I(N__19023));
    SRMux I__4442 (
            .O(N__19173),
            .I(N__19023));
    SRMux I__4441 (
            .O(N__19172),
            .I(N__19023));
    SRMux I__4440 (
            .O(N__19171),
            .I(N__19023));
    SRMux I__4439 (
            .O(N__19170),
            .I(N__19023));
    SRMux I__4438 (
            .O(N__19169),
            .I(N__19023));
    SRMux I__4437 (
            .O(N__19168),
            .I(N__19023));
    SRMux I__4436 (
            .O(N__19167),
            .I(N__19023));
    SRMux I__4435 (
            .O(N__19166),
            .I(N__19023));
    Glb2LocalMux I__4434 (
            .O(N__19163),
            .I(N__19023));
    Glb2LocalMux I__4433 (
            .O(N__19160),
            .I(N__19023));
    GlobalMux I__4432 (
            .O(N__19023),
            .I(N__19020));
    gio2CtrlBuf I__4431 (
            .O(N__19020),
            .I(rst_g));
    InMux I__4430 (
            .O(N__19017),
            .I(N__19014));
    LocalMux I__4429 (
            .O(N__19014),
            .I(N__19011));
    Span4Mux_v I__4428 (
            .O(N__19011),
            .I(N__19006));
    InMux I__4427 (
            .O(N__19010),
            .I(N__19003));
    InMux I__4426 (
            .O(N__19009),
            .I(N__19000));
    IoSpan4Mux I__4425 (
            .O(N__19006),
            .I(N__18994));
    LocalMux I__4424 (
            .O(N__19003),
            .I(N__18994));
    LocalMux I__4423 (
            .O(N__19000),
            .I(N__18991));
    InMux I__4422 (
            .O(N__18999),
            .I(N__18988));
    Span4Mux_s2_h I__4421 (
            .O(N__18994),
            .I(N__18983));
    Span4Mux_v I__4420 (
            .O(N__18991),
            .I(N__18980));
    LocalMux I__4419 (
            .O(N__18988),
            .I(N__18977));
    InMux I__4418 (
            .O(N__18987),
            .I(N__18972));
    InMux I__4417 (
            .O(N__18986),
            .I(N__18972));
    Span4Mux_h I__4416 (
            .O(N__18983),
            .I(N__18969));
    Odrv4 I__4415 (
            .O(N__18980),
            .I(bu_rx_data_rdy));
    Odrv12 I__4414 (
            .O(N__18977),
            .I(bu_rx_data_rdy));
    LocalMux I__4413 (
            .O(N__18972),
            .I(bu_rx_data_rdy));
    Odrv4 I__4412 (
            .O(N__18969),
            .I(bu_rx_data_rdy));
    CascadeMux I__4411 (
            .O(N__18960),
            .I(N__18957));
    InMux I__4410 (
            .O(N__18957),
            .I(N__18954));
    LocalMux I__4409 (
            .O(N__18954),
            .I(N__18951));
    Span4Mux_s1_h I__4408 (
            .O(N__18951),
            .I(N__18948));
    Odrv4 I__4407 (
            .O(N__18948),
            .I(\Lab_UT.dictrl.m25Z0Z_0 ));
    InMux I__4406 (
            .O(N__18945),
            .I(N__18937));
    InMux I__4405 (
            .O(N__18944),
            .I(N__18932));
    InMux I__4404 (
            .O(N__18943),
            .I(N__18932));
    InMux I__4403 (
            .O(N__18942),
            .I(N__18927));
    InMux I__4402 (
            .O(N__18941),
            .I(N__18927));
    InMux I__4401 (
            .O(N__18940),
            .I(N__18924));
    LocalMux I__4400 (
            .O(N__18937),
            .I(N__18917));
    LocalMux I__4399 (
            .O(N__18932),
            .I(N__18917));
    LocalMux I__4398 (
            .O(N__18927),
            .I(N__18917));
    LocalMux I__4397 (
            .O(N__18924),
            .I(bu_rx_data_fast_2));
    Odrv4 I__4396 (
            .O(N__18917),
            .I(bu_rx_data_fast_2));
    InMux I__4395 (
            .O(N__18912),
            .I(N__18905));
    InMux I__4394 (
            .O(N__18911),
            .I(N__18905));
    CascadeMux I__4393 (
            .O(N__18910),
            .I(N__18902));
    LocalMux I__4392 (
            .O(N__18905),
            .I(N__18896));
    InMux I__4391 (
            .O(N__18902),
            .I(N__18893));
    InMux I__4390 (
            .O(N__18901),
            .I(N__18886));
    InMux I__4389 (
            .O(N__18900),
            .I(N__18886));
    InMux I__4388 (
            .O(N__18899),
            .I(N__18886));
    Span4Mux_v I__4387 (
            .O(N__18896),
            .I(N__18879));
    LocalMux I__4386 (
            .O(N__18893),
            .I(N__18879));
    LocalMux I__4385 (
            .O(N__18886),
            .I(N__18879));
    Odrv4 I__4384 (
            .O(N__18879),
            .I(buart__rx_shifter_fast_5));
    InMux I__4383 (
            .O(N__18876),
            .I(N__18869));
    InMux I__4382 (
            .O(N__18875),
            .I(N__18869));
    InMux I__4381 (
            .O(N__18874),
            .I(N__18863));
    LocalMux I__4380 (
            .O(N__18869),
            .I(N__18860));
    InMux I__4379 (
            .O(N__18868),
            .I(N__18855));
    InMux I__4378 (
            .O(N__18867),
            .I(N__18855));
    CascadeMux I__4377 (
            .O(N__18866),
            .I(N__18847));
    LocalMux I__4376 (
            .O(N__18863),
            .I(N__18843));
    Span4Mux_h I__4375 (
            .O(N__18860),
            .I(N__18838));
    LocalMux I__4374 (
            .O(N__18855),
            .I(N__18838));
    InMux I__4373 (
            .O(N__18854),
            .I(N__18833));
    InMux I__4372 (
            .O(N__18853),
            .I(N__18833));
    InMux I__4371 (
            .O(N__18852),
            .I(N__18830));
    InMux I__4370 (
            .O(N__18851),
            .I(N__18827));
    InMux I__4369 (
            .O(N__18850),
            .I(N__18820));
    InMux I__4368 (
            .O(N__18847),
            .I(N__18820));
    InMux I__4367 (
            .O(N__18846),
            .I(N__18820));
    Span4Mux_v I__4366 (
            .O(N__18843),
            .I(N__18817));
    Span4Mux_h I__4365 (
            .O(N__18838),
            .I(N__18814));
    LocalMux I__4364 (
            .O(N__18833),
            .I(N__18811));
    LocalMux I__4363 (
            .O(N__18830),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4362 (
            .O(N__18827),
            .I(bu_rx_data_2_rep1));
    LocalMux I__4361 (
            .O(N__18820),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4360 (
            .O(N__18817),
            .I(bu_rx_data_2_rep1));
    Odrv4 I__4359 (
            .O(N__18814),
            .I(bu_rx_data_2_rep1));
    Odrv12 I__4358 (
            .O(N__18811),
            .I(bu_rx_data_2_rep1));
    InMux I__4357 (
            .O(N__18798),
            .I(N__18795));
    LocalMux I__4356 (
            .O(N__18795),
            .I(N__18792));
    Span4Mux_s3_h I__4355 (
            .O(N__18792),
            .I(N__18783));
    InMux I__4354 (
            .O(N__18791),
            .I(N__18780));
    InMux I__4353 (
            .O(N__18790),
            .I(N__18777));
    InMux I__4352 (
            .O(N__18789),
            .I(N__18772));
    InMux I__4351 (
            .O(N__18788),
            .I(N__18772));
    InMux I__4350 (
            .O(N__18787),
            .I(N__18767));
    InMux I__4349 (
            .O(N__18786),
            .I(N__18767));
    Odrv4 I__4348 (
            .O(N__18783),
            .I(\Lab_UT.dictrl.N_103_mux ));
    LocalMux I__4347 (
            .O(N__18780),
            .I(\Lab_UT.dictrl.N_103_mux ));
    LocalMux I__4346 (
            .O(N__18777),
            .I(\Lab_UT.dictrl.N_103_mux ));
    LocalMux I__4345 (
            .O(N__18772),
            .I(\Lab_UT.dictrl.N_103_mux ));
    LocalMux I__4344 (
            .O(N__18767),
            .I(\Lab_UT.dictrl.N_103_mux ));
    CascadeMux I__4343 (
            .O(N__18756),
            .I(\Lab_UT.dictrl.N_4_0_cascade_ ));
    InMux I__4342 (
            .O(N__18753),
            .I(N__18744));
    InMux I__4341 (
            .O(N__18752),
            .I(N__18739));
    InMux I__4340 (
            .O(N__18751),
            .I(N__18739));
    CascadeMux I__4339 (
            .O(N__18750),
            .I(N__18735));
    InMux I__4338 (
            .O(N__18749),
            .I(N__18730));
    InMux I__4337 (
            .O(N__18748),
            .I(N__18730));
    InMux I__4336 (
            .O(N__18747),
            .I(N__18727));
    LocalMux I__4335 (
            .O(N__18744),
            .I(N__18724));
    LocalMux I__4334 (
            .O(N__18739),
            .I(N__18721));
    InMux I__4333 (
            .O(N__18738),
            .I(N__18716));
    InMux I__4332 (
            .O(N__18735),
            .I(N__18713));
    LocalMux I__4331 (
            .O(N__18730),
            .I(N__18710));
    LocalMux I__4330 (
            .O(N__18727),
            .I(N__18703));
    Span4Mux_h I__4329 (
            .O(N__18724),
            .I(N__18703));
    Span4Mux_h I__4328 (
            .O(N__18721),
            .I(N__18703));
    InMux I__4327 (
            .O(N__18720),
            .I(N__18698));
    InMux I__4326 (
            .O(N__18719),
            .I(N__18698));
    LocalMux I__4325 (
            .O(N__18716),
            .I(N__18695));
    LocalMux I__4324 (
            .O(N__18713),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    Odrv4 I__4323 (
            .O(N__18710),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    Odrv4 I__4322 (
            .O(N__18703),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    LocalMux I__4321 (
            .O(N__18698),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    Odrv12 I__4320 (
            .O(N__18695),
            .I(\Lab_UT.dictrl.state_1_rep1 ));
    InMux I__4319 (
            .O(N__18684),
            .I(N__18681));
    LocalMux I__4318 (
            .O(N__18681),
            .I(N__18678));
    Span4Mux_h I__4317 (
            .O(N__18678),
            .I(N__18675));
    Odrv4 I__4316 (
            .O(N__18675),
            .I(\Lab_UT.dictrl.N_12_0 ));
    InMux I__4315 (
            .O(N__18672),
            .I(N__18669));
    LocalMux I__4314 (
            .O(N__18669),
            .I(N__18666));
    Odrv12 I__4313 (
            .O(N__18666),
            .I(\Lab_UT.LdASones ));
    CEMux I__4312 (
            .O(N__18663),
            .I(N__18659));
    CEMux I__4311 (
            .O(N__18662),
            .I(N__18656));
    LocalMux I__4310 (
            .O(N__18659),
            .I(N__18653));
    LocalMux I__4309 (
            .O(N__18656),
            .I(N__18650));
    Sp12to4 I__4308 (
            .O(N__18653),
            .I(N__18647));
    Span4Mux_v I__4307 (
            .O(N__18650),
            .I(N__18644));
    Span12Mux_v I__4306 (
            .O(N__18647),
            .I(N__18641));
    Span4Mux_v I__4305 (
            .O(N__18644),
            .I(N__18638));
    Odrv12 I__4304 (
            .O(N__18641),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    Odrv4 I__4303 (
            .O(N__18638),
            .I(\Lab_UT.didp.regrce1.LdASones_0 ));
    CascadeMux I__4302 (
            .O(N__18633),
            .I(N__18629));
    CascadeMux I__4301 (
            .O(N__18632),
            .I(N__18624));
    InMux I__4300 (
            .O(N__18629),
            .I(N__18621));
    CascadeMux I__4299 (
            .O(N__18628),
            .I(N__18618));
    InMux I__4298 (
            .O(N__18627),
            .I(N__18615));
    InMux I__4297 (
            .O(N__18624),
            .I(N__18612));
    LocalMux I__4296 (
            .O(N__18621),
            .I(N__18609));
    InMux I__4295 (
            .O(N__18618),
            .I(N__18606));
    LocalMux I__4294 (
            .O(N__18615),
            .I(N__18602));
    LocalMux I__4293 (
            .O(N__18612),
            .I(N__18599));
    Span4Mux_h I__4292 (
            .O(N__18609),
            .I(N__18594));
    LocalMux I__4291 (
            .O(N__18606),
            .I(N__18594));
    CascadeMux I__4290 (
            .O(N__18605),
            .I(N__18591));
    Span12Mux_s5_h I__4289 (
            .O(N__18602),
            .I(N__18588));
    Span4Mux_h I__4288 (
            .O(N__18599),
            .I(N__18585));
    Span4Mux_v I__4287 (
            .O(N__18594),
            .I(N__18582));
    InMux I__4286 (
            .O(N__18591),
            .I(N__18579));
    Odrv12 I__4285 (
            .O(N__18588),
            .I(bu_rx_data_7_rep1));
    Odrv4 I__4284 (
            .O(N__18585),
            .I(bu_rx_data_7_rep1));
    Odrv4 I__4283 (
            .O(N__18582),
            .I(bu_rx_data_7_rep1));
    LocalMux I__4282 (
            .O(N__18579),
            .I(bu_rx_data_7_rep1));
    InMux I__4281 (
            .O(N__18570),
            .I(N__18567));
    LocalMux I__4280 (
            .O(N__18567),
            .I(shifter_7_rep1_RNIG7Q01));
    CascadeMux I__4279 (
            .O(N__18564),
            .I(\Lab_UT.dictrl.N_77_cascade_ ));
    InMux I__4278 (
            .O(N__18561),
            .I(N__18558));
    LocalMux I__4277 (
            .O(N__18558),
            .I(N__18555));
    Odrv4 I__4276 (
            .O(N__18555),
            .I(\Lab_UT.dictrl.m73Z0Z_1 ));
    InMux I__4275 (
            .O(N__18552),
            .I(N__18549));
    LocalMux I__4274 (
            .O(N__18549),
            .I(\Lab_UT.dictrl.m77_ns_1 ));
    CascadeMux I__4273 (
            .O(N__18546),
            .I(\Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_ ));
    InMux I__4272 (
            .O(N__18543),
            .I(N__18539));
    InMux I__4271 (
            .O(N__18542),
            .I(N__18536));
    LocalMux I__4270 (
            .O(N__18539),
            .I(N__18533));
    LocalMux I__4269 (
            .O(N__18536),
            .I(N__18530));
    Span4Mux_h I__4268 (
            .O(N__18533),
            .I(N__18527));
    Odrv4 I__4267 (
            .O(N__18530),
            .I(\Lab_UT.dictrl.i9_mux_0_0 ));
    Odrv4 I__4266 (
            .O(N__18527),
            .I(\Lab_UT.dictrl.i9_mux_0_0 ));
    InMux I__4265 (
            .O(N__18522),
            .I(N__18516));
    InMux I__4264 (
            .O(N__18521),
            .I(N__18516));
    LocalMux I__4263 (
            .O(N__18516),
            .I(N__18512));
    InMux I__4262 (
            .O(N__18515),
            .I(N__18509));
    Odrv4 I__4261 (
            .O(N__18512),
            .I(\Lab_UT.dictrl.N_106_mux ));
    LocalMux I__4260 (
            .O(N__18509),
            .I(\Lab_UT.dictrl.N_106_mux ));
    InMux I__4259 (
            .O(N__18504),
            .I(N__18501));
    LocalMux I__4258 (
            .O(N__18501),
            .I(N__18498));
    Odrv4 I__4257 (
            .O(N__18498),
            .I(\Lab_UT.dictrl.m51_0 ));
    InMux I__4256 (
            .O(N__18495),
            .I(N__18490));
    InMux I__4255 (
            .O(N__18494),
            .I(N__18487));
    InMux I__4254 (
            .O(N__18493),
            .I(N__18484));
    LocalMux I__4253 (
            .O(N__18490),
            .I(N__18481));
    LocalMux I__4252 (
            .O(N__18487),
            .I(N__18478));
    LocalMux I__4251 (
            .O(N__18484),
            .I(N__18472));
    Span4Mux_v I__4250 (
            .O(N__18481),
            .I(N__18472));
    Span4Mux_v I__4249 (
            .O(N__18478),
            .I(N__18469));
    CascadeMux I__4248 (
            .O(N__18477),
            .I(N__18466));
    Span4Mux_v I__4247 (
            .O(N__18472),
            .I(N__18461));
    Span4Mux_v I__4246 (
            .O(N__18469),
            .I(N__18461));
    InMux I__4245 (
            .O(N__18466),
            .I(N__18458));
    Odrv4 I__4244 (
            .O(N__18461),
            .I(\Lab_UT.dictrl.state_i_3_1 ));
    LocalMux I__4243 (
            .O(N__18458),
            .I(\Lab_UT.dictrl.state_i_3_1 ));
    CascadeMux I__4242 (
            .O(N__18453),
            .I(\Lab_UT.dictrl.N_118_mux_cascade_ ));
    InMux I__4241 (
            .O(N__18450),
            .I(N__18447));
    LocalMux I__4240 (
            .O(N__18447),
            .I(N__18444));
    Odrv4 I__4239 (
            .O(N__18444),
            .I(\Lab_UT.dictrl.next_state_latmux_3_1_1 ));
    InMux I__4238 (
            .O(N__18441),
            .I(N__18438));
    LocalMux I__4237 (
            .O(N__18438),
            .I(N__18435));
    Span4Mux_h I__4236 (
            .O(N__18435),
            .I(N__18432));
    Odrv4 I__4235 (
            .O(N__18432),
            .I(\Lab_UT.dictrl.g0_17_a6_3Z0Z_7 ));
    CascadeMux I__4234 (
            .O(N__18429),
            .I(N__18425));
    InMux I__4233 (
            .O(N__18428),
            .I(N__18420));
    InMux I__4232 (
            .O(N__18425),
            .I(N__18414));
    InMux I__4231 (
            .O(N__18424),
            .I(N__18414));
    InMux I__4230 (
            .O(N__18423),
            .I(N__18411));
    LocalMux I__4229 (
            .O(N__18420),
            .I(N__18408));
    InMux I__4228 (
            .O(N__18419),
            .I(N__18405));
    LocalMux I__4227 (
            .O(N__18414),
            .I(N__18402));
    LocalMux I__4226 (
            .O(N__18411),
            .I(N__18399));
    Span4Mux_h I__4225 (
            .O(N__18408),
            .I(N__18396));
    LocalMux I__4224 (
            .O(N__18405),
            .I(N__18391));
    Span4Mux_h I__4223 (
            .O(N__18402),
            .I(N__18391));
    Odrv4 I__4222 (
            .O(N__18399),
            .I(buart__rx_shifter_fast_0));
    Odrv4 I__4221 (
            .O(N__18396),
            .I(buart__rx_shifter_fast_0));
    Odrv4 I__4220 (
            .O(N__18391),
            .I(buart__rx_shifter_fast_0));
    CascadeMux I__4219 (
            .O(N__18384),
            .I(N__18376));
    InMux I__4218 (
            .O(N__18383),
            .I(N__18370));
    InMux I__4217 (
            .O(N__18382),
            .I(N__18370));
    InMux I__4216 (
            .O(N__18381),
            .I(N__18365));
    InMux I__4215 (
            .O(N__18380),
            .I(N__18365));
    InMux I__4214 (
            .O(N__18379),
            .I(N__18362));
    InMux I__4213 (
            .O(N__18376),
            .I(N__18359));
    InMux I__4212 (
            .O(N__18375),
            .I(N__18356));
    LocalMux I__4211 (
            .O(N__18370),
            .I(N__18348));
    LocalMux I__4210 (
            .O(N__18365),
            .I(N__18348));
    LocalMux I__4209 (
            .O(N__18362),
            .I(N__18343));
    LocalMux I__4208 (
            .O(N__18359),
            .I(N__18343));
    LocalMux I__4207 (
            .O(N__18356),
            .I(N__18340));
    InMux I__4206 (
            .O(N__18355),
            .I(N__18337));
    InMux I__4205 (
            .O(N__18354),
            .I(N__18332));
    InMux I__4204 (
            .O(N__18353),
            .I(N__18332));
    Span4Mux_h I__4203 (
            .O(N__18348),
            .I(N__18329));
    Span4Mux_s3_h I__4202 (
            .O(N__18343),
            .I(N__18326));
    Odrv4 I__4201 (
            .O(N__18340),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4200 (
            .O(N__18337),
            .I(bu_rx_data_1_rep1));
    LocalMux I__4199 (
            .O(N__18332),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__4198 (
            .O(N__18329),
            .I(bu_rx_data_1_rep1));
    Odrv4 I__4197 (
            .O(N__18326),
            .I(bu_rx_data_1_rep1));
    CascadeMux I__4196 (
            .O(N__18315),
            .I(N__18311));
    InMux I__4195 (
            .O(N__18314),
            .I(N__18303));
    InMux I__4194 (
            .O(N__18311),
            .I(N__18303));
    InMux I__4193 (
            .O(N__18310),
            .I(N__18303));
    LocalMux I__4192 (
            .O(N__18303),
            .I(N__18299));
    InMux I__4191 (
            .O(N__18302),
            .I(N__18294));
    Span4Mux_v I__4190 (
            .O(N__18299),
            .I(N__18291));
    CascadeMux I__4189 (
            .O(N__18298),
            .I(N__18288));
    InMux I__4188 (
            .O(N__18297),
            .I(N__18283));
    LocalMux I__4187 (
            .O(N__18294),
            .I(N__18278));
    Sp12to4 I__4186 (
            .O(N__18291),
            .I(N__18278));
    InMux I__4185 (
            .O(N__18288),
            .I(N__18271));
    InMux I__4184 (
            .O(N__18287),
            .I(N__18271));
    InMux I__4183 (
            .O(N__18286),
            .I(N__18271));
    LocalMux I__4182 (
            .O(N__18283),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    Odrv12 I__4181 (
            .O(N__18278),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    LocalMux I__4180 (
            .O(N__18271),
            .I(\Lab_UT.dictrl.next_state_1_3 ));
    InMux I__4179 (
            .O(N__18264),
            .I(N__18261));
    LocalMux I__4178 (
            .O(N__18261),
            .I(\Lab_UT.dictrl.P6_mux_0 ));
    CascadeMux I__4177 (
            .O(N__18258),
            .I(N__18254));
    InMux I__4176 (
            .O(N__18257),
            .I(N__18250));
    InMux I__4175 (
            .O(N__18254),
            .I(N__18247));
    InMux I__4174 (
            .O(N__18253),
            .I(N__18244));
    LocalMux I__4173 (
            .O(N__18250),
            .I(N__18241));
    LocalMux I__4172 (
            .O(N__18247),
            .I(N__18238));
    LocalMux I__4171 (
            .O(N__18244),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv4 I__4170 (
            .O(N__18241),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    Odrv4 I__4169 (
            .O(N__18238),
            .I(\Lab_UT.dictrl.state_i_3_2 ));
    CascadeMux I__4168 (
            .O(N__18231),
            .I(N__18228));
    InMux I__4167 (
            .O(N__18228),
            .I(N__18225));
    LocalMux I__4166 (
            .O(N__18225),
            .I(N__18222));
    Odrv4 I__4165 (
            .O(N__18222),
            .I(\Lab_UT.dictrl.N_114_mux ));
    InMux I__4164 (
            .O(N__18219),
            .I(N__18216));
    LocalMux I__4163 (
            .O(N__18216),
            .I(\Lab_UT.dictrl.N_69 ));
    CascadeMux I__4162 (
            .O(N__18213),
            .I(N__18209));
    InMux I__4161 (
            .O(N__18212),
            .I(N__18204));
    InMux I__4160 (
            .O(N__18209),
            .I(N__18204));
    LocalMux I__4159 (
            .O(N__18204),
            .I(\Lab_UT.dictrl.i10_mux ));
    CascadeMux I__4158 (
            .O(N__18201),
            .I(\Lab_UT.dictrl.N_69_cascade_ ));
    InMux I__4157 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__4156 (
            .O(N__18195),
            .I(N__18192));
    Span4Mux_v I__4155 (
            .O(N__18192),
            .I(N__18189));
    Odrv4 I__4154 (
            .O(N__18189),
            .I(\Lab_UT.dictrl.next_state_1_0_3 ));
    InMux I__4153 (
            .O(N__18186),
            .I(N__18183));
    LocalMux I__4152 (
            .O(N__18183),
            .I(N__18180));
    Odrv4 I__4151 (
            .O(N__18180),
            .I(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1 ));
    CascadeMux I__4150 (
            .O(N__18177),
            .I(N__18171));
    CascadeMux I__4149 (
            .O(N__18176),
            .I(N__18168));
    CascadeMux I__4148 (
            .O(N__18175),
            .I(N__18165));
    InMux I__4147 (
            .O(N__18174),
            .I(N__18158));
    InMux I__4146 (
            .O(N__18171),
            .I(N__18158));
    InMux I__4145 (
            .O(N__18168),
            .I(N__18158));
    InMux I__4144 (
            .O(N__18165),
            .I(N__18155));
    LocalMux I__4143 (
            .O(N__18158),
            .I(N__18150));
    LocalMux I__4142 (
            .O(N__18155),
            .I(N__18150));
    Span4Mux_h I__4141 (
            .O(N__18150),
            .I(N__18147));
    Odrv4 I__4140 (
            .O(N__18147),
            .I(\Lab_UT.dictrl.g0_17_a6_0_1 ));
    CascadeMux I__4139 (
            .O(N__18144),
            .I(N__18141));
    InMux I__4138 (
            .O(N__18141),
            .I(N__18138));
    LocalMux I__4137 (
            .O(N__18138),
            .I(\Lab_UT.dictrl.P6_mux ));
    InMux I__4136 (
            .O(N__18135),
            .I(N__18128));
    InMux I__4135 (
            .O(N__18134),
            .I(N__18128));
    InMux I__4134 (
            .O(N__18133),
            .I(N__18125));
    LocalMux I__4133 (
            .O(N__18128),
            .I(N__18122));
    LocalMux I__4132 (
            .O(N__18125),
            .I(N__18119));
    Span4Mux_h I__4131 (
            .O(N__18122),
            .I(N__18116));
    Span4Mux_h I__4130 (
            .O(N__18119),
            .I(N__18113));
    Odrv4 I__4129 (
            .O(N__18116),
            .I(\Lab_UT.dictrl.N_189 ));
    Odrv4 I__4128 (
            .O(N__18113),
            .I(\Lab_UT.dictrl.N_189 ));
    CascadeMux I__4127 (
            .O(N__18108),
            .I(N__18105));
    InMux I__4126 (
            .O(N__18105),
            .I(N__18098));
    InMux I__4125 (
            .O(N__18104),
            .I(N__18098));
    InMux I__4124 (
            .O(N__18103),
            .I(N__18095));
    LocalMux I__4123 (
            .O(N__18098),
            .I(\Lab_UT.dictrl.m40_N_5_mux ));
    LocalMux I__4122 (
            .O(N__18095),
            .I(\Lab_UT.dictrl.m40_N_5_mux ));
    InMux I__4121 (
            .O(N__18090),
            .I(N__18086));
    InMux I__4120 (
            .O(N__18089),
            .I(N__18083));
    LocalMux I__4119 (
            .O(N__18086),
            .I(\Lab_UT.dictrl.N_77 ));
    LocalMux I__4118 (
            .O(N__18083),
            .I(\Lab_UT.dictrl.N_77 ));
    InMux I__4117 (
            .O(N__18078),
            .I(N__18072));
    InMux I__4116 (
            .O(N__18077),
            .I(N__18072));
    LocalMux I__4115 (
            .O(N__18072),
            .I(\Lab_UT.dictrl.alarmstate8Z0Z_4 ));
    InMux I__4114 (
            .O(N__18069),
            .I(N__18065));
    CascadeMux I__4113 (
            .O(N__18068),
            .I(N__18062));
    LocalMux I__4112 (
            .O(N__18065),
            .I(N__18057));
    InMux I__4111 (
            .O(N__18062),
            .I(N__18054));
    InMux I__4110 (
            .O(N__18061),
            .I(N__18051));
    InMux I__4109 (
            .O(N__18060),
            .I(N__18048));
    Span4Mux_s3_h I__4108 (
            .O(N__18057),
            .I(N__18041));
    LocalMux I__4107 (
            .O(N__18054),
            .I(N__18041));
    LocalMux I__4106 (
            .O(N__18051),
            .I(N__18036));
    LocalMux I__4105 (
            .O(N__18048),
            .I(N__18036));
    InMux I__4104 (
            .O(N__18047),
            .I(N__18029));
    InMux I__4103 (
            .O(N__18046),
            .I(N__18029));
    Span4Mux_h I__4102 (
            .O(N__18041),
            .I(N__18026));
    Span4Mux_v I__4101 (
            .O(N__18036),
            .I(N__18023));
    InMux I__4100 (
            .O(N__18035),
            .I(N__18020));
    InMux I__4099 (
            .O(N__18034),
            .I(N__18017));
    LocalMux I__4098 (
            .O(N__18029),
            .I(\Lab_UT.didp.di_Sones_0 ));
    Odrv4 I__4097 (
            .O(N__18026),
            .I(\Lab_UT.didp.di_Sones_0 ));
    Odrv4 I__4096 (
            .O(N__18023),
            .I(\Lab_UT.didp.di_Sones_0 ));
    LocalMux I__4095 (
            .O(N__18020),
            .I(\Lab_UT.didp.di_Sones_0 ));
    LocalMux I__4094 (
            .O(N__18017),
            .I(\Lab_UT.didp.di_Sones_0 ));
    InMux I__4093 (
            .O(N__18006),
            .I(N__18003));
    LocalMux I__4092 (
            .O(N__18003),
            .I(N__17999));
    CascadeMux I__4091 (
            .O(N__18002),
            .I(N__17995));
    Span4Mux_h I__4090 (
            .O(N__17999),
            .I(N__17991));
    InMux I__4089 (
            .O(N__17998),
            .I(N__17988));
    InMux I__4088 (
            .O(N__17995),
            .I(N__17985));
    CascadeMux I__4087 (
            .O(N__17994),
            .I(N__17982));
    Span4Mux_h I__4086 (
            .O(N__17991),
            .I(N__17977));
    LocalMux I__4085 (
            .O(N__17988),
            .I(N__17977));
    LocalMux I__4084 (
            .O(N__17985),
            .I(N__17974));
    InMux I__4083 (
            .O(N__17982),
            .I(N__17971));
    Odrv4 I__4082 (
            .O(N__17977),
            .I(\Lab_UT.LdSones ));
    Odrv4 I__4081 (
            .O(N__17974),
            .I(\Lab_UT.LdSones ));
    LocalMux I__4080 (
            .O(N__17971),
            .I(\Lab_UT.LdSones ));
    InMux I__4079 (
            .O(N__17964),
            .I(N__17961));
    LocalMux I__4078 (
            .O(N__17961),
            .I(N__17957));
    CascadeMux I__4077 (
            .O(N__17960),
            .I(N__17953));
    Span4Mux_h I__4076 (
            .O(N__17957),
            .I(N__17946));
    CascadeMux I__4075 (
            .O(N__17956),
            .I(N__17943));
    InMux I__4074 (
            .O(N__17953),
            .I(N__17940));
    InMux I__4073 (
            .O(N__17952),
            .I(N__17937));
    InMux I__4072 (
            .O(N__17951),
            .I(N__17932));
    InMux I__4071 (
            .O(N__17950),
            .I(N__17932));
    InMux I__4070 (
            .O(N__17949),
            .I(N__17929));
    Span4Mux_s3_h I__4069 (
            .O(N__17946),
            .I(N__17926));
    InMux I__4068 (
            .O(N__17943),
            .I(N__17923));
    LocalMux I__4067 (
            .O(N__17940),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__4066 (
            .O(N__17937),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__4065 (
            .O(N__17932),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__4064 (
            .O(N__17929),
            .I(\Lab_UT.didp.di_Sones_1 ));
    Odrv4 I__4063 (
            .O(N__17926),
            .I(\Lab_UT.didp.di_Sones_1 ));
    LocalMux I__4062 (
            .O(N__17923),
            .I(\Lab_UT.didp.di_Sones_1 ));
    InMux I__4061 (
            .O(N__17910),
            .I(N__17907));
    LocalMux I__4060 (
            .O(N__17907),
            .I(\Lab_UT.didp.countrce1.q_5_1 ));
    CascadeMux I__4059 (
            .O(N__17904),
            .I(\Lab_UT.dictrl.N_4_cascade_ ));
    InMux I__4058 (
            .O(N__17901),
            .I(N__17898));
    LocalMux I__4057 (
            .O(N__17898),
            .I(N__17892));
    InMux I__4056 (
            .O(N__17897),
            .I(N__17885));
    InMux I__4055 (
            .O(N__17896),
            .I(N__17885));
    InMux I__4054 (
            .O(N__17895),
            .I(N__17885));
    Span4Mux_h I__4053 (
            .O(N__17892),
            .I(N__17882));
    LocalMux I__4052 (
            .O(N__17885),
            .I(\Lab_UT.dictrl.N_12 ));
    Odrv4 I__4051 (
            .O(N__17882),
            .I(\Lab_UT.dictrl.N_12 ));
    InMux I__4050 (
            .O(N__17877),
            .I(N__17873));
    CascadeMux I__4049 (
            .O(N__17876),
            .I(N__17870));
    LocalMux I__4048 (
            .O(N__17873),
            .I(N__17867));
    InMux I__4047 (
            .O(N__17870),
            .I(N__17864));
    Odrv12 I__4046 (
            .O(N__17867),
            .I(\Lab_UT.dictrl.N_81 ));
    LocalMux I__4045 (
            .O(N__17864),
            .I(\Lab_UT.dictrl.N_81 ));
    InMux I__4044 (
            .O(N__17859),
            .I(N__17856));
    LocalMux I__4043 (
            .O(N__17856),
            .I(\Lab_UT.dictrl.next_state_i_1_2 ));
    CascadeMux I__4042 (
            .O(N__17853),
            .I(N__17850));
    InMux I__4041 (
            .O(N__17850),
            .I(N__17847));
    LocalMux I__4040 (
            .O(N__17847),
            .I(N__17844));
    Span4Mux_v I__4039 (
            .O(N__17844),
            .I(N__17841));
    Span4Mux_v I__4038 (
            .O(N__17841),
            .I(N__17838));
    Odrv4 I__4037 (
            .O(N__17838),
            .I(\Lab_UT.dictrl.P8_mux ));
    InMux I__4036 (
            .O(N__17835),
            .I(N__17831));
    InMux I__4035 (
            .O(N__17834),
            .I(N__17828));
    LocalMux I__4034 (
            .O(N__17831),
            .I(N__17821));
    LocalMux I__4033 (
            .O(N__17828),
            .I(N__17816));
    InMux I__4032 (
            .O(N__17827),
            .I(N__17810));
    InMux I__4031 (
            .O(N__17826),
            .I(N__17807));
    InMux I__4030 (
            .O(N__17825),
            .I(N__17802));
    InMux I__4029 (
            .O(N__17824),
            .I(N__17802));
    Span4Mux_v I__4028 (
            .O(N__17821),
            .I(N__17799));
    InMux I__4027 (
            .O(N__17820),
            .I(N__17794));
    InMux I__4026 (
            .O(N__17819),
            .I(N__17794));
    Span4Mux_h I__4025 (
            .O(N__17816),
            .I(N__17791));
    InMux I__4024 (
            .O(N__17815),
            .I(N__17784));
    InMux I__4023 (
            .O(N__17814),
            .I(N__17784));
    InMux I__4022 (
            .O(N__17813),
            .I(N__17784));
    LocalMux I__4021 (
            .O(N__17810),
            .I(G_183));
    LocalMux I__4020 (
            .O(N__17807),
            .I(G_183));
    LocalMux I__4019 (
            .O(N__17802),
            .I(G_183));
    Odrv4 I__4018 (
            .O(N__17799),
            .I(G_183));
    LocalMux I__4017 (
            .O(N__17794),
            .I(G_183));
    Odrv4 I__4016 (
            .O(N__17791),
            .I(G_183));
    LocalMux I__4015 (
            .O(N__17784),
            .I(G_183));
    InMux I__4014 (
            .O(N__17769),
            .I(N__17764));
    InMux I__4013 (
            .O(N__17768),
            .I(N__17758));
    InMux I__4012 (
            .O(N__17767),
            .I(N__17752));
    LocalMux I__4011 (
            .O(N__17764),
            .I(N__17749));
    InMux I__4010 (
            .O(N__17763),
            .I(N__17742));
    InMux I__4009 (
            .O(N__17762),
            .I(N__17742));
    InMux I__4008 (
            .O(N__17761),
            .I(N__17742));
    LocalMux I__4007 (
            .O(N__17758),
            .I(N__17739));
    InMux I__4006 (
            .O(N__17757),
            .I(N__17731));
    InMux I__4005 (
            .O(N__17756),
            .I(N__17731));
    InMux I__4004 (
            .O(N__17755),
            .I(N__17728));
    LocalMux I__4003 (
            .O(N__17752),
            .I(N__17719));
    Span4Mux_h I__4002 (
            .O(N__17749),
            .I(N__17719));
    LocalMux I__4001 (
            .O(N__17742),
            .I(N__17719));
    Span4Mux_v I__4000 (
            .O(N__17739),
            .I(N__17719));
    InMux I__3999 (
            .O(N__17738),
            .I(N__17712));
    InMux I__3998 (
            .O(N__17737),
            .I(N__17712));
    InMux I__3997 (
            .O(N__17736),
            .I(N__17712));
    LocalMux I__3996 (
            .O(N__17731),
            .I(G_185));
    LocalMux I__3995 (
            .O(N__17728),
            .I(G_185));
    Odrv4 I__3994 (
            .O(N__17719),
            .I(G_185));
    LocalMux I__3993 (
            .O(N__17712),
            .I(G_185));
    CascadeMux I__3992 (
            .O(N__17703),
            .I(\Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ));
    InMux I__3991 (
            .O(N__17700),
            .I(N__17697));
    LocalMux I__3990 (
            .O(N__17697),
            .I(\Lab_UT.dictrl.m3_0 ));
    CascadeMux I__3989 (
            .O(N__17694),
            .I(\Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_ ));
    InMux I__3988 (
            .O(N__17691),
            .I(N__17688));
    LocalMux I__3987 (
            .O(N__17688),
            .I(G_188));
    InMux I__3986 (
            .O(N__17685),
            .I(N__17682));
    LocalMux I__3985 (
            .O(N__17682),
            .I(\Lab_UT.dictrl.alarmstate8Z0Z_3 ));
    CascadeMux I__3984 (
            .O(N__17679),
            .I(G_188_cascade_));
    InMux I__3983 (
            .O(N__17676),
            .I(N__17673));
    LocalMux I__3982 (
            .O(N__17673),
            .I(G_187));
    CascadeMux I__3981 (
            .O(N__17670),
            .I(N__17666));
    InMux I__3980 (
            .O(N__17669),
            .I(N__17661));
    InMux I__3979 (
            .O(N__17666),
            .I(N__17661));
    LocalMux I__3978 (
            .O(N__17661),
            .I(N__17658));
    Odrv12 I__3977 (
            .O(N__17658),
            .I(G_186));
    CascadeMux I__3976 (
            .O(N__17655),
            .I(G_187_cascade_));
    InMux I__3975 (
            .O(N__17652),
            .I(N__17643));
    InMux I__3974 (
            .O(N__17651),
            .I(N__17643));
    InMux I__3973 (
            .O(N__17650),
            .I(N__17643));
    LocalMux I__3972 (
            .O(N__17643),
            .I(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ));
    InMux I__3971 (
            .O(N__17640),
            .I(N__17637));
    LocalMux I__3970 (
            .O(N__17637),
            .I(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ));
    InMux I__3969 (
            .O(N__17634),
            .I(N__17625));
    InMux I__3968 (
            .O(N__17633),
            .I(N__17616));
    InMux I__3967 (
            .O(N__17632),
            .I(N__17616));
    InMux I__3966 (
            .O(N__17631),
            .I(N__17616));
    InMux I__3965 (
            .O(N__17630),
            .I(N__17616));
    CascadeMux I__3964 (
            .O(N__17629),
            .I(N__17613));
    CascadeMux I__3963 (
            .O(N__17628),
            .I(N__17610));
    LocalMux I__3962 (
            .O(N__17625),
            .I(N__17607));
    LocalMux I__3961 (
            .O(N__17616),
            .I(N__17604));
    InMux I__3960 (
            .O(N__17613),
            .I(N__17601));
    InMux I__3959 (
            .O(N__17610),
            .I(N__17598));
    Odrv4 I__3958 (
            .O(N__17607),
            .I(\Lab_UT.state_i_3_0 ));
    Odrv4 I__3957 (
            .O(N__17604),
            .I(\Lab_UT.state_i_3_0 ));
    LocalMux I__3956 (
            .O(N__17601),
            .I(\Lab_UT.state_i_3_0 ));
    LocalMux I__3955 (
            .O(N__17598),
            .I(\Lab_UT.state_i_3_0 ));
    CascadeMux I__3954 (
            .O(N__17589),
            .I(\Lab_UT.dictrl.g0_2Z0Z_2_cascade_ ));
    InMux I__3953 (
            .O(N__17586),
            .I(N__17583));
    LocalMux I__3952 (
            .O(N__17583),
            .I(N__17580));
    Odrv4 I__3951 (
            .O(N__17580),
            .I(\Lab_UT.dictrl.m40_N_5_mux_1 ));
    InMux I__3950 (
            .O(N__17577),
            .I(N__17574));
    LocalMux I__3949 (
            .O(N__17574),
            .I(N__17570));
    InMux I__3948 (
            .O(N__17573),
            .I(N__17567));
    Span4Mux_v I__3947 (
            .O(N__17570),
            .I(N__17561));
    LocalMux I__3946 (
            .O(N__17567),
            .I(N__17561));
    InMux I__3945 (
            .O(N__17566),
            .I(N__17557));
    Span4Mux_h I__3944 (
            .O(N__17561),
            .I(N__17554));
    InMux I__3943 (
            .O(N__17560),
            .I(N__17551));
    LocalMux I__3942 (
            .O(N__17557),
            .I(\Lab_UT.di_AStens_2 ));
    Odrv4 I__3941 (
            .O(N__17554),
            .I(\Lab_UT.di_AStens_2 ));
    LocalMux I__3940 (
            .O(N__17551),
            .I(\Lab_UT.di_AStens_2 ));
    InMux I__3939 (
            .O(N__17544),
            .I(N__17539));
    InMux I__3938 (
            .O(N__17543),
            .I(N__17536));
    CascadeMux I__3937 (
            .O(N__17542),
            .I(N__17532));
    LocalMux I__3936 (
            .O(N__17539),
            .I(N__17529));
    LocalMux I__3935 (
            .O(N__17536),
            .I(N__17526));
    InMux I__3934 (
            .O(N__17535),
            .I(N__17523));
    InMux I__3933 (
            .O(N__17532),
            .I(N__17520));
    Span4Mux_h I__3932 (
            .O(N__17529),
            .I(N__17517));
    Span4Mux_h I__3931 (
            .O(N__17526),
            .I(N__17512));
    LocalMux I__3930 (
            .O(N__17523),
            .I(N__17512));
    LocalMux I__3929 (
            .O(N__17520),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv4 I__3928 (
            .O(N__17517),
            .I(\Lab_UT.di_AStens_3 ));
    Odrv4 I__3927 (
            .O(N__17512),
            .I(\Lab_UT.di_AStens_3 ));
    InMux I__3926 (
            .O(N__17505),
            .I(N__17500));
    InMux I__3925 (
            .O(N__17504),
            .I(N__17497));
    CascadeMux I__3924 (
            .O(N__17503),
            .I(N__17494));
    LocalMux I__3923 (
            .O(N__17500),
            .I(N__17490));
    LocalMux I__3922 (
            .O(N__17497),
            .I(N__17487));
    InMux I__3921 (
            .O(N__17494),
            .I(N__17484));
    InMux I__3920 (
            .O(N__17493),
            .I(N__17481));
    Span4Mux_h I__3919 (
            .O(N__17490),
            .I(N__17476));
    Span4Mux_v I__3918 (
            .O(N__17487),
            .I(N__17476));
    LocalMux I__3917 (
            .O(N__17484),
            .I(N__17473));
    LocalMux I__3916 (
            .O(N__17481),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__3915 (
            .O(N__17476),
            .I(\Lab_UT.di_AMones_0 ));
    Odrv4 I__3914 (
            .O(N__17473),
            .I(\Lab_UT.di_AMones_0 ));
    InMux I__3913 (
            .O(N__17466),
            .I(N__17459));
    InMux I__3912 (
            .O(N__17465),
            .I(N__17459));
    CascadeMux I__3911 (
            .O(N__17464),
            .I(N__17456));
    LocalMux I__3910 (
            .O(N__17459),
            .I(N__17453));
    InMux I__3909 (
            .O(N__17456),
            .I(N__17449));
    Span4Mux_v I__3908 (
            .O(N__17453),
            .I(N__17446));
    InMux I__3907 (
            .O(N__17452),
            .I(N__17443));
    LocalMux I__3906 (
            .O(N__17449),
            .I(\Lab_UT.di_AMones_1 ));
    Odrv4 I__3905 (
            .O(N__17446),
            .I(\Lab_UT.di_AMones_1 ));
    LocalMux I__3904 (
            .O(N__17443),
            .I(\Lab_UT.di_AMones_1 ));
    InMux I__3903 (
            .O(N__17436),
            .I(N__17432));
    InMux I__3902 (
            .O(N__17435),
            .I(N__17429));
    LocalMux I__3901 (
            .O(N__17432),
            .I(N__17425));
    LocalMux I__3900 (
            .O(N__17429),
            .I(N__17422));
    InMux I__3899 (
            .O(N__17428),
            .I(N__17418));
    Span4Mux_h I__3898 (
            .O(N__17425),
            .I(N__17413));
    Span4Mux_h I__3897 (
            .O(N__17422),
            .I(N__17413));
    InMux I__3896 (
            .O(N__17421),
            .I(N__17410));
    LocalMux I__3895 (
            .O(N__17418),
            .I(\Lab_UT.di_AMones_2 ));
    Odrv4 I__3894 (
            .O(N__17413),
            .I(\Lab_UT.di_AMones_2 ));
    LocalMux I__3893 (
            .O(N__17410),
            .I(\Lab_UT.di_AMones_2 ));
    CascadeMux I__3892 (
            .O(N__17403),
            .I(N__17396));
    CascadeMux I__3891 (
            .O(N__17402),
            .I(N__17392));
    CascadeMux I__3890 (
            .O(N__17401),
            .I(N__17388));
    CascadeMux I__3889 (
            .O(N__17400),
            .I(N__17384));
    InMux I__3888 (
            .O(N__17399),
            .I(N__17367));
    InMux I__3887 (
            .O(N__17396),
            .I(N__17367));
    InMux I__3886 (
            .O(N__17395),
            .I(N__17367));
    InMux I__3885 (
            .O(N__17392),
            .I(N__17367));
    InMux I__3884 (
            .O(N__17391),
            .I(N__17367));
    InMux I__3883 (
            .O(N__17388),
            .I(N__17367));
    InMux I__3882 (
            .O(N__17387),
            .I(N__17367));
    InMux I__3881 (
            .O(N__17384),
            .I(N__17367));
    LocalMux I__3880 (
            .O(N__17367),
            .I(N__17364));
    Span4Mux_h I__3879 (
            .O(N__17364),
            .I(N__17361));
    Odrv4 I__3878 (
            .O(N__17361),
            .I(\Lab_UT.N_13_0 ));
    InMux I__3877 (
            .O(N__17358),
            .I(N__17354));
    InMux I__3876 (
            .O(N__17357),
            .I(N__17350));
    LocalMux I__3875 (
            .O(N__17354),
            .I(N__17347));
    CascadeMux I__3874 (
            .O(N__17353),
            .I(N__17344));
    LocalMux I__3873 (
            .O(N__17350),
            .I(N__17341));
    Span4Mux_s0_v I__3872 (
            .O(N__17347),
            .I(N__17338));
    InMux I__3871 (
            .O(N__17344),
            .I(N__17334));
    Span4Mux_v I__3870 (
            .O(N__17341),
            .I(N__17329));
    Span4Mux_v I__3869 (
            .O(N__17338),
            .I(N__17329));
    InMux I__3868 (
            .O(N__17337),
            .I(N__17326));
    LocalMux I__3867 (
            .O(N__17334),
            .I(\Lab_UT.di_AMones_3 ));
    Odrv4 I__3866 (
            .O(N__17329),
            .I(\Lab_UT.di_AMones_3 ));
    LocalMux I__3865 (
            .O(N__17326),
            .I(\Lab_UT.di_AMones_3 ));
    InMux I__3864 (
            .O(N__17319),
            .I(N__17315));
    InMux I__3863 (
            .O(N__17318),
            .I(N__17312));
    LocalMux I__3862 (
            .O(N__17315),
            .I(N__17309));
    LocalMux I__3861 (
            .O(N__17312),
            .I(N__17303));
    Span12Mux_s5_v I__3860 (
            .O(N__17309),
            .I(N__17303));
    InMux I__3859 (
            .O(N__17308),
            .I(N__17300));
    Odrv12 I__3858 (
            .O(N__17303),
            .I(\Lab_UT.di_ASones_1 ));
    LocalMux I__3857 (
            .O(N__17300),
            .I(\Lab_UT.di_ASones_1 ));
    InMux I__3856 (
            .O(N__17295),
            .I(N__17291));
    InMux I__3855 (
            .O(N__17294),
            .I(N__17288));
    LocalMux I__3854 (
            .O(N__17291),
            .I(N__17285));
    LocalMux I__3853 (
            .O(N__17288),
            .I(N__17279));
    Span4Mux_v I__3852 (
            .O(N__17285),
            .I(N__17279));
    InMux I__3851 (
            .O(N__17284),
            .I(N__17276));
    Span4Mux_h I__3850 (
            .O(N__17279),
            .I(N__17273));
    LocalMux I__3849 (
            .O(N__17276),
            .I(N__17270));
    Odrv4 I__3848 (
            .O(N__17273),
            .I(\Lab_UT.di_ASones_2 ));
    Odrv4 I__3847 (
            .O(N__17270),
            .I(\Lab_UT.di_ASones_2 ));
    InMux I__3846 (
            .O(N__17265),
            .I(N__17260));
    InMux I__3845 (
            .O(N__17264),
            .I(N__17257));
    CascadeMux I__3844 (
            .O(N__17263),
            .I(N__17254));
    LocalMux I__3843 (
            .O(N__17260),
            .I(N__17251));
    LocalMux I__3842 (
            .O(N__17257),
            .I(N__17248));
    InMux I__3841 (
            .O(N__17254),
            .I(N__17245));
    Span4Mux_h I__3840 (
            .O(N__17251),
            .I(N__17242));
    Span4Mux_h I__3839 (
            .O(N__17248),
            .I(N__17237));
    LocalMux I__3838 (
            .O(N__17245),
            .I(N__17237));
    Odrv4 I__3837 (
            .O(N__17242),
            .I(\Lab_UT.di_ASones_3 ));
    Odrv4 I__3836 (
            .O(N__17237),
            .I(\Lab_UT.di_ASones_3 ));
    InMux I__3835 (
            .O(N__17232),
            .I(N__17228));
    InMux I__3834 (
            .O(N__17231),
            .I(N__17225));
    LocalMux I__3833 (
            .O(N__17228),
            .I(N__17220));
    LocalMux I__3832 (
            .O(N__17225),
            .I(N__17220));
    Odrv4 I__3831 (
            .O(N__17220),
            .I(\Lab_UT.didp.ceZ0Z_2 ));
    InMux I__3830 (
            .O(N__17217),
            .I(N__17214));
    LocalMux I__3829 (
            .O(N__17214),
            .I(N__17211));
    Odrv4 I__3828 (
            .O(N__17211),
            .I(\Lab_UT.didp.countrce3.q_5_0 ));
    InMux I__3827 (
            .O(N__17208),
            .I(N__17198));
    InMux I__3826 (
            .O(N__17207),
            .I(N__17198));
    InMux I__3825 (
            .O(N__17206),
            .I(N__17192));
    InMux I__3824 (
            .O(N__17205),
            .I(N__17192));
    InMux I__3823 (
            .O(N__17204),
            .I(N__17187));
    InMux I__3822 (
            .O(N__17203),
            .I(N__17187));
    LocalMux I__3821 (
            .O(N__17198),
            .I(N__17184));
    InMux I__3820 (
            .O(N__17197),
            .I(N__17181));
    LocalMux I__3819 (
            .O(N__17192),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    LocalMux I__3818 (
            .O(N__17187),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    Odrv4 I__3817 (
            .O(N__17184),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    LocalMux I__3816 (
            .O(N__17181),
            .I(\Lab_UT.didp.di_Mtens_0 ));
    InMux I__3815 (
            .O(N__17172),
            .I(N__17168));
    InMux I__3814 (
            .O(N__17171),
            .I(N__17165));
    LocalMux I__3813 (
            .O(N__17168),
            .I(N__17162));
    LocalMux I__3812 (
            .O(N__17165),
            .I(N__17159));
    Span4Mux_h I__3811 (
            .O(N__17162),
            .I(N__17155));
    Span4Mux_s2_v I__3810 (
            .O(N__17159),
            .I(N__17152));
    InMux I__3809 (
            .O(N__17158),
            .I(N__17149));
    Odrv4 I__3808 (
            .O(N__17155),
            .I(\Lab_UT.di_AMtens_0 ));
    Odrv4 I__3807 (
            .O(N__17152),
            .I(\Lab_UT.di_AMtens_0 ));
    LocalMux I__3806 (
            .O(N__17149),
            .I(\Lab_UT.di_AMtens_0 ));
    InMux I__3805 (
            .O(N__17142),
            .I(N__17139));
    LocalMux I__3804 (
            .O(N__17139),
            .I(N__17136));
    Span4Mux_h I__3803 (
            .O(N__17136),
            .I(N__17133));
    Odrv4 I__3802 (
            .O(N__17133),
            .I(\Lab_UT.didp.regrce4.did_alarmMatch_6 ));
    CascadeMux I__3801 (
            .O(N__17130),
            .I(N__17124));
    InMux I__3800 (
            .O(N__17129),
            .I(N__17115));
    InMux I__3799 (
            .O(N__17128),
            .I(N__17115));
    InMux I__3798 (
            .O(N__17127),
            .I(N__17115));
    InMux I__3797 (
            .O(N__17124),
            .I(N__17115));
    LocalMux I__3796 (
            .O(N__17115),
            .I(N__17112));
    Span4Mux_v I__3795 (
            .O(N__17112),
            .I(N__17109));
    Odrv4 I__3794 (
            .O(N__17109),
            .I(\Lab_UT.didp.resetZ0Z_2 ));
    CascadeMux I__3793 (
            .O(N__17106),
            .I(N__17103));
    InMux I__3792 (
            .O(N__17103),
            .I(N__17100));
    LocalMux I__3791 (
            .O(N__17100),
            .I(\Lab_UT.didp.countrce3.q_5_3 ));
    InMux I__3790 (
            .O(N__17097),
            .I(N__17091));
    InMux I__3789 (
            .O(N__17096),
            .I(N__17091));
    LocalMux I__3788 (
            .O(N__17091),
            .I(\Lab_UT.didp.un1_dicLdMones_0 ));
    InMux I__3787 (
            .O(N__17088),
            .I(N__17084));
    InMux I__3786 (
            .O(N__17087),
            .I(N__17080));
    LocalMux I__3785 (
            .O(N__17084),
            .I(N__17077));
    InMux I__3784 (
            .O(N__17083),
            .I(N__17072));
    LocalMux I__3783 (
            .O(N__17080),
            .I(N__17069));
    Span4Mux_s3_v I__3782 (
            .O(N__17077),
            .I(N__17066));
    InMux I__3781 (
            .O(N__17076),
            .I(N__17061));
    InMux I__3780 (
            .O(N__17075),
            .I(N__17061));
    LocalMux I__3779 (
            .O(N__17072),
            .I(\Lab_UT.didp.di_Mones_3 ));
    Odrv4 I__3778 (
            .O(N__17069),
            .I(\Lab_UT.didp.di_Mones_3 ));
    Odrv4 I__3777 (
            .O(N__17066),
            .I(\Lab_UT.didp.di_Mones_3 ));
    LocalMux I__3776 (
            .O(N__17061),
            .I(\Lab_UT.didp.di_Mones_3 ));
    InMux I__3775 (
            .O(N__17052),
            .I(N__17046));
    InMux I__3774 (
            .O(N__17051),
            .I(N__17043));
    InMux I__3773 (
            .O(N__17050),
            .I(N__17040));
    InMux I__3772 (
            .O(N__17049),
            .I(N__17036));
    LocalMux I__3771 (
            .O(N__17046),
            .I(N__17029));
    LocalMux I__3770 (
            .O(N__17043),
            .I(N__17029));
    LocalMux I__3769 (
            .O(N__17040),
            .I(N__17029));
    InMux I__3768 (
            .O(N__17039),
            .I(N__17024));
    LocalMux I__3767 (
            .O(N__17036),
            .I(N__17021));
    Span4Mux_s3_v I__3766 (
            .O(N__17029),
            .I(N__17018));
    InMux I__3765 (
            .O(N__17028),
            .I(N__17013));
    InMux I__3764 (
            .O(N__17027),
            .I(N__17013));
    LocalMux I__3763 (
            .O(N__17024),
            .I(\Lab_UT.didp.di_Mones_0 ));
    Odrv4 I__3762 (
            .O(N__17021),
            .I(\Lab_UT.didp.di_Mones_0 ));
    Odrv4 I__3761 (
            .O(N__17018),
            .I(\Lab_UT.didp.di_Mones_0 ));
    LocalMux I__3760 (
            .O(N__17013),
            .I(\Lab_UT.didp.di_Mones_0 ));
    InMux I__3759 (
            .O(N__17004),
            .I(N__16997));
    InMux I__3758 (
            .O(N__17003),
            .I(N__16997));
    InMux I__3757 (
            .O(N__17002),
            .I(N__16993));
    LocalMux I__3756 (
            .O(N__16997),
            .I(N__16987));
    CascadeMux I__3755 (
            .O(N__16996),
            .I(N__16984));
    LocalMux I__3754 (
            .O(N__16993),
            .I(N__16981));
    InMux I__3753 (
            .O(N__16992),
            .I(N__16978));
    InMux I__3752 (
            .O(N__16991),
            .I(N__16973));
    InMux I__3751 (
            .O(N__16990),
            .I(N__16973));
    Span4Mux_h I__3750 (
            .O(N__16987),
            .I(N__16970));
    InMux I__3749 (
            .O(N__16984),
            .I(N__16967));
    Odrv4 I__3748 (
            .O(N__16981),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3747 (
            .O(N__16978),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3746 (
            .O(N__16973),
            .I(\Lab_UT.didp.di_Mones_1 ));
    Odrv4 I__3745 (
            .O(N__16970),
            .I(\Lab_UT.didp.di_Mones_1 ));
    LocalMux I__3744 (
            .O(N__16967),
            .I(\Lab_UT.didp.di_Mones_1 ));
    InMux I__3743 (
            .O(N__16956),
            .I(N__16946));
    InMux I__3742 (
            .O(N__16955),
            .I(N__16946));
    InMux I__3741 (
            .O(N__16954),
            .I(N__16946));
    CascadeMux I__3740 (
            .O(N__16953),
            .I(N__16943));
    LocalMux I__3739 (
            .O(N__16946),
            .I(N__16938));
    InMux I__3738 (
            .O(N__16943),
            .I(N__16935));
    InMux I__3737 (
            .O(N__16942),
            .I(N__16932));
    InMux I__3736 (
            .O(N__16941),
            .I(N__16929));
    Span4Mux_v I__3735 (
            .O(N__16938),
            .I(N__16926));
    LocalMux I__3734 (
            .O(N__16935),
            .I(N__16923));
    LocalMux I__3733 (
            .O(N__16932),
            .I(N__16920));
    LocalMux I__3732 (
            .O(N__16929),
            .I(N__16917));
    Odrv4 I__3731 (
            .O(N__16926),
            .I(\Lab_UT.LdMones ));
    Odrv12 I__3730 (
            .O(N__16923),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3729 (
            .O(N__16920),
            .I(\Lab_UT.LdMones ));
    Odrv4 I__3728 (
            .O(N__16917),
            .I(\Lab_UT.LdMones ));
    CascadeMux I__3727 (
            .O(N__16908),
            .I(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ));
    CascadeMux I__3726 (
            .O(N__16905),
            .I(N__16901));
    InMux I__3725 (
            .O(N__16904),
            .I(N__16895));
    InMux I__3724 (
            .O(N__16901),
            .I(N__16892));
    InMux I__3723 (
            .O(N__16900),
            .I(N__16889));
    InMux I__3722 (
            .O(N__16899),
            .I(N__16886));
    InMux I__3721 (
            .O(N__16898),
            .I(N__16883));
    LocalMux I__3720 (
            .O(N__16895),
            .I(N__16880));
    LocalMux I__3719 (
            .O(N__16892),
            .I(N__16876));
    LocalMux I__3718 (
            .O(N__16889),
            .I(N__16867));
    LocalMux I__3717 (
            .O(N__16886),
            .I(N__16867));
    LocalMux I__3716 (
            .O(N__16883),
            .I(N__16867));
    Span4Mux_s3_v I__3715 (
            .O(N__16880),
            .I(N__16867));
    InMux I__3714 (
            .O(N__16879),
            .I(N__16864));
    Odrv4 I__3713 (
            .O(N__16876),
            .I(\Lab_UT.didp.di_Mones_2 ));
    Odrv4 I__3712 (
            .O(N__16867),
            .I(\Lab_UT.didp.di_Mones_2 ));
    LocalMux I__3711 (
            .O(N__16864),
            .I(\Lab_UT.didp.di_Mones_2 ));
    CascadeMux I__3710 (
            .O(N__16857),
            .I(N__16854));
    InMux I__3709 (
            .O(N__16854),
            .I(N__16851));
    LocalMux I__3708 (
            .O(N__16851),
            .I(\Lab_UT.didp.countrce3.q_5_2 ));
    CascadeMux I__3707 (
            .O(N__16848),
            .I(N__16845));
    InMux I__3706 (
            .O(N__16845),
            .I(N__16835));
    InMux I__3705 (
            .O(N__16844),
            .I(N__16835));
    InMux I__3704 (
            .O(N__16843),
            .I(N__16835));
    InMux I__3703 (
            .O(N__16842),
            .I(N__16832));
    LocalMux I__3702 (
            .O(N__16835),
            .I(N__16829));
    LocalMux I__3701 (
            .O(N__16832),
            .I(\Lab_UT.di_AStens_0 ));
    Odrv12 I__3700 (
            .O(N__16829),
            .I(\Lab_UT.di_AStens_0 ));
    InMux I__3699 (
            .O(N__16824),
            .I(N__16819));
    InMux I__3698 (
            .O(N__16823),
            .I(N__16816));
    CascadeMux I__3697 (
            .O(N__16822),
            .I(N__16812));
    LocalMux I__3696 (
            .O(N__16819),
            .I(N__16809));
    LocalMux I__3695 (
            .O(N__16816),
            .I(N__16806));
    CascadeMux I__3694 (
            .O(N__16815),
            .I(N__16803));
    InMux I__3693 (
            .O(N__16812),
            .I(N__16800));
    Span4Mux_v I__3692 (
            .O(N__16809),
            .I(N__16795));
    Span4Mux_v I__3691 (
            .O(N__16806),
            .I(N__16795));
    InMux I__3690 (
            .O(N__16803),
            .I(N__16792));
    LocalMux I__3689 (
            .O(N__16800),
            .I(\Lab_UT.di_AStens_1 ));
    Odrv4 I__3688 (
            .O(N__16795),
            .I(\Lab_UT.di_AStens_1 ));
    LocalMux I__3687 (
            .O(N__16792),
            .I(\Lab_UT.di_AStens_1 ));
    CascadeMux I__3686 (
            .O(N__16785),
            .I(N__16782));
    InMux I__3685 (
            .O(N__16782),
            .I(N__16774));
    InMux I__3684 (
            .O(N__16781),
            .I(N__16769));
    InMux I__3683 (
            .O(N__16780),
            .I(N__16769));
    InMux I__3682 (
            .O(N__16779),
            .I(N__16766));
    InMux I__3681 (
            .O(N__16778),
            .I(N__16761));
    InMux I__3680 (
            .O(N__16777),
            .I(N__16761));
    LocalMux I__3679 (
            .O(N__16774),
            .I(bu_rx_data_fast_1));
    LocalMux I__3678 (
            .O(N__16769),
            .I(bu_rx_data_fast_1));
    LocalMux I__3677 (
            .O(N__16766),
            .I(bu_rx_data_fast_1));
    LocalMux I__3676 (
            .O(N__16761),
            .I(bu_rx_data_fast_1));
    CascadeMux I__3675 (
            .O(N__16752),
            .I(N__16747));
    CascadeMux I__3674 (
            .O(N__16751),
            .I(N__16742));
    InMux I__3673 (
            .O(N__16750),
            .I(N__16739));
    InMux I__3672 (
            .O(N__16747),
            .I(N__16736));
    CascadeMux I__3671 (
            .O(N__16746),
            .I(N__16733));
    InMux I__3670 (
            .O(N__16745),
            .I(N__16726));
    InMux I__3669 (
            .O(N__16742),
            .I(N__16726));
    LocalMux I__3668 (
            .O(N__16739),
            .I(N__16721));
    LocalMux I__3667 (
            .O(N__16736),
            .I(N__16721));
    InMux I__3666 (
            .O(N__16733),
            .I(N__16717));
    InMux I__3665 (
            .O(N__16732),
            .I(N__16714));
    CascadeMux I__3664 (
            .O(N__16731),
            .I(N__16711));
    LocalMux I__3663 (
            .O(N__16726),
            .I(N__16707));
    Span4Mux_h I__3662 (
            .O(N__16721),
            .I(N__16704));
    InMux I__3661 (
            .O(N__16720),
            .I(N__16701));
    LocalMux I__3660 (
            .O(N__16717),
            .I(N__16696));
    LocalMux I__3659 (
            .O(N__16714),
            .I(N__16696));
    InMux I__3658 (
            .O(N__16711),
            .I(N__16691));
    InMux I__3657 (
            .O(N__16710),
            .I(N__16691));
    Odrv4 I__3656 (
            .O(N__16707),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__3655 (
            .O(N__16704),
            .I(bu_rx_data_3_rep1));
    LocalMux I__3654 (
            .O(N__16701),
            .I(bu_rx_data_3_rep1));
    Odrv4 I__3653 (
            .O(N__16696),
            .I(bu_rx_data_3_rep1));
    LocalMux I__3652 (
            .O(N__16691),
            .I(bu_rx_data_3_rep1));
    InMux I__3651 (
            .O(N__16680),
            .I(N__16677));
    LocalMux I__3650 (
            .O(N__16677),
            .I(N__16674));
    Odrv4 I__3649 (
            .O(N__16674),
            .I(\Lab_UT.dictrl.g1_1Z0Z_1 ));
    InMux I__3648 (
            .O(N__16671),
            .I(N__16668));
    LocalMux I__3647 (
            .O(N__16668),
            .I(N__16665));
    Odrv4 I__3646 (
            .O(N__16665),
            .I(\Lab_UT.dictrl.g2_1_0 ));
    InMux I__3645 (
            .O(N__16662),
            .I(N__16659));
    LocalMux I__3644 (
            .O(N__16659),
            .I(N__16656));
    Odrv4 I__3643 (
            .O(N__16656),
            .I(\Lab_UT.dictrl.g2 ));
    InMux I__3642 (
            .O(N__16653),
            .I(N__16646));
    InMux I__3641 (
            .O(N__16652),
            .I(N__16646));
    InMux I__3640 (
            .O(N__16651),
            .I(N__16643));
    LocalMux I__3639 (
            .O(N__16646),
            .I(\Lab_UT.didp.countrce3.ce_12_2_3 ));
    LocalMux I__3638 (
            .O(N__16643),
            .I(\Lab_UT.didp.countrce3.ce_12_2_3 ));
    InMux I__3637 (
            .O(N__16638),
            .I(N__16635));
    LocalMux I__3636 (
            .O(N__16635),
            .I(N__16631));
    InMux I__3635 (
            .O(N__16634),
            .I(N__16628));
    Span4Mux_h I__3634 (
            .O(N__16631),
            .I(N__16624));
    LocalMux I__3633 (
            .O(N__16628),
            .I(N__16621));
    CascadeMux I__3632 (
            .O(N__16627),
            .I(N__16618));
    Span4Mux_v I__3631 (
            .O(N__16624),
            .I(N__16613));
    Span4Mux_s2_v I__3630 (
            .O(N__16621),
            .I(N__16613));
    InMux I__3629 (
            .O(N__16618),
            .I(N__16610));
    Odrv4 I__3628 (
            .O(N__16613),
            .I(\Lab_UT.di_AMtens_3 ));
    LocalMux I__3627 (
            .O(N__16610),
            .I(\Lab_UT.di_AMtens_3 ));
    CEMux I__3626 (
            .O(N__16605),
            .I(N__16601));
    CEMux I__3625 (
            .O(N__16604),
            .I(N__16598));
    LocalMux I__3624 (
            .O(N__16601),
            .I(N__16595));
    LocalMux I__3623 (
            .O(N__16598),
            .I(N__16592));
    Span4Mux_h I__3622 (
            .O(N__16595),
            .I(N__16589));
    Span4Mux_h I__3621 (
            .O(N__16592),
            .I(N__16586));
    Span4Mux_v I__3620 (
            .O(N__16589),
            .I(N__16583));
    Span4Mux_h I__3619 (
            .O(N__16586),
            .I(N__16580));
    Odrv4 I__3618 (
            .O(N__16583),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    Odrv4 I__3617 (
            .O(N__16580),
            .I(\Lab_UT.didp.regrce4.LdAMtens_0 ));
    CascadeMux I__3616 (
            .O(N__16575),
            .I(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ));
    InMux I__3615 (
            .O(N__16572),
            .I(N__16569));
    LocalMux I__3614 (
            .O(N__16569),
            .I(N__16566));
    Span4Mux_h I__3613 (
            .O(N__16566),
            .I(N__16563));
    Odrv4 I__3612 (
            .O(N__16563),
            .I(\Lab_UT.didp.countrce3.q_5_1 ));
    InMux I__3611 (
            .O(N__16560),
            .I(N__16557));
    LocalMux I__3610 (
            .O(N__16557),
            .I(\Lab_UT.dictrl.g0_2Z0Z_4 ));
    CascadeMux I__3609 (
            .O(N__16554),
            .I(\Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ));
    InMux I__3608 (
            .O(N__16551),
            .I(N__16548));
    LocalMux I__3607 (
            .O(N__16548),
            .I(\Lab_UT.dictrl.N_77_1_0 ));
    CascadeMux I__3606 (
            .O(N__16545),
            .I(\Lab_UT.dictrl.N_77_1_0_cascade_ ));
    InMux I__3605 (
            .O(N__16542),
            .I(N__16539));
    LocalMux I__3604 (
            .O(N__16539),
            .I(\Lab_UT.dictrl.N_2353_0_0 ));
    CascadeMux I__3603 (
            .O(N__16536),
            .I(N__16528));
    CascadeMux I__3602 (
            .O(N__16535),
            .I(N__16525));
    InMux I__3601 (
            .O(N__16534),
            .I(N__16520));
    InMux I__3600 (
            .O(N__16533),
            .I(N__16520));
    InMux I__3599 (
            .O(N__16532),
            .I(N__16510));
    InMux I__3598 (
            .O(N__16531),
            .I(N__16510));
    InMux I__3597 (
            .O(N__16528),
            .I(N__16510));
    InMux I__3596 (
            .O(N__16525),
            .I(N__16510));
    LocalMux I__3595 (
            .O(N__16520),
            .I(N__16507));
    CascadeMux I__3594 (
            .O(N__16519),
            .I(N__16504));
    LocalMux I__3593 (
            .O(N__16510),
            .I(N__16501));
    Span4Mux_h I__3592 (
            .O(N__16507),
            .I(N__16498));
    InMux I__3591 (
            .O(N__16504),
            .I(N__16495));
    Span4Mux_h I__3590 (
            .O(N__16501),
            .I(N__16492));
    Odrv4 I__3589 (
            .O(N__16498),
            .I(buart__rx_shifter_fast_6));
    LocalMux I__3588 (
            .O(N__16495),
            .I(buart__rx_shifter_fast_6));
    Odrv4 I__3587 (
            .O(N__16492),
            .I(buart__rx_shifter_fast_6));
    CascadeMux I__3586 (
            .O(N__16485),
            .I(N__16481));
    InMux I__3585 (
            .O(N__16484),
            .I(N__16470));
    InMux I__3584 (
            .O(N__16481),
            .I(N__16470));
    InMux I__3583 (
            .O(N__16480),
            .I(N__16470));
    InMux I__3582 (
            .O(N__16479),
            .I(N__16470));
    LocalMux I__3581 (
            .O(N__16470),
            .I(N__16466));
    InMux I__3580 (
            .O(N__16469),
            .I(N__16463));
    Span4Mux_h I__3579 (
            .O(N__16466),
            .I(N__16460));
    LocalMux I__3578 (
            .O(N__16463),
            .I(bu_rx_data_fast_7));
    Odrv4 I__3577 (
            .O(N__16460),
            .I(bu_rx_data_fast_7));
    InMux I__3576 (
            .O(N__16455),
            .I(N__16452));
    LocalMux I__3575 (
            .O(N__16452),
            .I(\Lab_UT.dictrl.state_fast_3 ));
    InMux I__3574 (
            .O(N__16449),
            .I(N__16443));
    InMux I__3573 (
            .O(N__16448),
            .I(N__16443));
    LocalMux I__3572 (
            .O(N__16443),
            .I(N__16440));
    Odrv4 I__3571 (
            .O(N__16440),
            .I(\Lab_UT.dictrl.g1_6 ));
    CascadeMux I__3570 (
            .O(N__16437),
            .I(\Lab_UT.dictrl.m47_xZ0Z0_cascade_ ));
    InMux I__3569 (
            .O(N__16434),
            .I(N__16429));
    InMux I__3568 (
            .O(N__16433),
            .I(N__16424));
    InMux I__3567 (
            .O(N__16432),
            .I(N__16424));
    LocalMux I__3566 (
            .O(N__16429),
            .I(N__16417));
    LocalMux I__3565 (
            .O(N__16424),
            .I(N__16417));
    InMux I__3564 (
            .O(N__16423),
            .I(N__16412));
    InMux I__3563 (
            .O(N__16422),
            .I(N__16412));
    Odrv4 I__3562 (
            .O(N__16417),
            .I(bu_rx_data_fast_4));
    LocalMux I__3561 (
            .O(N__16412),
            .I(bu_rx_data_fast_4));
    InMux I__3560 (
            .O(N__16407),
            .I(N__16401));
    InMux I__3559 (
            .O(N__16406),
            .I(N__16401));
    LocalMux I__3558 (
            .O(N__16401),
            .I(N__16398));
    Odrv4 I__3557 (
            .O(N__16398),
            .I(\Lab_UT.dictrl.m30Z0Z_1 ));
    InMux I__3556 (
            .O(N__16395),
            .I(N__16392));
    LocalMux I__3555 (
            .O(N__16392),
            .I(\Lab_UT.dictrl.N_81_0 ));
    CascadeMux I__3554 (
            .O(N__16389),
            .I(\Lab_UT.dictrl.N_16_mux_0_cascade_ ));
    InMux I__3553 (
            .O(N__16386),
            .I(N__16383));
    LocalMux I__3552 (
            .O(N__16383),
            .I(\Lab_UT.dictrl.N_113_0_0 ));
    InMux I__3551 (
            .O(N__16380),
            .I(N__16373));
    InMux I__3550 (
            .O(N__16379),
            .I(N__16368));
    InMux I__3549 (
            .O(N__16378),
            .I(N__16368));
    InMux I__3548 (
            .O(N__16377),
            .I(N__16363));
    CascadeMux I__3547 (
            .O(N__16376),
            .I(N__16360));
    LocalMux I__3546 (
            .O(N__16373),
            .I(N__16356));
    LocalMux I__3545 (
            .O(N__16368),
            .I(N__16353));
    InMux I__3544 (
            .O(N__16367),
            .I(N__16350));
    InMux I__3543 (
            .O(N__16366),
            .I(N__16347));
    LocalMux I__3542 (
            .O(N__16363),
            .I(N__16344));
    InMux I__3541 (
            .O(N__16360),
            .I(N__16339));
    InMux I__3540 (
            .O(N__16359),
            .I(N__16339));
    Span4Mux_v I__3539 (
            .O(N__16356),
            .I(N__16332));
    Span4Mux_h I__3538 (
            .O(N__16353),
            .I(N__16332));
    LocalMux I__3537 (
            .O(N__16350),
            .I(N__16332));
    LocalMux I__3536 (
            .O(N__16347),
            .I(N__16325));
    Span4Mux_v I__3535 (
            .O(N__16344),
            .I(N__16325));
    LocalMux I__3534 (
            .O(N__16339),
            .I(N__16325));
    Span4Mux_v I__3533 (
            .O(N__16332),
            .I(N__16322));
    Odrv4 I__3532 (
            .O(N__16325),
            .I(\Lab_UT.dictrl.state_2_rep1 ));
    Odrv4 I__3531 (
            .O(N__16322),
            .I(\Lab_UT.dictrl.state_2_rep1 ));
    CascadeMux I__3530 (
            .O(N__16317),
            .I(\Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_ ));
    InMux I__3529 (
            .O(N__16314),
            .I(N__16311));
    LocalMux I__3528 (
            .O(N__16311),
            .I(\Lab_UT.dictrl.N_5_0 ));
    CascadeMux I__3527 (
            .O(N__16308),
            .I(\Lab_UT.dictrl.g2_2_cascade_ ));
    InMux I__3526 (
            .O(N__16305),
            .I(N__16302));
    LocalMux I__3525 (
            .O(N__16302),
            .I(N__16298));
    InMux I__3524 (
            .O(N__16301),
            .I(N__16295));
    Odrv12 I__3523 (
            .O(N__16298),
            .I(\Lab_UT.dictrl.i9_mux_0 ));
    LocalMux I__3522 (
            .O(N__16295),
            .I(\Lab_UT.dictrl.i9_mux_0 ));
    InMux I__3521 (
            .O(N__16290),
            .I(N__16287));
    LocalMux I__3520 (
            .O(N__16287),
            .I(N__16284));
    Span4Mux_h I__3519 (
            .O(N__16284),
            .I(N__16280));
    InMux I__3518 (
            .O(N__16283),
            .I(N__16277));
    Odrv4 I__3517 (
            .O(N__16280),
            .I(\Lab_UT.dictrl.N_77_0 ));
    LocalMux I__3516 (
            .O(N__16277),
            .I(\Lab_UT.dictrl.N_77_0 ));
    InMux I__3515 (
            .O(N__16272),
            .I(N__16267));
    InMux I__3514 (
            .O(N__16271),
            .I(N__16264));
    InMux I__3513 (
            .O(N__16270),
            .I(N__16261));
    LocalMux I__3512 (
            .O(N__16267),
            .I(N__16253));
    LocalMux I__3511 (
            .O(N__16264),
            .I(N__16253));
    LocalMux I__3510 (
            .O(N__16261),
            .I(N__16250));
    InMux I__3509 (
            .O(N__16260),
            .I(N__16247));
    InMux I__3508 (
            .O(N__16259),
            .I(N__16242));
    InMux I__3507 (
            .O(N__16258),
            .I(N__16242));
    Odrv4 I__3506 (
            .O(N__16253),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    Odrv4 I__3505 (
            .O(N__16250),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    LocalMux I__3504 (
            .O(N__16247),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    LocalMux I__3503 (
            .O(N__16242),
            .I(\Lab_UT.dictrl.state_3_rep1 ));
    InMux I__3502 (
            .O(N__16233),
            .I(N__16230));
    LocalMux I__3501 (
            .O(N__16230),
            .I(\Lab_UT.dictrl.g0_0Z0Z_1 ));
    InMux I__3500 (
            .O(N__16227),
            .I(N__16224));
    LocalMux I__3499 (
            .O(N__16224),
            .I(N__16220));
    InMux I__3498 (
            .O(N__16223),
            .I(N__16217));
    Span12Mux_s6_h I__3497 (
            .O(N__16220),
            .I(N__16214));
    LocalMux I__3496 (
            .O(N__16217),
            .I(N__16211));
    Odrv12 I__3495 (
            .O(N__16214),
            .I(\Lab_UT.dictrl.m30_0Z0Z_0 ));
    Odrv12 I__3494 (
            .O(N__16211),
            .I(\Lab_UT.dictrl.m30_0Z0Z_0 ));
    CascadeMux I__3493 (
            .O(N__16206),
            .I(\Lab_UT.dictrl.m25Z0Z_0_cascade_ ));
    InMux I__3492 (
            .O(N__16203),
            .I(N__16200));
    LocalMux I__3491 (
            .O(N__16200),
            .I(N__16197));
    Span4Mux_h I__3490 (
            .O(N__16197),
            .I(N__16194));
    Odrv4 I__3489 (
            .O(N__16194),
            .I(\Lab_UT.dictrl.m59_ns_1_xZ0Z1 ));
    CascadeMux I__3488 (
            .O(N__16191),
            .I(\Lab_UT.dictrl.N_81_1_cascade_ ));
    InMux I__3487 (
            .O(N__16188),
            .I(N__16185));
    LocalMux I__3486 (
            .O(N__16185),
            .I(\Lab_UT.dictrl.N_113_1 ));
    CascadeMux I__3485 (
            .O(N__16182),
            .I(\Lab_UT.dictrl.N_113_1_cascade_ ));
    InMux I__3484 (
            .O(N__16179),
            .I(N__16173));
    InMux I__3483 (
            .O(N__16178),
            .I(N__16166));
    InMux I__3482 (
            .O(N__16177),
            .I(N__16166));
    InMux I__3481 (
            .O(N__16176),
            .I(N__16166));
    LocalMux I__3480 (
            .O(N__16173),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    LocalMux I__3479 (
            .O(N__16166),
            .I(\Lab_UT.dictrl.next_stateZ0Z_0 ));
    InMux I__3478 (
            .O(N__16161),
            .I(N__16156));
    InMux I__3477 (
            .O(N__16160),
            .I(N__16153));
    InMux I__3476 (
            .O(N__16159),
            .I(N__16150));
    LocalMux I__3475 (
            .O(N__16156),
            .I(N__16145));
    LocalMux I__3474 (
            .O(N__16153),
            .I(N__16145));
    LocalMux I__3473 (
            .O(N__16150),
            .I(N__16142));
    Span4Mux_v I__3472 (
            .O(N__16145),
            .I(N__16139));
    Span4Mux_v I__3471 (
            .O(N__16142),
            .I(N__16136));
    Odrv4 I__3470 (
            .O(N__16139),
            .I(\Lab_UT.dictrl.m59_ns_1 ));
    Odrv4 I__3469 (
            .O(N__16136),
            .I(\Lab_UT.dictrl.m59_ns_1 ));
    InMux I__3468 (
            .O(N__16131),
            .I(N__16128));
    LocalMux I__3467 (
            .O(N__16128),
            .I(N__16125));
    Span4Mux_v I__3466 (
            .O(N__16125),
            .I(N__16122));
    Odrv4 I__3465 (
            .O(N__16122),
            .I(\Lab_UT.dictrl.state_fast_2 ));
    CascadeMux I__3464 (
            .O(N__16119),
            .I(N__16116));
    InMux I__3463 (
            .O(N__16116),
            .I(N__16107));
    InMux I__3462 (
            .O(N__16115),
            .I(N__16107));
    InMux I__3461 (
            .O(N__16114),
            .I(N__16107));
    LocalMux I__3460 (
            .O(N__16107),
            .I(N__16103));
    InMux I__3459 (
            .O(N__16106),
            .I(N__16100));
    Span4Mux_h I__3458 (
            .O(N__16103),
            .I(N__16097));
    LocalMux I__3457 (
            .O(N__16100),
            .I(N__16094));
    Span4Mux_v I__3456 (
            .O(N__16097),
            .I(N__16091));
    Sp12to4 I__3455 (
            .O(N__16094),
            .I(N__16088));
    Odrv4 I__3454 (
            .O(N__16091),
            .I(\Lab_UT.dictrl.g0_17_0 ));
    Odrv12 I__3453 (
            .O(N__16088),
            .I(\Lab_UT.dictrl.g0_17_0 ));
    InMux I__3452 (
            .O(N__16083),
            .I(N__16074));
    InMux I__3451 (
            .O(N__16082),
            .I(N__16074));
    InMux I__3450 (
            .O(N__16081),
            .I(N__16074));
    LocalMux I__3449 (
            .O(N__16074),
            .I(N__16070));
    InMux I__3448 (
            .O(N__16073),
            .I(N__16067));
    Span4Mux_h I__3447 (
            .O(N__16070),
            .I(N__16064));
    LocalMux I__3446 (
            .O(N__16067),
            .I(N__16061));
    Span4Mux_v I__3445 (
            .O(N__16064),
            .I(N__16057));
    Span4Mux_v I__3444 (
            .O(N__16061),
            .I(N__16054));
    InMux I__3443 (
            .O(N__16060),
            .I(N__16051));
    Odrv4 I__3442 (
            .O(N__16057),
            .I(\Lab_UT.dictrl.g0_17_1 ));
    Odrv4 I__3441 (
            .O(N__16054),
            .I(\Lab_UT.dictrl.g0_17_1 ));
    LocalMux I__3440 (
            .O(N__16051),
            .I(\Lab_UT.dictrl.g0_17_1 ));
    InMux I__3439 (
            .O(N__16044),
            .I(N__16040));
    InMux I__3438 (
            .O(N__16043),
            .I(N__16036));
    LocalMux I__3437 (
            .O(N__16040),
            .I(N__16031));
    InMux I__3436 (
            .O(N__16039),
            .I(N__16027));
    LocalMux I__3435 (
            .O(N__16036),
            .I(N__16024));
    InMux I__3434 (
            .O(N__16035),
            .I(N__16021));
    InMux I__3433 (
            .O(N__16034),
            .I(N__16018));
    Span4Mux_h I__3432 (
            .O(N__16031),
            .I(N__16015));
    InMux I__3431 (
            .O(N__16030),
            .I(N__16012));
    LocalMux I__3430 (
            .O(N__16027),
            .I(\Lab_UT.didp.di_Sones_2 ));
    Odrv4 I__3429 (
            .O(N__16024),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__3428 (
            .O(N__16021),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__3427 (
            .O(N__16018),
            .I(\Lab_UT.didp.di_Sones_2 ));
    Odrv4 I__3426 (
            .O(N__16015),
            .I(\Lab_UT.didp.di_Sones_2 ));
    LocalMux I__3425 (
            .O(N__16012),
            .I(\Lab_UT.didp.di_Sones_2 ));
    InMux I__3424 (
            .O(N__15999),
            .I(N__15995));
    InMux I__3423 (
            .O(N__15998),
            .I(N__15990));
    LocalMux I__3422 (
            .O(N__15995),
            .I(N__15987));
    InMux I__3421 (
            .O(N__15994),
            .I(N__15983));
    InMux I__3420 (
            .O(N__15993),
            .I(N__15980));
    LocalMux I__3419 (
            .O(N__15990),
            .I(N__15977));
    Span4Mux_h I__3418 (
            .O(N__15987),
            .I(N__15974));
    InMux I__3417 (
            .O(N__15986),
            .I(N__15971));
    LocalMux I__3416 (
            .O(N__15983),
            .I(\Lab_UT.didp.di_Sones_3 ));
    LocalMux I__3415 (
            .O(N__15980),
            .I(\Lab_UT.didp.di_Sones_3 ));
    Odrv4 I__3414 (
            .O(N__15977),
            .I(\Lab_UT.didp.di_Sones_3 ));
    Odrv4 I__3413 (
            .O(N__15974),
            .I(\Lab_UT.didp.di_Sones_3 ));
    LocalMux I__3412 (
            .O(N__15971),
            .I(\Lab_UT.didp.di_Sones_3 ));
    InMux I__3411 (
            .O(N__15960),
            .I(N__15942));
    InMux I__3410 (
            .O(N__15959),
            .I(N__15942));
    InMux I__3409 (
            .O(N__15958),
            .I(N__15942));
    InMux I__3408 (
            .O(N__15957),
            .I(N__15942));
    InMux I__3407 (
            .O(N__15956),
            .I(N__15942));
    InMux I__3406 (
            .O(N__15955),
            .I(N__15942));
    LocalMux I__3405 (
            .O(N__15942),
            .I(N__15938));
    InMux I__3404 (
            .O(N__15941),
            .I(N__15935));
    Span4Mux_v I__3403 (
            .O(N__15938),
            .I(N__15932));
    LocalMux I__3402 (
            .O(N__15935),
            .I(\Lab_UT.didp.un18_ce ));
    Odrv4 I__3401 (
            .O(N__15932),
            .I(\Lab_UT.didp.un18_ce ));
    InMux I__3400 (
            .O(N__15927),
            .I(N__15924));
    LocalMux I__3399 (
            .O(N__15924),
            .I(N__15921));
    Odrv4 I__3398 (
            .O(N__15921),
            .I(\Lab_UT.LdSones_i_3 ));
    InMux I__3397 (
            .O(N__15918),
            .I(N__15914));
    InMux I__3396 (
            .O(N__15917),
            .I(N__15911));
    LocalMux I__3395 (
            .O(N__15914),
            .I(N__15908));
    LocalMux I__3394 (
            .O(N__15911),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    Odrv4 I__3393 (
            .O(N__15908),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1 ));
    CascadeMux I__3392 (
            .O(N__15903),
            .I(N__15898));
    CascadeMux I__3391 (
            .O(N__15902),
            .I(N__15894));
    InMux I__3390 (
            .O(N__15901),
            .I(N__15887));
    InMux I__3389 (
            .O(N__15898),
            .I(N__15887));
    InMux I__3388 (
            .O(N__15897),
            .I(N__15887));
    InMux I__3387 (
            .O(N__15894),
            .I(N__15884));
    LocalMux I__3386 (
            .O(N__15887),
            .I(N__15881));
    LocalMux I__3385 (
            .O(N__15884),
            .I(N__15878));
    Odrv12 I__3384 (
            .O(N__15881),
            .I(\Lab_UT.LdStens ));
    Odrv4 I__3383 (
            .O(N__15878),
            .I(\Lab_UT.LdStens ));
    CEMux I__3382 (
            .O(N__15873),
            .I(N__15858));
    CEMux I__3381 (
            .O(N__15872),
            .I(N__15858));
    CEMux I__3380 (
            .O(N__15871),
            .I(N__15858));
    CEMux I__3379 (
            .O(N__15870),
            .I(N__15858));
    CEMux I__3378 (
            .O(N__15869),
            .I(N__15858));
    GlobalMux I__3377 (
            .O(N__15858),
            .I(N__15855));
    gio2CtrlBuf I__3376 (
            .O(N__15855),
            .I(bu_rx_data_rdy_0_g));
    InMux I__3375 (
            .O(N__15852),
            .I(N__15849));
    LocalMux I__3374 (
            .O(N__15849),
            .I(\Lab_UT.didp.countrce1.un13_qPone ));
    CascadeMux I__3373 (
            .O(N__15846),
            .I(\Lab_UT.didp.countrce1.q_5_2_cascade_ ));
    InMux I__3372 (
            .O(N__15843),
            .I(N__15839));
    InMux I__3371 (
            .O(N__15842),
            .I(N__15836));
    LocalMux I__3370 (
            .O(N__15839),
            .I(N__15833));
    LocalMux I__3369 (
            .O(N__15836),
            .I(N__15828));
    Span4Mux_v I__3368 (
            .O(N__15833),
            .I(N__15825));
    InMux I__3367 (
            .O(N__15832),
            .I(N__15820));
    InMux I__3366 (
            .O(N__15831),
            .I(N__15820));
    Span4Mux_h I__3365 (
            .O(N__15828),
            .I(N__15817));
    Odrv4 I__3364 (
            .O(N__15825),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    LocalMux I__3363 (
            .O(N__15820),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    Odrv4 I__3362 (
            .O(N__15817),
            .I(\Lab_UT.didp.un1_dicLdSones_0 ));
    InMux I__3361 (
            .O(N__15810),
            .I(N__15807));
    LocalMux I__3360 (
            .O(N__15807),
            .I(N__15803));
    InMux I__3359 (
            .O(N__15806),
            .I(N__15798));
    Span4Mux_v I__3358 (
            .O(N__15803),
            .I(N__15795));
    InMux I__3357 (
            .O(N__15802),
            .I(N__15790));
    InMux I__3356 (
            .O(N__15801),
            .I(N__15790));
    LocalMux I__3355 (
            .O(N__15798),
            .I(N__15787));
    Span4Mux_s1_v I__3354 (
            .O(N__15795),
            .I(N__15784));
    LocalMux I__3353 (
            .O(N__15790),
            .I(N__15779));
    Sp12to4 I__3352 (
            .O(N__15787),
            .I(N__15779));
    Odrv4 I__3351 (
            .O(N__15784),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    Odrv12 I__3350 (
            .O(N__15779),
            .I(\Lab_UT.didp.resetZ0Z_0 ));
    InMux I__3349 (
            .O(N__15774),
            .I(N__15771));
    LocalMux I__3348 (
            .O(N__15771),
            .I(N__15768));
    Odrv4 I__3347 (
            .O(N__15768),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0 ));
    InMux I__3346 (
            .O(N__15765),
            .I(N__15762));
    LocalMux I__3345 (
            .O(N__15762),
            .I(\Lab_UT.un1_idle_5_0_iclkZ0 ));
    CascadeMux I__3344 (
            .O(N__15759),
            .I(N__15756));
    InMux I__3343 (
            .O(N__15756),
            .I(N__15753));
    LocalMux I__3342 (
            .O(N__15753),
            .I(N__15748));
    InMux I__3341 (
            .O(N__15752),
            .I(N__15745));
    InMux I__3340 (
            .O(N__15751),
            .I(N__15741));
    Span4Mux_v I__3339 (
            .O(N__15748),
            .I(N__15736));
    LocalMux I__3338 (
            .O(N__15745),
            .I(N__15736));
    SRMux I__3337 (
            .O(N__15744),
            .I(N__15733));
    LocalMux I__3336 (
            .O(N__15741),
            .I(N__15730));
    Span4Mux_v I__3335 (
            .O(N__15736),
            .I(N__15724));
    LocalMux I__3334 (
            .O(N__15733),
            .I(N__15724));
    Span12Mux_v I__3333 (
            .O(N__15730),
            .I(N__15721));
    IoInMux I__3332 (
            .O(N__15729),
            .I(N__15718));
    Span4Mux_h I__3331 (
            .O(N__15724),
            .I(N__15715));
    Odrv12 I__3330 (
            .O(N__15721),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3329 (
            .O(N__15718),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3328 (
            .O(N__15715),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__3327 (
            .O(N__15708),
            .I(\Lab_UT.un1_armed_2_0_iso_iZ0_cascade_ ));
    InMux I__3326 (
            .O(N__15705),
            .I(N__15701));
    InMux I__3325 (
            .O(N__15704),
            .I(N__15698));
    LocalMux I__3324 (
            .O(N__15701),
            .I(G_192));
    LocalMux I__3323 (
            .O(N__15698),
            .I(G_192));
    CascadeMux I__3322 (
            .O(N__15693),
            .I(\Lab_UT.dictrl.N_113_cascade_ ));
    InMux I__3321 (
            .O(N__15690),
            .I(N__15687));
    LocalMux I__3320 (
            .O(N__15687),
            .I(N__15684));
    Span4Mux_h I__3319 (
            .O(N__15684),
            .I(N__15681));
    Odrv4 I__3318 (
            .O(N__15681),
            .I(\Lab_UT.didp.did_alarmMatch_7 ));
    CascadeMux I__3317 (
            .O(N__15678),
            .I(\Lab_UT.didp.did_alarmMatch_4_cascade_ ));
    InMux I__3316 (
            .O(N__15675),
            .I(N__15672));
    LocalMux I__3315 (
            .O(N__15672),
            .I(\Lab_UT.didp.did_alarmMatch_5 ));
    CascadeMux I__3314 (
            .O(N__15669),
            .I(\Lab_UT.did_alarmMatch_13_cascade_ ));
    CascadeMux I__3313 (
            .O(N__15666),
            .I(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ));
    InMux I__3312 (
            .O(N__15663),
            .I(N__15660));
    LocalMux I__3311 (
            .O(N__15660),
            .I(\Lab_UT.did_alarmMatch_13 ));
    CascadeMux I__3310 (
            .O(N__15657),
            .I(G_183_cascade_));
    InMux I__3309 (
            .O(N__15654),
            .I(N__15648));
    InMux I__3308 (
            .O(N__15653),
            .I(N__15648));
    LocalMux I__3307 (
            .O(N__15648),
            .I(N__15645));
    Odrv4 I__3306 (
            .O(N__15645),
            .I(\Lab_UT.did_alarmMatch_12 ));
    InMux I__3305 (
            .O(N__15642),
            .I(N__15639));
    LocalMux I__3304 (
            .O(N__15639),
            .I(N__15636));
    Odrv4 I__3303 (
            .O(N__15636),
            .I(\Lab_UT.didp.countrce2.un13_qPone ));
    InMux I__3302 (
            .O(N__15633),
            .I(N__15628));
    InMux I__3301 (
            .O(N__15632),
            .I(N__15622));
    InMux I__3300 (
            .O(N__15631),
            .I(N__15622));
    LocalMux I__3299 (
            .O(N__15628),
            .I(N__15619));
    InMux I__3298 (
            .O(N__15627),
            .I(N__15614));
    LocalMux I__3297 (
            .O(N__15622),
            .I(N__15611));
    Span4Mux_h I__3296 (
            .O(N__15619),
            .I(N__15608));
    InMux I__3295 (
            .O(N__15618),
            .I(N__15603));
    InMux I__3294 (
            .O(N__15617),
            .I(N__15603));
    LocalMux I__3293 (
            .O(N__15614),
            .I(\Lab_UT.didp.di_Stens_2 ));
    Odrv4 I__3292 (
            .O(N__15611),
            .I(\Lab_UT.didp.di_Stens_2 ));
    Odrv4 I__3291 (
            .O(N__15608),
            .I(\Lab_UT.didp.di_Stens_2 ));
    LocalMux I__3290 (
            .O(N__15603),
            .I(\Lab_UT.didp.di_Stens_2 ));
    InMux I__3289 (
            .O(N__15594),
            .I(N__15591));
    LocalMux I__3288 (
            .O(N__15591),
            .I(N__15588));
    Odrv4 I__3287 (
            .O(N__15588),
            .I(\Lab_UT.didp.countrce2.q_5_2 ));
    IoInMux I__3286 (
            .O(N__15585),
            .I(N__15579));
    InMux I__3285 (
            .O(N__15584),
            .I(N__15575));
    InMux I__3284 (
            .O(N__15583),
            .I(N__15571));
    InMux I__3283 (
            .O(N__15582),
            .I(N__15568));
    LocalMux I__3282 (
            .O(N__15579),
            .I(N__15565));
    InMux I__3281 (
            .O(N__15578),
            .I(N__15562));
    LocalMux I__3280 (
            .O(N__15575),
            .I(N__15559));
    InMux I__3279 (
            .O(N__15574),
            .I(N__15556));
    LocalMux I__3278 (
            .O(N__15571),
            .I(N__15553));
    LocalMux I__3277 (
            .O(N__15568),
            .I(N__15550));
    Span4Mux_s0_h I__3276 (
            .O(N__15565),
            .I(N__15547));
    LocalMux I__3275 (
            .O(N__15562),
            .I(N__15544));
    Span4Mux_v I__3274 (
            .O(N__15559),
            .I(N__15541));
    LocalMux I__3273 (
            .O(N__15556),
            .I(N__15538));
    Span4Mux_v I__3272 (
            .O(N__15553),
            .I(N__15533));
    Span4Mux_v I__3271 (
            .O(N__15550),
            .I(N__15533));
    Span4Mux_h I__3270 (
            .O(N__15547),
            .I(N__15530));
    Span4Mux_v I__3269 (
            .O(N__15544),
            .I(N__15527));
    Odrv4 I__3268 (
            .O(N__15541),
            .I(rst));
    Odrv12 I__3267 (
            .O(N__15538),
            .I(rst));
    Odrv4 I__3266 (
            .O(N__15533),
            .I(rst));
    Odrv4 I__3265 (
            .O(N__15530),
            .I(rst));
    Odrv4 I__3264 (
            .O(N__15527),
            .I(rst));
    CascadeMux I__3263 (
            .O(N__15516),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ));
    InMux I__3262 (
            .O(N__15513),
            .I(N__15509));
    InMux I__3261 (
            .O(N__15512),
            .I(N__15506));
    LocalMux I__3260 (
            .O(N__15509),
            .I(G_184));
    LocalMux I__3259 (
            .O(N__15506),
            .I(G_184));
    CascadeMux I__3258 (
            .O(N__15501),
            .I(N__15497));
    InMux I__3257 (
            .O(N__15500),
            .I(N__15494));
    InMux I__3256 (
            .O(N__15497),
            .I(N__15490));
    LocalMux I__3255 (
            .O(N__15494),
            .I(N__15487));
    InMux I__3254 (
            .O(N__15493),
            .I(N__15484));
    LocalMux I__3253 (
            .O(N__15490),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    Odrv4 I__3252 (
            .O(N__15487),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    LocalMux I__3251 (
            .O(N__15484),
            .I(\Lab_UT.alarmstate_0_sqmuxa_1 ));
    InMux I__3250 (
            .O(N__15477),
            .I(N__15473));
    InMux I__3249 (
            .O(N__15476),
            .I(N__15470));
    LocalMux I__3248 (
            .O(N__15473),
            .I(N__15462));
    LocalMux I__3247 (
            .O(N__15470),
            .I(N__15462));
    InMux I__3246 (
            .O(N__15469),
            .I(N__15455));
    InMux I__3245 (
            .O(N__15468),
            .I(N__15455));
    InMux I__3244 (
            .O(N__15467),
            .I(N__15455));
    Odrv4 I__3243 (
            .O(N__15462),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    LocalMux I__3242 (
            .O(N__15455),
            .I(\Lab_UT.didp.di_Mtens_3 ));
    InMux I__3241 (
            .O(N__15450),
            .I(N__15447));
    LocalMux I__3240 (
            .O(N__15447),
            .I(\Lab_UT.didp.countrce2.q_5_3 ));
    InMux I__3239 (
            .O(N__15444),
            .I(N__15441));
    LocalMux I__3238 (
            .O(N__15441),
            .I(N__15438));
    Odrv4 I__3237 (
            .O(N__15438),
            .I(\Lab_UT.didp.countrce2.q_5_0 ));
    CascadeMux I__3236 (
            .O(N__15435),
            .I(N__15427));
    CascadeMux I__3235 (
            .O(N__15434),
            .I(N__15423));
    InMux I__3234 (
            .O(N__15433),
            .I(N__15414));
    InMux I__3233 (
            .O(N__15432),
            .I(N__15414));
    InMux I__3232 (
            .O(N__15431),
            .I(N__15414));
    InMux I__3231 (
            .O(N__15430),
            .I(N__15414));
    InMux I__3230 (
            .O(N__15427),
            .I(N__15408));
    InMux I__3229 (
            .O(N__15426),
            .I(N__15408));
    InMux I__3228 (
            .O(N__15423),
            .I(N__15405));
    LocalMux I__3227 (
            .O(N__15414),
            .I(N__15402));
    InMux I__3226 (
            .O(N__15413),
            .I(N__15399));
    LocalMux I__3225 (
            .O(N__15408),
            .I(N__15396));
    LocalMux I__3224 (
            .O(N__15405),
            .I(\Lab_UT.didp.di_Stens_0 ));
    Odrv4 I__3223 (
            .O(N__15402),
            .I(\Lab_UT.didp.di_Stens_0 ));
    LocalMux I__3222 (
            .O(N__15399),
            .I(\Lab_UT.didp.di_Stens_0 ));
    Odrv4 I__3221 (
            .O(N__15396),
            .I(\Lab_UT.didp.di_Stens_0 ));
    CascadeMux I__3220 (
            .O(N__15387),
            .I(N__15382));
    InMux I__3219 (
            .O(N__15386),
            .I(N__15375));
    InMux I__3218 (
            .O(N__15385),
            .I(N__15372));
    InMux I__3217 (
            .O(N__15382),
            .I(N__15369));
    InMux I__3216 (
            .O(N__15381),
            .I(N__15364));
    InMux I__3215 (
            .O(N__15380),
            .I(N__15364));
    InMux I__3214 (
            .O(N__15379),
            .I(N__15359));
    InMux I__3213 (
            .O(N__15378),
            .I(N__15359));
    LocalMux I__3212 (
            .O(N__15375),
            .I(N__15356));
    LocalMux I__3211 (
            .O(N__15372),
            .I(N__15353));
    LocalMux I__3210 (
            .O(N__15369),
            .I(\Lab_UT.didp.di_Stens_1 ));
    LocalMux I__3209 (
            .O(N__15364),
            .I(\Lab_UT.didp.di_Stens_1 ));
    LocalMux I__3208 (
            .O(N__15359),
            .I(\Lab_UT.didp.di_Stens_1 ));
    Odrv12 I__3207 (
            .O(N__15356),
            .I(\Lab_UT.didp.di_Stens_1 ));
    Odrv4 I__3206 (
            .O(N__15353),
            .I(\Lab_UT.didp.di_Stens_1 ));
    InMux I__3205 (
            .O(N__15342),
            .I(N__15335));
    InMux I__3204 (
            .O(N__15341),
            .I(N__15332));
    InMux I__3203 (
            .O(N__15340),
            .I(N__15329));
    InMux I__3202 (
            .O(N__15339),
            .I(N__15326));
    InMux I__3201 (
            .O(N__15338),
            .I(N__15323));
    LocalMux I__3200 (
            .O(N__15335),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3199 (
            .O(N__15332),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3198 (
            .O(N__15329),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3197 (
            .O(N__15326),
            .I(\Lab_UT.didp.di_Stens_3 ));
    LocalMux I__3196 (
            .O(N__15323),
            .I(\Lab_UT.didp.di_Stens_3 ));
    InMux I__3195 (
            .O(N__15312),
            .I(N__15309));
    LocalMux I__3194 (
            .O(N__15309),
            .I(\Lab_UT.didp.regrce3.did_alarmMatch_3 ));
    InMux I__3193 (
            .O(N__15306),
            .I(N__15303));
    LocalMux I__3192 (
            .O(N__15303),
            .I(\Lab_UT.didp.did_alarmMatch_0 ));
    CascadeMux I__3191 (
            .O(N__15300),
            .I(\Lab_UT.didp.did_alarmMatch_1_cascade_ ));
    InMux I__3190 (
            .O(N__15297),
            .I(N__15294));
    LocalMux I__3189 (
            .O(N__15294),
            .I(N__15291));
    Odrv4 I__3188 (
            .O(N__15291),
            .I(\Lab_UT.didp.did_alarmMatch_2 ));
    CascadeMux I__3187 (
            .O(N__15288),
            .I(N__15283));
    InMux I__3186 (
            .O(N__15287),
            .I(N__15277));
    InMux I__3185 (
            .O(N__15286),
            .I(N__15277));
    InMux I__3184 (
            .O(N__15283),
            .I(N__15272));
    InMux I__3183 (
            .O(N__15282),
            .I(N__15272));
    LocalMux I__3182 (
            .O(N__15277),
            .I(N__15267));
    LocalMux I__3181 (
            .O(N__15272),
            .I(N__15267));
    Span4Mux_v I__3180 (
            .O(N__15267),
            .I(N__15264));
    Odrv4 I__3179 (
            .O(N__15264),
            .I(\Lab_UT.didp.un1_dicLdStens_0 ));
    CascadeMux I__3178 (
            .O(N__15261),
            .I(N__15256));
    CascadeMux I__3177 (
            .O(N__15260),
            .I(N__15253));
    InMux I__3176 (
            .O(N__15259),
            .I(N__15247));
    InMux I__3175 (
            .O(N__15256),
            .I(N__15247));
    InMux I__3174 (
            .O(N__15253),
            .I(N__15242));
    InMux I__3173 (
            .O(N__15252),
            .I(N__15242));
    LocalMux I__3172 (
            .O(N__15247),
            .I(N__15239));
    LocalMux I__3171 (
            .O(N__15242),
            .I(N__15236));
    Span4Mux_h I__3170 (
            .O(N__15239),
            .I(N__15233));
    Odrv4 I__3169 (
            .O(N__15236),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    Odrv4 I__3168 (
            .O(N__15233),
            .I(\Lab_UT.didp.resetZ0Z_1 ));
    CascadeMux I__3167 (
            .O(N__15228),
            .I(N__15223));
    CascadeMux I__3166 (
            .O(N__15227),
            .I(N__15220));
    CascadeMux I__3165 (
            .O(N__15226),
            .I(N__15215));
    InMux I__3164 (
            .O(N__15223),
            .I(N__15208));
    InMux I__3163 (
            .O(N__15220),
            .I(N__15208));
    InMux I__3162 (
            .O(N__15219),
            .I(N__15208));
    InMux I__3161 (
            .O(N__15218),
            .I(N__15203));
    InMux I__3160 (
            .O(N__15215),
            .I(N__15203));
    LocalMux I__3159 (
            .O(N__15208),
            .I(\Lab_UT.didp.un24_ce_2 ));
    LocalMux I__3158 (
            .O(N__15203),
            .I(\Lab_UT.didp.un24_ce_2 ));
    InMux I__3157 (
            .O(N__15198),
            .I(N__15193));
    InMux I__3156 (
            .O(N__15197),
            .I(N__15190));
    CascadeMux I__3155 (
            .O(N__15196),
            .I(N__15185));
    LocalMux I__3154 (
            .O(N__15193),
            .I(N__15179));
    LocalMux I__3153 (
            .O(N__15190),
            .I(N__15179));
    InMux I__3152 (
            .O(N__15189),
            .I(N__15176));
    InMux I__3151 (
            .O(N__15188),
            .I(N__15171));
    InMux I__3150 (
            .O(N__15185),
            .I(N__15171));
    InMux I__3149 (
            .O(N__15184),
            .I(N__15168));
    Span4Mux_s2_v I__3148 (
            .O(N__15179),
            .I(N__15163));
    LocalMux I__3147 (
            .O(N__15176),
            .I(N__15163));
    LocalMux I__3146 (
            .O(N__15171),
            .I(N__15158));
    LocalMux I__3145 (
            .O(N__15168),
            .I(N__15158));
    Odrv4 I__3144 (
            .O(N__15163),
            .I(\Lab_UT.LdMtens ));
    Odrv12 I__3143 (
            .O(N__15158),
            .I(\Lab_UT.LdMtens ));
    CascadeMux I__3142 (
            .O(N__15153),
            .I(N__15150));
    InMux I__3141 (
            .O(N__15150),
            .I(N__15147));
    LocalMux I__3140 (
            .O(N__15147),
            .I(N__15144));
    Span4Mux_h I__3139 (
            .O(N__15144),
            .I(N__15141));
    Odrv4 I__3138 (
            .O(N__15141),
            .I(\Lab_UT.didp.countrce4.un20_qPone ));
    InMux I__3137 (
            .O(N__15138),
            .I(N__15133));
    InMux I__3136 (
            .O(N__15137),
            .I(N__15130));
    InMux I__3135 (
            .O(N__15136),
            .I(N__15127));
    LocalMux I__3134 (
            .O(N__15133),
            .I(N__15124));
    LocalMux I__3133 (
            .O(N__15130),
            .I(N__15119));
    LocalMux I__3132 (
            .O(N__15127),
            .I(N__15119));
    Span4Mux_v I__3131 (
            .O(N__15124),
            .I(N__15113));
    Span4Mux_v I__3130 (
            .O(N__15119),
            .I(N__15113));
    InMux I__3129 (
            .O(N__15118),
            .I(N__15110));
    Odrv4 I__3128 (
            .O(N__15113),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    LocalMux I__3127 (
            .O(N__15110),
            .I(\Lab_UT.didp.resetZ0Z_3 ));
    CascadeMux I__3126 (
            .O(N__15105),
            .I(\Lab_UT.didp.countrce4.q_5_3_cascade_ ));
    InMux I__3125 (
            .O(N__15102),
            .I(N__15099));
    LocalMux I__3124 (
            .O(N__15099),
            .I(N__15094));
    InMux I__3123 (
            .O(N__15098),
            .I(N__15089));
    InMux I__3122 (
            .O(N__15097),
            .I(N__15089));
    Span4Mux_h I__3121 (
            .O(N__15094),
            .I(N__15086));
    LocalMux I__3120 (
            .O(N__15089),
            .I(N__15083));
    Odrv4 I__3119 (
            .O(N__15086),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    Odrv4 I__3118 (
            .O(N__15083),
            .I(\Lab_UT.didp.un1_dicLdMtens_0 ));
    InMux I__3117 (
            .O(N__15078),
            .I(N__15075));
    LocalMux I__3116 (
            .O(N__15075),
            .I(\Lab_UT.didp.countrce2.q_5_1 ));
    CascadeMux I__3115 (
            .O(N__15072),
            .I(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ));
    InMux I__3114 (
            .O(N__15069),
            .I(N__15066));
    LocalMux I__3113 (
            .O(N__15066),
            .I(\Lab_UT.didp.reset_12_1_3 ));
    InMux I__3112 (
            .O(N__15063),
            .I(N__15057));
    InMux I__3111 (
            .O(N__15062),
            .I(N__15052));
    InMux I__3110 (
            .O(N__15061),
            .I(N__15052));
    InMux I__3109 (
            .O(N__15060),
            .I(N__15047));
    LocalMux I__3108 (
            .O(N__15057),
            .I(N__15044));
    LocalMux I__3107 (
            .O(N__15052),
            .I(N__15041));
    InMux I__3106 (
            .O(N__15051),
            .I(N__15036));
    InMux I__3105 (
            .O(N__15050),
            .I(N__15036));
    LocalMux I__3104 (
            .O(N__15047),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    Odrv4 I__3103 (
            .O(N__15044),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    Odrv12 I__3102 (
            .O(N__15041),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    LocalMux I__3101 (
            .O(N__15036),
            .I(\Lab_UT.didp.di_Mtens_2 ));
    CascadeMux I__3100 (
            .O(N__15027),
            .I(\Lab_UT.didp.ce_12_3_cascade_ ));
    CascadeMux I__3099 (
            .O(N__15024),
            .I(N__15021));
    InMux I__3098 (
            .O(N__15021),
            .I(N__15006));
    InMux I__3097 (
            .O(N__15020),
            .I(N__15006));
    InMux I__3096 (
            .O(N__15019),
            .I(N__14992));
    InMux I__3095 (
            .O(N__15018),
            .I(N__14992));
    InMux I__3094 (
            .O(N__15017),
            .I(N__14992));
    InMux I__3093 (
            .O(N__15016),
            .I(N__14992));
    InMux I__3092 (
            .O(N__15015),
            .I(N__14992));
    InMux I__3091 (
            .O(N__15014),
            .I(N__14992));
    InMux I__3090 (
            .O(N__15013),
            .I(N__14989));
    InMux I__3089 (
            .O(N__15012),
            .I(N__14986));
    InMux I__3088 (
            .O(N__15011),
            .I(N__14983));
    LocalMux I__3087 (
            .O(N__15006),
            .I(N__14980));
    InMux I__3086 (
            .O(N__15005),
            .I(N__14977));
    LocalMux I__3085 (
            .O(N__14992),
            .I(N__14972));
    LocalMux I__3084 (
            .O(N__14989),
            .I(N__14972));
    LocalMux I__3083 (
            .O(N__14986),
            .I(N__14969));
    LocalMux I__3082 (
            .O(N__14983),
            .I(N__14966));
    Span4Mux_v I__3081 (
            .O(N__14980),
            .I(N__14960));
    LocalMux I__3080 (
            .O(N__14977),
            .I(N__14960));
    Span4Mux_s2_v I__3079 (
            .O(N__14972),
            .I(N__14957));
    Span4Mux_h I__3078 (
            .O(N__14969),
            .I(N__14952));
    Span4Mux_h I__3077 (
            .O(N__14966),
            .I(N__14952));
    InMux I__3076 (
            .O(N__14965),
            .I(N__14949));
    Span4Mux_h I__3075 (
            .O(N__14960),
            .I(N__14944));
    Span4Mux_h I__3074 (
            .O(N__14957),
            .I(N__14944));
    Odrv4 I__3073 (
            .O(N__14952),
            .I(oneSecStrb));
    LocalMux I__3072 (
            .O(N__14949),
            .I(oneSecStrb));
    Odrv4 I__3071 (
            .O(N__14944),
            .I(oneSecStrb));
    CascadeMux I__3070 (
            .O(N__14937),
            .I(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ));
    InMux I__3069 (
            .O(N__14934),
            .I(N__14931));
    LocalMux I__3068 (
            .O(N__14931),
            .I(\Lab_UT.didp.countrce4.q_5_0 ));
    CascadeMux I__3067 (
            .O(N__14928),
            .I(N__14925));
    InMux I__3066 (
            .O(N__14925),
            .I(N__14921));
    InMux I__3065 (
            .O(N__14924),
            .I(N__14918));
    LocalMux I__3064 (
            .O(N__14921),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    LocalMux I__3063 (
            .O(N__14918),
            .I(\Lab_UT.didp.ceZ0Z_3 ));
    CascadeMux I__3062 (
            .O(N__14913),
            .I(\Lab_UT.dictrl.g0_17_0_cascade_ ));
    InMux I__3061 (
            .O(N__14910),
            .I(N__14907));
    LocalMux I__3060 (
            .O(N__14907),
            .I(N__14904));
    Odrv4 I__3059 (
            .O(N__14904),
            .I(\Lab_UT.dictrl.g2_0_0 ));
    CascadeMux I__3058 (
            .O(N__14901),
            .I(N__14897));
    InMux I__3057 (
            .O(N__14900),
            .I(N__14891));
    InMux I__3056 (
            .O(N__14897),
            .I(N__14891));
    InMux I__3055 (
            .O(N__14896),
            .I(N__14888));
    LocalMux I__3054 (
            .O(N__14891),
            .I(N__14883));
    LocalMux I__3053 (
            .O(N__14888),
            .I(N__14883));
    Odrv4 I__3052 (
            .O(N__14883),
            .I(bu_rx_data_fast_3));
    CascadeMux I__3051 (
            .O(N__14880),
            .I(\Lab_UT.dictrl.g0_2Z0Z_5_cascade_ ));
    InMux I__3050 (
            .O(N__14877),
            .I(N__14874));
    LocalMux I__3049 (
            .O(N__14874),
            .I(N__14871));
    Odrv4 I__3048 (
            .O(N__14871),
            .I(\Lab_UT.dictrl.g2_0 ));
    InMux I__3047 (
            .O(N__14868),
            .I(N__14865));
    LocalMux I__3046 (
            .O(N__14865),
            .I(\Lab_UT.dictrl.g1_1 ));
    CascadeMux I__3045 (
            .O(N__14862),
            .I(\Lab_UT.dictrl.g2_0_cascade_ ));
    InMux I__3044 (
            .O(N__14859),
            .I(N__14856));
    LocalMux I__3043 (
            .O(N__14856),
            .I(\Lab_UT.dictrl.N_90_0_0_0 ));
    InMux I__3042 (
            .O(N__14853),
            .I(N__14850));
    LocalMux I__3041 (
            .O(N__14850),
            .I(\Lab_UT.dictrl.m40_N_5_mux_0 ));
    CascadeMux I__3040 (
            .O(N__14847),
            .I(\Lab_UT.dictrl.g2Z0Z_1_cascade_ ));
    InMux I__3039 (
            .O(N__14844),
            .I(N__14841));
    LocalMux I__3038 (
            .O(N__14841),
            .I(N__14838));
    Span4Mux_h I__3037 (
            .O(N__14838),
            .I(N__14834));
    InMux I__3036 (
            .O(N__14837),
            .I(N__14831));
    Odrv4 I__3035 (
            .O(N__14834),
            .I(\Lab_UT.dictrl.g1_0 ));
    LocalMux I__3034 (
            .O(N__14831),
            .I(\Lab_UT.dictrl.g1_0 ));
    InMux I__3033 (
            .O(N__14826),
            .I(N__14823));
    LocalMux I__3032 (
            .O(N__14823),
            .I(\Lab_UT.dictrl.g0_17_a6_2_1 ));
    InMux I__3031 (
            .O(N__14820),
            .I(N__14817));
    LocalMux I__3030 (
            .O(N__14817),
            .I(N__14814));
    Odrv12 I__3029 (
            .O(N__14814),
            .I(\Lab_UT.dictrl.g0_17_a6_3_6 ));
    InMux I__3028 (
            .O(N__14811),
            .I(N__14808));
    LocalMux I__3027 (
            .O(N__14808),
            .I(\Lab_UT.dictrl.g0_17_a6_3_8 ));
    CascadeMux I__3026 (
            .O(N__14805),
            .I(\Lab_UT.dictrl.N_22_cascade_ ));
    InMux I__3025 (
            .O(N__14802),
            .I(N__14790));
    InMux I__3024 (
            .O(N__14801),
            .I(N__14790));
    InMux I__3023 (
            .O(N__14800),
            .I(N__14790));
    InMux I__3022 (
            .O(N__14799),
            .I(N__14790));
    LocalMux I__3021 (
            .O(N__14790),
            .I(N__14787));
    Odrv4 I__3020 (
            .O(N__14787),
            .I(\Lab_UT.dictrl.N_90_0 ));
    CascadeMux I__3019 (
            .O(N__14784),
            .I(N__14778));
    CascadeMux I__3018 (
            .O(N__14783),
            .I(N__14775));
    CascadeMux I__3017 (
            .O(N__14782),
            .I(N__14772));
    CascadeMux I__3016 (
            .O(N__14781),
            .I(N__14769));
    InMux I__3015 (
            .O(N__14778),
            .I(N__14764));
    InMux I__3014 (
            .O(N__14775),
            .I(N__14764));
    InMux I__3013 (
            .O(N__14772),
            .I(N__14759));
    InMux I__3012 (
            .O(N__14769),
            .I(N__14759));
    LocalMux I__3011 (
            .O(N__14764),
            .I(N__14754));
    LocalMux I__3010 (
            .O(N__14759),
            .I(N__14754));
    Odrv12 I__3009 (
            .O(N__14754),
            .I(\Lab_UT.dictrl.N_95_0 ));
    CascadeMux I__3008 (
            .O(N__14751),
            .I(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ));
    InMux I__3007 (
            .O(N__14748),
            .I(N__14745));
    LocalMux I__3006 (
            .O(N__14745),
            .I(N__14742));
    Odrv12 I__3005 (
            .O(N__14742),
            .I(\Lab_UT.LdStens_i_3 ));
    CascadeMux I__3004 (
            .O(N__14739),
            .I(N__14735));
    CascadeMux I__3003 (
            .O(N__14738),
            .I(N__14731));
    InMux I__3002 (
            .O(N__14735),
            .I(N__14728));
    InMux I__3001 (
            .O(N__14734),
            .I(N__14725));
    InMux I__3000 (
            .O(N__14731),
            .I(N__14722));
    LocalMux I__2999 (
            .O(N__14728),
            .I(N__14717));
    LocalMux I__2998 (
            .O(N__14725),
            .I(N__14717));
    LocalMux I__2997 (
            .O(N__14722),
            .I(\Lab_UT.dictrl.state_fast_1 ));
    Odrv4 I__2996 (
            .O(N__14717),
            .I(\Lab_UT.dictrl.state_fast_1 ));
    CascadeMux I__2995 (
            .O(N__14712),
            .I(\Lab_UT.dictrl.N_95_0_0_cascade_ ));
    CascadeMux I__2994 (
            .O(N__14709),
            .I(\Lab_UT.dictrl.g0_3_0_cascade_ ));
    CascadeMux I__2993 (
            .O(N__14706),
            .I(\Lab_UT.dictrl.g4_cascade_ ));
    CascadeMux I__2992 (
            .O(N__14703),
            .I(\Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_ ));
    InMux I__2991 (
            .O(N__14700),
            .I(N__14697));
    LocalMux I__2990 (
            .O(N__14697),
            .I(\Lab_UT.dictrl.g2_5 ));
    InMux I__2989 (
            .O(N__14694),
            .I(N__14688));
    InMux I__2988 (
            .O(N__14693),
            .I(N__14681));
    InMux I__2987 (
            .O(N__14692),
            .I(N__14681));
    InMux I__2986 (
            .O(N__14691),
            .I(N__14681));
    LocalMux I__2985 (
            .O(N__14688),
            .I(N__14678));
    LocalMux I__2984 (
            .O(N__14681),
            .I(\Lab_UT.dicRun_2 ));
    Odrv4 I__2983 (
            .O(N__14678),
            .I(\Lab_UT.dicRun_2 ));
    InMux I__2982 (
            .O(N__14673),
            .I(N__14670));
    LocalMux I__2981 (
            .O(N__14670),
            .I(\Lab_UT.didp.ceZ0Z_0 ));
    InMux I__2980 (
            .O(N__14667),
            .I(N__14664));
    LocalMux I__2979 (
            .O(N__14664),
            .I(\Lab_UT.didp.ceZ0Z_1 ));
    InMux I__2978 (
            .O(N__14661),
            .I(N__14655));
    InMux I__2977 (
            .O(N__14660),
            .I(N__14655));
    LocalMux I__2976 (
            .O(N__14655),
            .I(N__14650));
    InMux I__2975 (
            .O(N__14654),
            .I(N__14647));
    InMux I__2974 (
            .O(N__14653),
            .I(N__14644));
    Span4Mux_h I__2973 (
            .O(N__14650),
            .I(N__14641));
    LocalMux I__2972 (
            .O(N__14647),
            .I(N__14636));
    LocalMux I__2971 (
            .O(N__14644),
            .I(N__14636));
    Span4Mux_h I__2970 (
            .O(N__14641),
            .I(N__14633));
    Span4Mux_h I__2969 (
            .O(N__14636),
            .I(N__14630));
    Odrv4 I__2968 (
            .O(N__14633),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    Odrv4 I__2967 (
            .O(N__14630),
            .I(\buart.Z_rx.hhZ0Z_1 ));
    InMux I__2966 (
            .O(N__14625),
            .I(N__14622));
    LocalMux I__2965 (
            .O(N__14622),
            .I(\Lab_UT.un1_idle_1_0_iclkZ0 ));
    CascadeMux I__2964 (
            .O(N__14619),
            .I(G_186_cascade_));
    InMux I__2963 (
            .O(N__14616),
            .I(N__14611));
    InMux I__2962 (
            .O(N__14615),
            .I(N__14606));
    InMux I__2961 (
            .O(N__14614),
            .I(N__14606));
    LocalMux I__2960 (
            .O(N__14611),
            .I(G_191));
    LocalMux I__2959 (
            .O(N__14606),
            .I(G_191));
    CascadeMux I__2958 (
            .O(N__14601),
            .I(\Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_ ));
    InMux I__2957 (
            .O(N__14598),
            .I(N__14595));
    LocalMux I__2956 (
            .O(N__14595),
            .I(N__14592));
    Odrv4 I__2955 (
            .O(N__14592),
            .I(\Lab_UT.dictrl.G_10_1 ));
    CascadeMux I__2954 (
            .O(N__14589),
            .I(\Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ));
    CascadeMux I__2953 (
            .O(N__14586),
            .I(\Lab_UT.dictrl.N_21_0_cascade_ ));
    InMux I__2952 (
            .O(N__14583),
            .I(N__14573));
    InMux I__2951 (
            .O(N__14582),
            .I(N__14573));
    InMux I__2950 (
            .O(N__14581),
            .I(N__14573));
    InMux I__2949 (
            .O(N__14580),
            .I(N__14558));
    LocalMux I__2948 (
            .O(N__14573),
            .I(N__14555));
    InMux I__2947 (
            .O(N__14572),
            .I(N__14548));
    InMux I__2946 (
            .O(N__14571),
            .I(N__14548));
    InMux I__2945 (
            .O(N__14570),
            .I(N__14548));
    InMux I__2944 (
            .O(N__14569),
            .I(N__14539));
    InMux I__2943 (
            .O(N__14568),
            .I(N__14539));
    InMux I__2942 (
            .O(N__14567),
            .I(N__14539));
    InMux I__2941 (
            .O(N__14566),
            .I(N__14539));
    InMux I__2940 (
            .O(N__14565),
            .I(N__14536));
    InMux I__2939 (
            .O(N__14564),
            .I(N__14531));
    InMux I__2938 (
            .O(N__14563),
            .I(N__14531));
    InMux I__2937 (
            .O(N__14562),
            .I(N__14526));
    InMux I__2936 (
            .O(N__14561),
            .I(N__14526));
    LocalMux I__2935 (
            .O(N__14558),
            .I(N__14521));
    Span4Mux_s1_v I__2934 (
            .O(N__14555),
            .I(N__14521));
    LocalMux I__2933 (
            .O(N__14548),
            .I(N__14518));
    LocalMux I__2932 (
            .O(N__14539),
            .I(N__14515));
    LocalMux I__2931 (
            .O(N__14536),
            .I(\Lab_UT.i16_mux ));
    LocalMux I__2930 (
            .O(N__14531),
            .I(\Lab_UT.i16_mux ));
    LocalMux I__2929 (
            .O(N__14526),
            .I(\Lab_UT.i16_mux ));
    Odrv4 I__2928 (
            .O(N__14521),
            .I(\Lab_UT.i16_mux ));
    Odrv12 I__2927 (
            .O(N__14518),
            .I(\Lab_UT.i16_mux ));
    Odrv12 I__2926 (
            .O(N__14515),
            .I(\Lab_UT.i16_mux ));
    InMux I__2925 (
            .O(N__14502),
            .I(N__14499));
    LocalMux I__2924 (
            .O(N__14499),
            .I(\Lab_UT.dictrl.i18_mux ));
    InMux I__2923 (
            .O(N__14496),
            .I(N__14493));
    LocalMux I__2922 (
            .O(N__14493),
            .I(\Lab_UT.dispString.dOut_RNO_1Z0Z_1 ));
    CascadeMux I__2921 (
            .O(N__14490),
            .I(N__14484));
    CascadeMux I__2920 (
            .O(N__14489),
            .I(N__14477));
    CascadeMux I__2919 (
            .O(N__14488),
            .I(N__14473));
    InMux I__2918 (
            .O(N__14487),
            .I(N__14466));
    InMux I__2917 (
            .O(N__14484),
            .I(N__14466));
    InMux I__2916 (
            .O(N__14483),
            .I(N__14459));
    InMux I__2915 (
            .O(N__14482),
            .I(N__14459));
    InMux I__2914 (
            .O(N__14481),
            .I(N__14459));
    InMux I__2913 (
            .O(N__14480),
            .I(N__14450));
    InMux I__2912 (
            .O(N__14477),
            .I(N__14447));
    InMux I__2911 (
            .O(N__14476),
            .I(N__14442));
    InMux I__2910 (
            .O(N__14473),
            .I(N__14442));
    InMux I__2909 (
            .O(N__14472),
            .I(N__14436));
    InMux I__2908 (
            .O(N__14471),
            .I(N__14436));
    LocalMux I__2907 (
            .O(N__14466),
            .I(N__14433));
    LocalMux I__2906 (
            .O(N__14459),
            .I(N__14430));
    InMux I__2905 (
            .O(N__14458),
            .I(N__14425));
    InMux I__2904 (
            .O(N__14457),
            .I(N__14425));
    InMux I__2903 (
            .O(N__14456),
            .I(N__14422));
    InMux I__2902 (
            .O(N__14455),
            .I(N__14415));
    InMux I__2901 (
            .O(N__14454),
            .I(N__14415));
    InMux I__2900 (
            .O(N__14453),
            .I(N__14415));
    LocalMux I__2899 (
            .O(N__14450),
            .I(N__14408));
    LocalMux I__2898 (
            .O(N__14447),
            .I(N__14408));
    LocalMux I__2897 (
            .O(N__14442),
            .I(N__14408));
    InMux I__2896 (
            .O(N__14441),
            .I(N__14404));
    LocalMux I__2895 (
            .O(N__14436),
            .I(N__14399));
    Span4Mux_h I__2894 (
            .O(N__14433),
            .I(N__14399));
    Span4Mux_h I__2893 (
            .O(N__14430),
            .I(N__14394));
    LocalMux I__2892 (
            .O(N__14425),
            .I(N__14394));
    LocalMux I__2891 (
            .O(N__14422),
            .I(N__14391));
    LocalMux I__2890 (
            .O(N__14415),
            .I(N__14386));
    Span4Mux_v I__2889 (
            .O(N__14408),
            .I(N__14386));
    InMux I__2888 (
            .O(N__14407),
            .I(N__14383));
    LocalMux I__2887 (
            .O(N__14404),
            .I(N__14376));
    Span4Mux_v I__2886 (
            .O(N__14399),
            .I(N__14376));
    Span4Mux_h I__2885 (
            .O(N__14394),
            .I(N__14376));
    Odrv12 I__2884 (
            .O(N__14391),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2883 (
            .O(N__14386),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    LocalMux I__2882 (
            .O(N__14383),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    Odrv4 I__2881 (
            .O(N__14376),
            .I(\Lab_UT.dispString.cntZ0Z_0 ));
    InMux I__2880 (
            .O(N__14367),
            .I(N__14358));
    CascadeMux I__2879 (
            .O(N__14366),
            .I(N__14353));
    InMux I__2878 (
            .O(N__14365),
            .I(N__14350));
    CascadeMux I__2877 (
            .O(N__14364),
            .I(N__14347));
    CascadeMux I__2876 (
            .O(N__14363),
            .I(N__14344));
    InMux I__2875 (
            .O(N__14362),
            .I(N__14341));
    CascadeMux I__2874 (
            .O(N__14361),
            .I(N__14337));
    LocalMux I__2873 (
            .O(N__14358),
            .I(N__14331));
    InMux I__2872 (
            .O(N__14357),
            .I(N__14324));
    InMux I__2871 (
            .O(N__14356),
            .I(N__14324));
    InMux I__2870 (
            .O(N__14353),
            .I(N__14324));
    LocalMux I__2869 (
            .O(N__14350),
            .I(N__14321));
    InMux I__2868 (
            .O(N__14347),
            .I(N__14316));
    InMux I__2867 (
            .O(N__14344),
            .I(N__14316));
    LocalMux I__2866 (
            .O(N__14341),
            .I(N__14313));
    InMux I__2865 (
            .O(N__14340),
            .I(N__14303));
    InMux I__2864 (
            .O(N__14337),
            .I(N__14303));
    InMux I__2863 (
            .O(N__14336),
            .I(N__14303));
    InMux I__2862 (
            .O(N__14335),
            .I(N__14298));
    InMux I__2861 (
            .O(N__14334),
            .I(N__14298));
    Span4Mux_h I__2860 (
            .O(N__14331),
            .I(N__14292));
    LocalMux I__2859 (
            .O(N__14324),
            .I(N__14292));
    Span4Mux_v I__2858 (
            .O(N__14321),
            .I(N__14287));
    LocalMux I__2857 (
            .O(N__14316),
            .I(N__14287));
    Span4Mux_h I__2856 (
            .O(N__14313),
            .I(N__14284));
    InMux I__2855 (
            .O(N__14312),
            .I(N__14277));
    InMux I__2854 (
            .O(N__14311),
            .I(N__14277));
    InMux I__2853 (
            .O(N__14310),
            .I(N__14277));
    LocalMux I__2852 (
            .O(N__14303),
            .I(N__14272));
    LocalMux I__2851 (
            .O(N__14298),
            .I(N__14272));
    InMux I__2850 (
            .O(N__14297),
            .I(N__14269));
    Span4Mux_v I__2849 (
            .O(N__14292),
            .I(N__14264));
    Span4Mux_h I__2848 (
            .O(N__14287),
            .I(N__14264));
    Odrv4 I__2847 (
            .O(N__14284),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2846 (
            .O(N__14277),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv12 I__2845 (
            .O(N__14272),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    LocalMux I__2844 (
            .O(N__14269),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    Odrv4 I__2843 (
            .O(N__14264),
            .I(\Lab_UT.dispString.cntZ0Z_1 ));
    InMux I__2842 (
            .O(N__14253),
            .I(N__14250));
    LocalMux I__2841 (
            .O(N__14250),
            .I(N__14247));
    Span4Mux_h I__2840 (
            .O(N__14247),
            .I(N__14244));
    Odrv4 I__2839 (
            .O(N__14244),
            .I(\Lab_UT.dispString.m49_ns_1 ));
    CascadeMux I__2838 (
            .O(N__14241),
            .I(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ));
    CascadeMux I__2837 (
            .O(N__14238),
            .I(\Lab_UT.didp.countrce1.q_5_3_cascade_ ));
    CascadeMux I__2836 (
            .O(N__14235),
            .I(N__14226));
    CascadeMux I__2835 (
            .O(N__14234),
            .I(N__14223));
    CascadeMux I__2834 (
            .O(N__14233),
            .I(N__14220));
    CascadeMux I__2833 (
            .O(N__14232),
            .I(N__14217));
    CascadeMux I__2832 (
            .O(N__14231),
            .I(N__14214));
    CascadeMux I__2831 (
            .O(N__14230),
            .I(N__14211));
    CascadeMux I__2830 (
            .O(N__14229),
            .I(N__14208));
    InMux I__2829 (
            .O(N__14226),
            .I(N__14199));
    InMux I__2828 (
            .O(N__14223),
            .I(N__14199));
    InMux I__2827 (
            .O(N__14220),
            .I(N__14199));
    InMux I__2826 (
            .O(N__14217),
            .I(N__14199));
    InMux I__2825 (
            .O(N__14214),
            .I(N__14196));
    InMux I__2824 (
            .O(N__14211),
            .I(N__14191));
    InMux I__2823 (
            .O(N__14208),
            .I(N__14191));
    LocalMux I__2822 (
            .O(N__14199),
            .I(\Lab_UT.sec1_3 ));
    LocalMux I__2821 (
            .O(N__14196),
            .I(\Lab_UT.sec1_3 ));
    LocalMux I__2820 (
            .O(N__14191),
            .I(\Lab_UT.sec1_3 ));
    InMux I__2819 (
            .O(N__14184),
            .I(N__14181));
    LocalMux I__2818 (
            .O(N__14181),
            .I(N__14176));
    InMux I__2817 (
            .O(N__14180),
            .I(N__14173));
    InMux I__2816 (
            .O(N__14179),
            .I(N__14170));
    Odrv4 I__2815 (
            .O(N__14176),
            .I(\Lab_UT.di_AMtens_1 ));
    LocalMux I__2814 (
            .O(N__14173),
            .I(\Lab_UT.di_AMtens_1 ));
    LocalMux I__2813 (
            .O(N__14170),
            .I(\Lab_UT.di_AMtens_1 ));
    InMux I__2812 (
            .O(N__14163),
            .I(N__14160));
    LocalMux I__2811 (
            .O(N__14160),
            .I(N__14156));
    InMux I__2810 (
            .O(N__14159),
            .I(N__14152));
    Span4Mux_s0_v I__2809 (
            .O(N__14156),
            .I(N__14149));
    InMux I__2808 (
            .O(N__14155),
            .I(N__14146));
    LocalMux I__2807 (
            .O(N__14152),
            .I(\Lab_UT.di_AMtens_2 ));
    Odrv4 I__2806 (
            .O(N__14149),
            .I(\Lab_UT.di_AMtens_2 ));
    LocalMux I__2805 (
            .O(N__14146),
            .I(\Lab_UT.di_AMtens_2 ));
    CascadeMux I__2804 (
            .O(N__14139),
            .I(\Lab_UT.didp.countrce4.q_5_1_cascade_ ));
    InMux I__2803 (
            .O(N__14136),
            .I(N__14129));
    InMux I__2802 (
            .O(N__14135),
            .I(N__14126));
    CascadeMux I__2801 (
            .O(N__14134),
            .I(N__14121));
    InMux I__2800 (
            .O(N__14133),
            .I(N__14116));
    InMux I__2799 (
            .O(N__14132),
            .I(N__14116));
    LocalMux I__2798 (
            .O(N__14129),
            .I(N__14111));
    LocalMux I__2797 (
            .O(N__14126),
            .I(N__14111));
    InMux I__2796 (
            .O(N__14125),
            .I(N__14108));
    InMux I__2795 (
            .O(N__14124),
            .I(N__14103));
    InMux I__2794 (
            .O(N__14121),
            .I(N__14103));
    LocalMux I__2793 (
            .O(N__14116),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    Odrv4 I__2792 (
            .O(N__14111),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__2791 (
            .O(N__14108),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    LocalMux I__2790 (
            .O(N__14103),
            .I(\Lab_UT.didp.di_Mtens_1 ));
    CascadeMux I__2789 (
            .O(N__14094),
            .I(\Lab_UT.didp.countrce4.un13_qPone_cascade_ ));
    CascadeMux I__2788 (
            .O(N__14091),
            .I(\Lab_UT.didp.countrce4.q_5_2_cascade_ ));
    CascadeMux I__2787 (
            .O(N__14088),
            .I(\Lab_UT.dictrl.N_95_cascade_ ));
    InMux I__2786 (
            .O(N__14085),
            .I(N__14081));
    InMux I__2785 (
            .O(N__14084),
            .I(N__14078));
    LocalMux I__2784 (
            .O(N__14081),
            .I(N__14073));
    LocalMux I__2783 (
            .O(N__14078),
            .I(N__14070));
    InMux I__2782 (
            .O(N__14077),
            .I(N__14067));
    InMux I__2781 (
            .O(N__14076),
            .I(N__14064));
    Span4Mux_v I__2780 (
            .O(N__14073),
            .I(N__14052));
    Span4Mux_s2_h I__2779 (
            .O(N__14070),
            .I(N__14052));
    LocalMux I__2778 (
            .O(N__14067),
            .I(N__14052));
    LocalMux I__2777 (
            .O(N__14064),
            .I(N__14049));
    InMux I__2776 (
            .O(N__14063),
            .I(N__14038));
    InMux I__2775 (
            .O(N__14062),
            .I(N__14038));
    InMux I__2774 (
            .O(N__14061),
            .I(N__14038));
    InMux I__2773 (
            .O(N__14060),
            .I(N__14038));
    InMux I__2772 (
            .O(N__14059),
            .I(N__14038));
    Odrv4 I__2771 (
            .O(N__14052),
            .I(\uu2.N_101 ));
    Odrv4 I__2770 (
            .O(N__14049),
            .I(\uu2.N_101 ));
    LocalMux I__2769 (
            .O(N__14038),
            .I(\uu2.N_101 ));
    CascadeMux I__2768 (
            .O(N__14031),
            .I(N__14027));
    CascadeMux I__2767 (
            .O(N__14030),
            .I(N__14024));
    InMux I__2766 (
            .O(N__14027),
            .I(N__14020));
    InMux I__2765 (
            .O(N__14024),
            .I(N__14015));
    InMux I__2764 (
            .O(N__14023),
            .I(N__14015));
    LocalMux I__2763 (
            .O(N__14020),
            .I(N__14012));
    LocalMux I__2762 (
            .O(N__14015),
            .I(N__14009));
    Span4Mux_s2_v I__2761 (
            .O(N__14012),
            .I(N__14006));
    Span4Mux_v I__2760 (
            .O(N__14009),
            .I(N__14003));
    Odrv4 I__2759 (
            .O(N__14006),
            .I(\uu2.N_111 ));
    Odrv4 I__2758 (
            .O(N__14003),
            .I(\uu2.N_111 ));
    InMux I__2757 (
            .O(N__13998),
            .I(N__13994));
    InMux I__2756 (
            .O(N__13997),
            .I(N__13991));
    LocalMux I__2755 (
            .O(N__13994),
            .I(N__13987));
    LocalMux I__2754 (
            .O(N__13991),
            .I(N__13984));
    InMux I__2753 (
            .O(N__13990),
            .I(N__13981));
    Span4Mux_h I__2752 (
            .O(N__13987),
            .I(N__13977));
    Span4Mux_s1_h I__2751 (
            .O(N__13984),
            .I(N__13972));
    LocalMux I__2750 (
            .O(N__13981),
            .I(N__13972));
    InMux I__2749 (
            .O(N__13980),
            .I(N__13969));
    Odrv4 I__2748 (
            .O(N__13977),
            .I(\uu2.un28_w_addr_user_i_0 ));
    Odrv4 I__2747 (
            .O(N__13972),
            .I(\uu2.un28_w_addr_user_i_0 ));
    LocalMux I__2746 (
            .O(N__13969),
            .I(\uu2.un28_w_addr_user_i_0 ));
    CascadeMux I__2745 (
            .O(N__13962),
            .I(N__13959));
    InMux I__2744 (
            .O(N__13959),
            .I(N__13956));
    LocalMux I__2743 (
            .O(N__13956),
            .I(N__13950));
    InMux I__2742 (
            .O(N__13955),
            .I(N__13945));
    InMux I__2741 (
            .O(N__13954),
            .I(N__13945));
    InMux I__2740 (
            .O(N__13953),
            .I(N__13942));
    Span4Mux_v I__2739 (
            .O(N__13950),
            .I(N__13937));
    LocalMux I__2738 (
            .O(N__13945),
            .I(N__13937));
    LocalMux I__2737 (
            .O(N__13942),
            .I(N__13932));
    Span4Mux_h I__2736 (
            .O(N__13937),
            .I(N__13932));
    Odrv4 I__2735 (
            .O(N__13932),
            .I(\uu2.w_addr_userZ0Z_7 ));
    InMux I__2734 (
            .O(N__13929),
            .I(N__13925));
    InMux I__2733 (
            .O(N__13928),
            .I(N__13922));
    LocalMux I__2732 (
            .O(N__13925),
            .I(N__13919));
    LocalMux I__2731 (
            .O(N__13922),
            .I(N__13912));
    Span4Mux_s3_v I__2730 (
            .O(N__13919),
            .I(N__13909));
    InMux I__2729 (
            .O(N__13918),
            .I(N__13906));
    InMux I__2728 (
            .O(N__13917),
            .I(N__13901));
    InMux I__2727 (
            .O(N__13916),
            .I(N__13901));
    InMux I__2726 (
            .O(N__13915),
            .I(N__13898));
    Span4Mux_h I__2725 (
            .O(N__13912),
            .I(N__13893));
    Span4Mux_h I__2724 (
            .O(N__13909),
            .I(N__13893));
    LocalMux I__2723 (
            .O(N__13906),
            .I(N__13888));
    LocalMux I__2722 (
            .O(N__13901),
            .I(N__13888));
    LocalMux I__2721 (
            .O(N__13898),
            .I(o_One_Sec_Pulse));
    Odrv4 I__2720 (
            .O(N__13893),
            .I(o_One_Sec_Pulse));
    Odrv12 I__2719 (
            .O(N__13888),
            .I(o_One_Sec_Pulse));
    InMux I__2718 (
            .O(N__13881),
            .I(N__13878));
    LocalMux I__2717 (
            .O(N__13878),
            .I(\uu2.bitmapZ0Z_111 ));
    InMux I__2716 (
            .O(N__13875),
            .I(N__13872));
    LocalMux I__2715 (
            .O(N__13872),
            .I(N__13868));
    InMux I__2714 (
            .O(N__13871),
            .I(N__13865));
    Span4Mux_h I__2713 (
            .O(N__13868),
            .I(N__13862));
    LocalMux I__2712 (
            .O(N__13865),
            .I(N__13857));
    Span4Mux_v I__2711 (
            .O(N__13862),
            .I(N__13854));
    InMux I__2710 (
            .O(N__13861),
            .I(N__13849));
    InMux I__2709 (
            .O(N__13860),
            .I(N__13849));
    Span12Mux_s9_v I__2708 (
            .O(N__13857),
            .I(N__13846));
    Odrv4 I__2707 (
            .O(N__13854),
            .I(\uu2.vram_rd_clkZ0 ));
    LocalMux I__2706 (
            .O(N__13849),
            .I(\uu2.vram_rd_clkZ0 ));
    Odrv12 I__2705 (
            .O(N__13846),
            .I(\uu2.vram_rd_clkZ0 ));
    InMux I__2704 (
            .O(N__13839),
            .I(N__13836));
    LocalMux I__2703 (
            .O(N__13836),
            .I(N__13832));
    InMux I__2702 (
            .O(N__13835),
            .I(N__13829));
    Span4Mux_v I__2701 (
            .O(N__13832),
            .I(N__13826));
    LocalMux I__2700 (
            .O(N__13829),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    Odrv4 I__2699 (
            .O(N__13826),
            .I(\uu2.vram_rd_clk_detZ0Z_0 ));
    InMux I__2698 (
            .O(N__13821),
            .I(N__13818));
    LocalMux I__2697 (
            .O(N__13818),
            .I(N__13815));
    Span4Mux_v I__2696 (
            .O(N__13815),
            .I(N__13812));
    Span4Mux_s2_v I__2695 (
            .O(N__13812),
            .I(N__13809));
    Odrv4 I__2694 (
            .O(N__13809),
            .I(\uu2.vram_rd_clk_detZ0Z_1 ));
    InMux I__2693 (
            .O(N__13806),
            .I(N__13803));
    LocalMux I__2692 (
            .O(N__13803),
            .I(N__13800));
    Span4Mux_v I__2691 (
            .O(N__13800),
            .I(N__13797));
    Span4Mux_s2_v I__2690 (
            .O(N__13797),
            .I(N__13794));
    Odrv4 I__2689 (
            .O(N__13794),
            .I(\uu2.bitmapZ0Z_180 ));
    CascadeMux I__2688 (
            .O(N__13791),
            .I(N__13788));
    InMux I__2687 (
            .O(N__13788),
            .I(N__13785));
    LocalMux I__2686 (
            .O(N__13785),
            .I(N__13782));
    Odrv4 I__2685 (
            .O(N__13782),
            .I(\uu2.bitmapZ0Z_215 ));
    InMux I__2684 (
            .O(N__13779),
            .I(N__13766));
    InMux I__2683 (
            .O(N__13778),
            .I(N__13766));
    InMux I__2682 (
            .O(N__13777),
            .I(N__13766));
    InMux I__2681 (
            .O(N__13776),
            .I(N__13757));
    InMux I__2680 (
            .O(N__13775),
            .I(N__13757));
    InMux I__2679 (
            .O(N__13774),
            .I(N__13757));
    InMux I__2678 (
            .O(N__13773),
            .I(N__13757));
    LocalMux I__2677 (
            .O(N__13766),
            .I(\Lab_UT.sec1_2 ));
    LocalMux I__2676 (
            .O(N__13757),
            .I(\Lab_UT.sec1_2 ));
    InMux I__2675 (
            .O(N__13752),
            .I(N__13743));
    InMux I__2674 (
            .O(N__13751),
            .I(N__13738));
    InMux I__2673 (
            .O(N__13750),
            .I(N__13738));
    InMux I__2672 (
            .O(N__13749),
            .I(N__13729));
    InMux I__2671 (
            .O(N__13748),
            .I(N__13729));
    InMux I__2670 (
            .O(N__13747),
            .I(N__13729));
    InMux I__2669 (
            .O(N__13746),
            .I(N__13729));
    LocalMux I__2668 (
            .O(N__13743),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__2667 (
            .O(N__13738),
            .I(\Lab_UT.sec1_1 ));
    LocalMux I__2666 (
            .O(N__13729),
            .I(\Lab_UT.sec1_1 ));
    InMux I__2665 (
            .O(N__13722),
            .I(N__13709));
    InMux I__2664 (
            .O(N__13721),
            .I(N__13709));
    InMux I__2663 (
            .O(N__13720),
            .I(N__13709));
    InMux I__2662 (
            .O(N__13719),
            .I(N__13700));
    InMux I__2661 (
            .O(N__13718),
            .I(N__13700));
    InMux I__2660 (
            .O(N__13717),
            .I(N__13700));
    InMux I__2659 (
            .O(N__13716),
            .I(N__13700));
    LocalMux I__2658 (
            .O(N__13709),
            .I(N__13697));
    LocalMux I__2657 (
            .O(N__13700),
            .I(N__13694));
    Odrv4 I__2656 (
            .O(N__13697),
            .I(\Lab_UT.sec1_0 ));
    Odrv4 I__2655 (
            .O(N__13694),
            .I(\Lab_UT.sec1_0 ));
    InMux I__2654 (
            .O(N__13689),
            .I(N__13686));
    LocalMux I__2653 (
            .O(N__13686),
            .I(N__13683));
    Odrv12 I__2652 (
            .O(N__13683),
            .I(\uu2.bitmapZ0Z_212 ));
    CascadeMux I__2651 (
            .O(N__13680),
            .I(N__13675));
    CascadeMux I__2650 (
            .O(N__13679),
            .I(N__13672));
    InMux I__2649 (
            .O(N__13678),
            .I(N__13659));
    InMux I__2648 (
            .O(N__13675),
            .I(N__13659));
    InMux I__2647 (
            .O(N__13672),
            .I(N__13659));
    InMux I__2646 (
            .O(N__13671),
            .I(N__13659));
    InMux I__2645 (
            .O(N__13670),
            .I(N__13659));
    LocalMux I__2644 (
            .O(N__13659),
            .I(N__13655));
    CascadeMux I__2643 (
            .O(N__13658),
            .I(N__13651));
    Span4Mux_s0_v I__2642 (
            .O(N__13655),
            .I(N__13648));
    InMux I__2641 (
            .O(N__13654),
            .I(N__13643));
    InMux I__2640 (
            .O(N__13651),
            .I(N__13643));
    Odrv4 I__2639 (
            .O(N__13648),
            .I(\Lab_UT.min1_2 ));
    LocalMux I__2638 (
            .O(N__13643),
            .I(\Lab_UT.min1_2 ));
    InMux I__2637 (
            .O(N__13638),
            .I(N__13623));
    InMux I__2636 (
            .O(N__13637),
            .I(N__13623));
    InMux I__2635 (
            .O(N__13636),
            .I(N__13623));
    InMux I__2634 (
            .O(N__13635),
            .I(N__13623));
    InMux I__2633 (
            .O(N__13634),
            .I(N__13623));
    LocalMux I__2632 (
            .O(N__13623),
            .I(N__13618));
    InMux I__2631 (
            .O(N__13622),
            .I(N__13613));
    InMux I__2630 (
            .O(N__13621),
            .I(N__13613));
    Odrv4 I__2629 (
            .O(N__13618),
            .I(\Lab_UT.min1_0 ));
    LocalMux I__2628 (
            .O(N__13613),
            .I(\Lab_UT.min1_0 ));
    CascadeMux I__2627 (
            .O(N__13608),
            .I(N__13604));
    InMux I__2626 (
            .O(N__13607),
            .I(N__13592));
    InMux I__2625 (
            .O(N__13604),
            .I(N__13592));
    InMux I__2624 (
            .O(N__13603),
            .I(N__13592));
    InMux I__2623 (
            .O(N__13602),
            .I(N__13583));
    InMux I__2622 (
            .O(N__13601),
            .I(N__13583));
    InMux I__2621 (
            .O(N__13600),
            .I(N__13583));
    InMux I__2620 (
            .O(N__13599),
            .I(N__13583));
    LocalMux I__2619 (
            .O(N__13592),
            .I(\Lab_UT.min2_1 ));
    LocalMux I__2618 (
            .O(N__13583),
            .I(\Lab_UT.min2_1 ));
    InMux I__2617 (
            .O(N__13578),
            .I(N__13565));
    InMux I__2616 (
            .O(N__13577),
            .I(N__13565));
    InMux I__2615 (
            .O(N__13576),
            .I(N__13565));
    InMux I__2614 (
            .O(N__13575),
            .I(N__13556));
    InMux I__2613 (
            .O(N__13574),
            .I(N__13556));
    InMux I__2612 (
            .O(N__13573),
            .I(N__13556));
    InMux I__2611 (
            .O(N__13572),
            .I(N__13556));
    LocalMux I__2610 (
            .O(N__13565),
            .I(\Lab_UT.min2_0 ));
    LocalMux I__2609 (
            .O(N__13556),
            .I(\Lab_UT.min2_0 ));
    CascadeMux I__2608 (
            .O(N__13551),
            .I(N__13544));
    CascadeMux I__2607 (
            .O(N__13550),
            .I(N__13541));
    CascadeMux I__2606 (
            .O(N__13549),
            .I(N__13538));
    CascadeMux I__2605 (
            .O(N__13548),
            .I(N__13534));
    CascadeMux I__2604 (
            .O(N__13547),
            .I(N__13531));
    InMux I__2603 (
            .O(N__13544),
            .I(N__13521));
    InMux I__2602 (
            .O(N__13541),
            .I(N__13521));
    InMux I__2601 (
            .O(N__13538),
            .I(N__13521));
    InMux I__2600 (
            .O(N__13537),
            .I(N__13521));
    InMux I__2599 (
            .O(N__13534),
            .I(N__13514));
    InMux I__2598 (
            .O(N__13531),
            .I(N__13514));
    InMux I__2597 (
            .O(N__13530),
            .I(N__13514));
    LocalMux I__2596 (
            .O(N__13521),
            .I(\Lab_UT.min2_2 ));
    LocalMux I__2595 (
            .O(N__13514),
            .I(\Lab_UT.min2_2 ));
    CascadeMux I__2594 (
            .O(N__13509),
            .I(\Lab_UT.dispString.N_18_0_cascade_ ));
    InMux I__2593 (
            .O(N__13506),
            .I(N__13503));
    LocalMux I__2592 (
            .O(N__13503),
            .I(N__13500));
    Span4Mux_v I__2591 (
            .O(N__13500),
            .I(N__13497));
    Span4Mux_h I__2590 (
            .O(N__13497),
            .I(N__13494));
    Odrv4 I__2589 (
            .O(N__13494),
            .I(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ));
    InMux I__2588 (
            .O(N__13491),
            .I(N__13488));
    LocalMux I__2587 (
            .O(N__13488),
            .I(\Lab_UT.dictrl.g0_17_a6_1_7 ));
    InMux I__2586 (
            .O(N__13485),
            .I(N__13482));
    LocalMux I__2585 (
            .O(N__13482),
            .I(\Lab_UT.dictrl.g0_17_a6_1Z0Z_6 ));
    CascadeMux I__2584 (
            .O(N__13479),
            .I(\Lab_UT.dictrl.g0_17_a6_1_5_cascade_ ));
    CascadeMux I__2583 (
            .O(N__13476),
            .I(\Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_ ));
    InMux I__2582 (
            .O(N__13473),
            .I(N__13470));
    LocalMux I__2581 (
            .O(N__13470),
            .I(\Lab_UT.dictrl.g0_17_a6_2 ));
    InMux I__2580 (
            .O(N__13467),
            .I(N__13464));
    LocalMux I__2579 (
            .O(N__13464),
            .I(\Lab_UT.dictrl.N_19 ));
    InMux I__2578 (
            .O(N__13461),
            .I(N__13458));
    LocalMux I__2577 (
            .O(N__13458),
            .I(\Lab_UT.dictrl.g0_17_o6_1Z0Z_5 ));
    CascadeMux I__2576 (
            .O(N__13455),
            .I(N__13449));
    InMux I__2575 (
            .O(N__13454),
            .I(N__13440));
    InMux I__2574 (
            .O(N__13453),
            .I(N__13440));
    InMux I__2573 (
            .O(N__13452),
            .I(N__13440));
    InMux I__2572 (
            .O(N__13449),
            .I(N__13440));
    LocalMux I__2571 (
            .O(N__13440),
            .I(N__13434));
    InMux I__2570 (
            .O(N__13439),
            .I(N__13427));
    InMux I__2569 (
            .O(N__13438),
            .I(N__13427));
    InMux I__2568 (
            .O(N__13437),
            .I(N__13427));
    Odrv4 I__2567 (
            .O(N__13434),
            .I(\Lab_UT.min2_3 ));
    LocalMux I__2566 (
            .O(N__13427),
            .I(\Lab_UT.min2_3 ));
    CascadeMux I__2565 (
            .O(N__13422),
            .I(N__13416));
    CascadeMux I__2564 (
            .O(N__13421),
            .I(N__13411));
    CascadeMux I__2563 (
            .O(N__13420),
            .I(N__13408));
    CascadeMux I__2562 (
            .O(N__13419),
            .I(N__13405));
    InMux I__2561 (
            .O(N__13416),
            .I(N__13393));
    InMux I__2560 (
            .O(N__13415),
            .I(N__13393));
    InMux I__2559 (
            .O(N__13414),
            .I(N__13393));
    InMux I__2558 (
            .O(N__13411),
            .I(N__13393));
    InMux I__2557 (
            .O(N__13408),
            .I(N__13393));
    InMux I__2556 (
            .O(N__13405),
            .I(N__13388));
    InMux I__2555 (
            .O(N__13404),
            .I(N__13388));
    LocalMux I__2554 (
            .O(N__13393),
            .I(N__13385));
    LocalMux I__2553 (
            .O(N__13388),
            .I(N__13382));
    Odrv4 I__2552 (
            .O(N__13385),
            .I(\Lab_UT.min1_3 ));
    Odrv4 I__2551 (
            .O(N__13382),
            .I(\Lab_UT.min1_3 ));
    InMux I__2550 (
            .O(N__13377),
            .I(N__13374));
    LocalMux I__2549 (
            .O(N__13374),
            .I(\Lab_UT.dictrl.g1Z0Z_5 ));
    CascadeMux I__2548 (
            .O(N__13371),
            .I(\Lab_UT.dictrl.g1_cascade_ ));
    CascadeMux I__2547 (
            .O(N__13368),
            .I(\Lab_UT.dictrl.g0_2_3_cascade_ ));
    InMux I__2546 (
            .O(N__13365),
            .I(N__13361));
    InMux I__2545 (
            .O(N__13364),
            .I(N__13358));
    LocalMux I__2544 (
            .O(N__13361),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__2543 (
            .O(N__13358),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ));
    InMux I__2542 (
            .O(N__13353),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ));
    InMux I__2541 (
            .O(N__13350),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ));
    InMux I__2540 (
            .O(N__13347),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ));
    InMux I__2539 (
            .O(N__13344),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ));
    InMux I__2538 (
            .O(N__13341),
            .I(N__13331));
    InMux I__2537 (
            .O(N__13340),
            .I(N__13331));
    InMux I__2536 (
            .O(N__13339),
            .I(N__13331));
    InMux I__2535 (
            .O(N__13338),
            .I(N__13328));
    LocalMux I__2534 (
            .O(N__13331),
            .I(\buart.Z_tx.ser_clk ));
    LocalMux I__2533 (
            .O(N__13328),
            .I(\buart.Z_tx.ser_clk ));
    InMux I__2532 (
            .O(N__13323),
            .I(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ));
    CascadeMux I__2531 (
            .O(N__13320),
            .I(N__13317));
    InMux I__2530 (
            .O(N__13317),
            .I(N__13311));
    InMux I__2529 (
            .O(N__13316),
            .I(N__13311));
    LocalMux I__2528 (
            .O(N__13311),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ));
    CascadeMux I__2527 (
            .O(N__13308),
            .I(N__13305));
    InMux I__2526 (
            .O(N__13305),
            .I(N__13299));
    InMux I__2525 (
            .O(N__13304),
            .I(N__13299));
    LocalMux I__2524 (
            .O(N__13299),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ));
    CascadeMux I__2523 (
            .O(N__13296),
            .I(N__13292));
    InMux I__2522 (
            .O(N__13295),
            .I(N__13289));
    InMux I__2521 (
            .O(N__13292),
            .I(N__13286));
    LocalMux I__2520 (
            .O(N__13289),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    LocalMux I__2519 (
            .O(N__13286),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ));
    InMux I__2518 (
            .O(N__13281),
            .I(N__13275));
    InMux I__2517 (
            .O(N__13280),
            .I(N__13275));
    LocalMux I__2516 (
            .O(N__13275),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ));
    InMux I__2515 (
            .O(N__13272),
            .I(N__13269));
    LocalMux I__2514 (
            .O(N__13269),
            .I(\buart.Z_tx.Z_baudgen.ser_clk_4 ));
    InMux I__2513 (
            .O(N__13266),
            .I(N__13263));
    LocalMux I__2512 (
            .O(N__13263),
            .I(N__13260));
    Span4Mux_s2_h I__2511 (
            .O(N__13260),
            .I(N__13257));
    Span4Mux_v I__2510 (
            .O(N__13257),
            .I(N__13252));
    InMux I__2509 (
            .O(N__13256),
            .I(N__13249));
    InMux I__2508 (
            .O(N__13255),
            .I(N__13246));
    Odrv4 I__2507 (
            .O(N__13252),
            .I(L3_tx_data_1));
    LocalMux I__2506 (
            .O(N__13249),
            .I(L3_tx_data_1));
    LocalMux I__2505 (
            .O(N__13246),
            .I(L3_tx_data_1));
    InMux I__2504 (
            .O(N__13239),
            .I(N__13236));
    LocalMux I__2503 (
            .O(N__13236),
            .I(\Lab_UT.dispString.m42_ns_1 ));
    InMux I__2502 (
            .O(N__13233),
            .I(N__13230));
    LocalMux I__2501 (
            .O(N__13230),
            .I(N__13227));
    Odrv4 I__2500 (
            .O(N__13227),
            .I(vbuf_tx_data_6));
    InMux I__2499 (
            .O(N__13224),
            .I(N__13221));
    LocalMux I__2498 (
            .O(N__13221),
            .I(\buart.Z_tx.shifterZ0Z_7 ));
    CascadeMux I__2497 (
            .O(N__13218),
            .I(N__13213));
    InMux I__2496 (
            .O(N__13217),
            .I(N__13207));
    InMux I__2495 (
            .O(N__13216),
            .I(N__13207));
    InMux I__2494 (
            .O(N__13213),
            .I(N__13202));
    InMux I__2493 (
            .O(N__13212),
            .I(N__13202));
    LocalMux I__2492 (
            .O(N__13207),
            .I(N__13194));
    LocalMux I__2491 (
            .O(N__13202),
            .I(N__13194));
    InMux I__2490 (
            .O(N__13201),
            .I(N__13189));
    InMux I__2489 (
            .O(N__13200),
            .I(N__13189));
    CascadeMux I__2488 (
            .O(N__13199),
            .I(N__13177));
    Span4Mux_h I__2487 (
            .O(N__13194),
            .I(N__13172));
    LocalMux I__2486 (
            .O(N__13189),
            .I(N__13172));
    InMux I__2485 (
            .O(N__13188),
            .I(N__13155));
    InMux I__2484 (
            .O(N__13187),
            .I(N__13155));
    InMux I__2483 (
            .O(N__13186),
            .I(N__13155));
    InMux I__2482 (
            .O(N__13185),
            .I(N__13155));
    InMux I__2481 (
            .O(N__13184),
            .I(N__13155));
    InMux I__2480 (
            .O(N__13183),
            .I(N__13155));
    InMux I__2479 (
            .O(N__13182),
            .I(N__13155));
    InMux I__2478 (
            .O(N__13181),
            .I(N__13155));
    InMux I__2477 (
            .O(N__13180),
            .I(N__13152));
    InMux I__2476 (
            .O(N__13177),
            .I(N__13149));
    Span4Mux_v I__2475 (
            .O(N__13172),
            .I(N__13146));
    LocalMux I__2474 (
            .O(N__13155),
            .I(N__13141));
    LocalMux I__2473 (
            .O(N__13152),
            .I(N__13141));
    LocalMux I__2472 (
            .O(N__13149),
            .I(vbuf_tx_data_rdy));
    Odrv4 I__2471 (
            .O(N__13146),
            .I(vbuf_tx_data_rdy));
    Odrv12 I__2470 (
            .O(N__13141),
            .I(vbuf_tx_data_rdy));
    InMux I__2469 (
            .O(N__13134),
            .I(N__13131));
    LocalMux I__2468 (
            .O(N__13131),
            .I(N__13128));
    Odrv4 I__2467 (
            .O(N__13128),
            .I(vbuf_tx_data_7));
    InMux I__2466 (
            .O(N__13125),
            .I(N__13122));
    LocalMux I__2465 (
            .O(N__13122),
            .I(\buart.Z_tx.shifterZ0Z_8 ));
    CEMux I__2464 (
            .O(N__13119),
            .I(N__13116));
    LocalMux I__2463 (
            .O(N__13116),
            .I(N__13112));
    CEMux I__2462 (
            .O(N__13115),
            .I(N__13109));
    Span4Mux_v I__2461 (
            .O(N__13112),
            .I(N__13106));
    LocalMux I__2460 (
            .O(N__13109),
            .I(N__13103));
    Span4Mux_v I__2459 (
            .O(N__13106),
            .I(N__13100));
    Span4Mux_v I__2458 (
            .O(N__13103),
            .I(N__13097));
    Odrv4 I__2457 (
            .O(N__13100),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    Odrv4 I__2456 (
            .O(N__13097),
            .I(\buart.Z_tx.un1_uart_wr_i_0_i ));
    CascadeMux I__2455 (
            .O(N__13092),
            .I(N__13086));
    CascadeMux I__2454 (
            .O(N__13091),
            .I(N__13081));
    InMux I__2453 (
            .O(N__13090),
            .I(N__13075));
    InMux I__2452 (
            .O(N__13089),
            .I(N__13070));
    InMux I__2451 (
            .O(N__13086),
            .I(N__13070));
    CascadeMux I__2450 (
            .O(N__13085),
            .I(N__13065));
    InMux I__2449 (
            .O(N__13084),
            .I(N__13056));
    InMux I__2448 (
            .O(N__13081),
            .I(N__13056));
    InMux I__2447 (
            .O(N__13080),
            .I(N__13056));
    InMux I__2446 (
            .O(N__13079),
            .I(N__13056));
    CascadeMux I__2445 (
            .O(N__13078),
            .I(N__13052));
    LocalMux I__2444 (
            .O(N__13075),
            .I(N__13049));
    LocalMux I__2443 (
            .O(N__13070),
            .I(N__13046));
    InMux I__2442 (
            .O(N__13069),
            .I(N__13039));
    InMux I__2441 (
            .O(N__13068),
            .I(N__13039));
    InMux I__2440 (
            .O(N__13065),
            .I(N__13039));
    LocalMux I__2439 (
            .O(N__13056),
            .I(N__13036));
    InMux I__2438 (
            .O(N__13055),
            .I(N__13031));
    InMux I__2437 (
            .O(N__13052),
            .I(N__13031));
    Span4Mux_h I__2436 (
            .O(N__13049),
            .I(N__13026));
    Span4Mux_h I__2435 (
            .O(N__13046),
            .I(N__13026));
    LocalMux I__2434 (
            .O(N__13039),
            .I(N__13023));
    Span4Mux_h I__2433 (
            .O(N__13036),
            .I(N__13020));
    LocalMux I__2432 (
            .O(N__13031),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2431 (
            .O(N__13026),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2430 (
            .O(N__13023),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    Odrv4 I__2429 (
            .O(N__13020),
            .I(\Lab_UT.dispString.cntZ0Z_2 ));
    CascadeMux I__2428 (
            .O(N__13011),
            .I(N__13005));
    InMux I__2427 (
            .O(N__13010),
            .I(N__13002));
    InMux I__2426 (
            .O(N__13009),
            .I(N__12995));
    InMux I__2425 (
            .O(N__13008),
            .I(N__12995));
    InMux I__2424 (
            .O(N__13005),
            .I(N__12995));
    LocalMux I__2423 (
            .O(N__13002),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2422 (
            .O(N__12995),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__2421 (
            .O(N__12990),
            .I(N__12987));
    InMux I__2420 (
            .O(N__12987),
            .I(N__12982));
    InMux I__2419 (
            .O(N__12986),
            .I(N__12977));
    InMux I__2418 (
            .O(N__12985),
            .I(N__12977));
    LocalMux I__2417 (
            .O(N__12982),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__2416 (
            .O(N__12977),
            .I(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ));
    InMux I__2415 (
            .O(N__12972),
            .I(N__12968));
    CascadeMux I__2414 (
            .O(N__12971),
            .I(N__12963));
    LocalMux I__2413 (
            .O(N__12968),
            .I(N__12959));
    InMux I__2412 (
            .O(N__12967),
            .I(N__12956));
    CascadeMux I__2411 (
            .O(N__12966),
            .I(N__12953));
    InMux I__2410 (
            .O(N__12963),
            .I(N__12950));
    InMux I__2409 (
            .O(N__12962),
            .I(N__12947));
    Span4Mux_v I__2408 (
            .O(N__12959),
            .I(N__12944));
    LocalMux I__2407 (
            .O(N__12956),
            .I(N__12941));
    InMux I__2406 (
            .O(N__12953),
            .I(N__12938));
    LocalMux I__2405 (
            .O(N__12950),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__2404 (
            .O(N__12947),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__2403 (
            .O(N__12944),
            .I(\uu2.w_addr_userZ0Z_6 ));
    Odrv4 I__2402 (
            .O(N__12941),
            .I(\uu2.w_addr_userZ0Z_6 ));
    LocalMux I__2401 (
            .O(N__12938),
            .I(\uu2.w_addr_userZ0Z_6 ));
    CascadeMux I__2400 (
            .O(N__12927),
            .I(N__12922));
    InMux I__2399 (
            .O(N__12926),
            .I(N__12916));
    InMux I__2398 (
            .O(N__12925),
            .I(N__12916));
    InMux I__2397 (
            .O(N__12922),
            .I(N__12913));
    InMux I__2396 (
            .O(N__12921),
            .I(N__12908));
    LocalMux I__2395 (
            .O(N__12916),
            .I(N__12905));
    LocalMux I__2394 (
            .O(N__12913),
            .I(N__12902));
    InMux I__2393 (
            .O(N__12912),
            .I(N__12897));
    InMux I__2392 (
            .O(N__12911),
            .I(N__12897));
    LocalMux I__2391 (
            .O(N__12908),
            .I(N__12888));
    Span4Mux_h I__2390 (
            .O(N__12905),
            .I(N__12888));
    Span4Mux_v I__2389 (
            .O(N__12902),
            .I(N__12888));
    LocalMux I__2388 (
            .O(N__12897),
            .I(N__12888));
    Odrv4 I__2387 (
            .O(N__12888),
            .I(\uu2.w_addr_userZ0Z_4 ));
    CascadeMux I__2386 (
            .O(N__12885),
            .I(N__12882));
    InMux I__2385 (
            .O(N__12882),
            .I(N__12878));
    CascadeMux I__2384 (
            .O(N__12881),
            .I(N__12874));
    LocalMux I__2383 (
            .O(N__12878),
            .I(N__12870));
    InMux I__2382 (
            .O(N__12877),
            .I(N__12865));
    InMux I__2381 (
            .O(N__12874),
            .I(N__12865));
    InMux I__2380 (
            .O(N__12873),
            .I(N__12862));
    Span4Mux_s2_h I__2379 (
            .O(N__12870),
            .I(N__12857));
    LocalMux I__2378 (
            .O(N__12865),
            .I(N__12857));
    LocalMux I__2377 (
            .O(N__12862),
            .I(\uu2.N_106 ));
    Odrv4 I__2376 (
            .O(N__12857),
            .I(\uu2.N_106 ));
    CascadeMux I__2375 (
            .O(N__12852),
            .I(N__12846));
    CascadeMux I__2374 (
            .O(N__12851),
            .I(N__12843));
    InMux I__2373 (
            .O(N__12850),
            .I(N__12839));
    InMux I__2372 (
            .O(N__12849),
            .I(N__12834));
    InMux I__2371 (
            .O(N__12846),
            .I(N__12834));
    InMux I__2370 (
            .O(N__12843),
            .I(N__12829));
    InMux I__2369 (
            .O(N__12842),
            .I(N__12829));
    LocalMux I__2368 (
            .O(N__12839),
            .I(N__12826));
    LocalMux I__2367 (
            .O(N__12834),
            .I(N__12823));
    LocalMux I__2366 (
            .O(N__12829),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__2365 (
            .O(N__12826),
            .I(\uu2.w_addr_userZ0Z_5 ));
    Odrv4 I__2364 (
            .O(N__12823),
            .I(\uu2.w_addr_userZ0Z_5 ));
    CEMux I__2363 (
            .O(N__12816),
            .I(N__12812));
    CEMux I__2362 (
            .O(N__12815),
            .I(N__12809));
    LocalMux I__2361 (
            .O(N__12812),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    LocalMux I__2360 (
            .O(N__12809),
            .I(\uu2.un28_w_addr_user_i_0_0 ));
    CascadeMux I__2359 (
            .O(N__12804),
            .I(N__12801));
    InMux I__2358 (
            .O(N__12801),
            .I(N__12798));
    LocalMux I__2357 (
            .O(N__12798),
            .I(G_193));
    CascadeMux I__2356 (
            .O(N__12795),
            .I(G_193_cascade_));
    InMux I__2355 (
            .O(N__12792),
            .I(N__12789));
    LocalMux I__2354 (
            .O(N__12789),
            .I(\Lab_UT.dispString.N_219 ));
    CascadeMux I__2353 (
            .O(N__12786),
            .I(\Lab_UT.dispString.N_222_cascade_ ));
    InMux I__2352 (
            .O(N__12783),
            .I(N__12780));
    LocalMux I__2351 (
            .O(N__12780),
            .I(N__12776));
    CascadeMux I__2350 (
            .O(N__12779),
            .I(N__12773));
    Span4Mux_s2_v I__2349 (
            .O(N__12776),
            .I(N__12770));
    InMux I__2348 (
            .O(N__12773),
            .I(N__12767));
    Span4Mux_h I__2347 (
            .O(N__12770),
            .I(N__12761));
    LocalMux I__2346 (
            .O(N__12767),
            .I(N__12761));
    InMux I__2345 (
            .O(N__12766),
            .I(N__12758));
    Odrv4 I__2344 (
            .O(N__12761),
            .I(L3_tx_data_3));
    LocalMux I__2343 (
            .O(N__12758),
            .I(L3_tx_data_3));
    CascadeMux I__2342 (
            .O(N__12753),
            .I(N__12750));
    InMux I__2341 (
            .O(N__12750),
            .I(N__12747));
    LocalMux I__2340 (
            .O(N__12747),
            .I(G_189));
    CascadeMux I__2339 (
            .O(N__12744),
            .I(G_189_cascade_));
    InMux I__2338 (
            .O(N__12741),
            .I(N__12738));
    LocalMux I__2337 (
            .O(N__12738),
            .I(\Lab_UT.dispString.un42_dOutP ));
    CascadeMux I__2336 (
            .O(N__12735),
            .I(N__12732));
    InMux I__2335 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__2334 (
            .O(N__12729),
            .I(N__12726));
    Span4Mux_s2_v I__2333 (
            .O(N__12726),
            .I(N__12722));
    CascadeMux I__2332 (
            .O(N__12725),
            .I(N__12718));
    Span4Mux_h I__2331 (
            .O(N__12722),
            .I(N__12715));
    InMux I__2330 (
            .O(N__12721),
            .I(N__12712));
    InMux I__2329 (
            .O(N__12718),
            .I(N__12709));
    Odrv4 I__2328 (
            .O(N__12715),
            .I(L3_tx_data_6));
    LocalMux I__2327 (
            .O(N__12712),
            .I(L3_tx_data_6));
    LocalMux I__2326 (
            .O(N__12709),
            .I(L3_tx_data_6));
    InMux I__2325 (
            .O(N__12702),
            .I(N__12698));
    InMux I__2324 (
            .O(N__12701),
            .I(N__12695));
    LocalMux I__2323 (
            .O(N__12698),
            .I(N__12692));
    LocalMux I__2322 (
            .O(N__12695),
            .I(N__12688));
    Span4Mux_h I__2321 (
            .O(N__12692),
            .I(N__12685));
    InMux I__2320 (
            .O(N__12691),
            .I(N__12682));
    Odrv4 I__2319 (
            .O(N__12688),
            .I(uu0_sec_clkD));
    Odrv4 I__2318 (
            .O(N__12685),
            .I(uu0_sec_clkD));
    LocalMux I__2317 (
            .O(N__12682),
            .I(uu0_sec_clkD));
    InMux I__2316 (
            .O(N__12675),
            .I(N__12672));
    LocalMux I__2315 (
            .O(N__12672),
            .I(\Lab_UT.dispString.m44_ns_1 ));
    InMux I__2314 (
            .O(N__12669),
            .I(N__12657));
    InMux I__2313 (
            .O(N__12668),
            .I(N__12657));
    InMux I__2312 (
            .O(N__12667),
            .I(N__12657));
    InMux I__2311 (
            .O(N__12666),
            .I(N__12657));
    LocalMux I__2310 (
            .O(N__12657),
            .I(N__12654));
    Span4Mux_v I__2309 (
            .O(N__12654),
            .I(N__12648));
    InMux I__2308 (
            .O(N__12653),
            .I(N__12641));
    InMux I__2307 (
            .O(N__12652),
            .I(N__12641));
    InMux I__2306 (
            .O(N__12651),
            .I(N__12641));
    Odrv4 I__2305 (
            .O(N__12648),
            .I(\Lab_UT.sec2_0 ));
    LocalMux I__2304 (
            .O(N__12641),
            .I(\Lab_UT.sec2_0 ));
    InMux I__2303 (
            .O(N__12636),
            .I(N__12632));
    InMux I__2302 (
            .O(N__12635),
            .I(N__12629));
    LocalMux I__2301 (
            .O(N__12632),
            .I(G_190));
    LocalMux I__2300 (
            .O(N__12629),
            .I(G_190));
    CascadeMux I__2299 (
            .O(N__12624),
            .I(G_190_cascade_));
    InMux I__2298 (
            .O(N__12621),
            .I(N__12618));
    LocalMux I__2297 (
            .O(N__12618),
            .I(\Lab_UT.dispString.i21_mux ));
    CascadeMux I__2296 (
            .O(N__12615),
            .I(\Lab_UT.dispString.m28_ns_1_cascade_ ));
    InMux I__2295 (
            .O(N__12612),
            .I(N__12609));
    LocalMux I__2294 (
            .O(N__12609),
            .I(\Lab_UT.dispString.N_204 ));
    CascadeMux I__2293 (
            .O(N__12606),
            .I(N__12601));
    InMux I__2292 (
            .O(N__12605),
            .I(N__12596));
    InMux I__2291 (
            .O(N__12604),
            .I(N__12596));
    InMux I__2290 (
            .O(N__12601),
            .I(N__12593));
    LocalMux I__2289 (
            .O(N__12596),
            .I(\Lab_UT.di_ASones_0 ));
    LocalMux I__2288 (
            .O(N__12593),
            .I(\Lab_UT.di_ASones_0 ));
    InMux I__2287 (
            .O(N__12588),
            .I(N__12585));
    LocalMux I__2286 (
            .O(N__12585),
            .I(\uu2.bitmapZ0Z_52 ));
    CascadeMux I__2285 (
            .O(N__12582),
            .I(N__12575));
    CascadeMux I__2284 (
            .O(N__12581),
            .I(N__12572));
    InMux I__2283 (
            .O(N__12580),
            .I(N__12568));
    CascadeMux I__2282 (
            .O(N__12579),
            .I(N__12564));
    InMux I__2281 (
            .O(N__12578),
            .I(N__12561));
    InMux I__2280 (
            .O(N__12575),
            .I(N__12551));
    InMux I__2279 (
            .O(N__12572),
            .I(N__12551));
    InMux I__2278 (
            .O(N__12571),
            .I(N__12551));
    LocalMux I__2277 (
            .O(N__12568),
            .I(N__12548));
    CascadeMux I__2276 (
            .O(N__12567),
            .I(N__12544));
    InMux I__2275 (
            .O(N__12564),
            .I(N__12541));
    LocalMux I__2274 (
            .O(N__12561),
            .I(N__12538));
    InMux I__2273 (
            .O(N__12560),
            .I(N__12531));
    InMux I__2272 (
            .O(N__12559),
            .I(N__12531));
    InMux I__2271 (
            .O(N__12558),
            .I(N__12531));
    LocalMux I__2270 (
            .O(N__12551),
            .I(N__12528));
    Span4Mux_h I__2269 (
            .O(N__12548),
            .I(N__12525));
    InMux I__2268 (
            .O(N__12547),
            .I(N__12520));
    InMux I__2267 (
            .O(N__12544),
            .I(N__12520));
    LocalMux I__2266 (
            .O(N__12541),
            .I(N__12515));
    Span4Mux_h I__2265 (
            .O(N__12538),
            .I(N__12515));
    LocalMux I__2264 (
            .O(N__12531),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2263 (
            .O(N__12528),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2262 (
            .O(N__12525),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    LocalMux I__2261 (
            .O(N__12520),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    Odrv4 I__2260 (
            .O(N__12515),
            .I(\uu2.w_addr_displayingZ0Z_7 ));
    InMux I__2259 (
            .O(N__12504),
            .I(N__12501));
    LocalMux I__2258 (
            .O(N__12501),
            .I(\uu2.bitmapZ0Z_84 ));
    CascadeMux I__2257 (
            .O(N__12498),
            .I(N__12495));
    InMux I__2256 (
            .O(N__12495),
            .I(N__12492));
    LocalMux I__2255 (
            .O(N__12492),
            .I(\uu2.bitmapZ0Z_87 ));
    InMux I__2254 (
            .O(N__12489),
            .I(N__12483));
    CascadeMux I__2253 (
            .O(N__12488),
            .I(N__12480));
    InMux I__2252 (
            .O(N__12487),
            .I(N__12476));
    InMux I__2251 (
            .O(N__12486),
            .I(N__12472));
    LocalMux I__2250 (
            .O(N__12483),
            .I(N__12469));
    InMux I__2249 (
            .O(N__12480),
            .I(N__12464));
    InMux I__2248 (
            .O(N__12479),
            .I(N__12464));
    LocalMux I__2247 (
            .O(N__12476),
            .I(N__12461));
    InMux I__2246 (
            .O(N__12475),
            .I(N__12458));
    LocalMux I__2245 (
            .O(N__12472),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__2244 (
            .O(N__12469),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__2243 (
            .O(N__12464),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    Odrv4 I__2242 (
            .O(N__12461),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    LocalMux I__2241 (
            .O(N__12458),
            .I(\uu2.w_addr_displaying_fastZ0Z_0 ));
    InMux I__2240 (
            .O(N__12447),
            .I(N__12444));
    LocalMux I__2239 (
            .O(N__12444),
            .I(\uu2.bitmap_pmux_24_am_1 ));
    InMux I__2238 (
            .O(N__12441),
            .I(N__12424));
    InMux I__2237 (
            .O(N__12440),
            .I(N__12424));
    InMux I__2236 (
            .O(N__12439),
            .I(N__12424));
    InMux I__2235 (
            .O(N__12438),
            .I(N__12424));
    InMux I__2234 (
            .O(N__12437),
            .I(N__12424));
    InMux I__2233 (
            .O(N__12436),
            .I(N__12419));
    InMux I__2232 (
            .O(N__12435),
            .I(N__12419));
    LocalMux I__2231 (
            .O(N__12424),
            .I(N__12414));
    LocalMux I__2230 (
            .O(N__12419),
            .I(N__12414));
    Odrv4 I__2229 (
            .O(N__12414),
            .I(\Lab_UT.min1_1 ));
    InMux I__2228 (
            .O(N__12411),
            .I(N__12408));
    LocalMux I__2227 (
            .O(N__12408),
            .I(N__12405));
    Odrv4 I__2226 (
            .O(N__12405),
            .I(\Lab_UT.dispString.un46_dOutP_2 ));
    InMux I__2225 (
            .O(N__12402),
            .I(N__12399));
    LocalMux I__2224 (
            .O(N__12399),
            .I(\uu2.bitmap_pmux_24_bm_1 ));
    InMux I__2223 (
            .O(N__12396),
            .I(N__12393));
    LocalMux I__2222 (
            .O(N__12393),
            .I(\uu2.bitmapZ0Z_72 ));
    CascadeMux I__2221 (
            .O(N__12390),
            .I(N__12387));
    InMux I__2220 (
            .O(N__12387),
            .I(N__12384));
    LocalMux I__2219 (
            .O(N__12384),
            .I(\uu2.bitmapZ0Z_200 ));
    InMux I__2218 (
            .O(N__12381),
            .I(N__12378));
    LocalMux I__2217 (
            .O(N__12378),
            .I(N__12370));
    InMux I__2216 (
            .O(N__12377),
            .I(N__12363));
    InMux I__2215 (
            .O(N__12376),
            .I(N__12363));
    InMux I__2214 (
            .O(N__12375),
            .I(N__12363));
    InMux I__2213 (
            .O(N__12374),
            .I(N__12355));
    InMux I__2212 (
            .O(N__12373),
            .I(N__12352));
    Span4Mux_v I__2211 (
            .O(N__12370),
            .I(N__12347));
    LocalMux I__2210 (
            .O(N__12363),
            .I(N__12347));
    InMux I__2209 (
            .O(N__12362),
            .I(N__12344));
    InMux I__2208 (
            .O(N__12361),
            .I(N__12341));
    InMux I__2207 (
            .O(N__12360),
            .I(N__12338));
    InMux I__2206 (
            .O(N__12359),
            .I(N__12333));
    InMux I__2205 (
            .O(N__12358),
            .I(N__12333));
    LocalMux I__2204 (
            .O(N__12355),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2203 (
            .O(N__12352),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    Odrv4 I__2202 (
            .O(N__12347),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2201 (
            .O(N__12344),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2200 (
            .O(N__12341),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2199 (
            .O(N__12338),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    LocalMux I__2198 (
            .O(N__12333),
            .I(\uu2.w_addr_displayingZ0Z_0 ));
    InMux I__2197 (
            .O(N__12318),
            .I(N__12315));
    LocalMux I__2196 (
            .O(N__12315),
            .I(N__12312));
    Span4Mux_h I__2195 (
            .O(N__12312),
            .I(N__12309));
    Odrv4 I__2194 (
            .O(N__12309),
            .I(\uu2.bitmap_RNI5T9T1Z0Z_72 ));
    InMux I__2193 (
            .O(N__12306),
            .I(N__12303));
    LocalMux I__2192 (
            .O(N__12303),
            .I(N__12300));
    Odrv12 I__2191 (
            .O(N__12300),
            .I(\uu2.bitmap_pmux_sn_N_54_mux ));
    InMux I__2190 (
            .O(N__12297),
            .I(N__12294));
    LocalMux I__2189 (
            .O(N__12294),
            .I(\uu2.N_237 ));
    InMux I__2188 (
            .O(N__12291),
            .I(N__12288));
    LocalMux I__2187 (
            .O(N__12288),
            .I(N__12285));
    Odrv4 I__2186 (
            .O(N__12285),
            .I(\uu2.bitmap_pmux_sn_N_15 ));
    CascadeMux I__2185 (
            .O(N__12282),
            .I(\uu2.N_395_cascade_ ));
    InMux I__2184 (
            .O(N__12279),
            .I(N__12276));
    LocalMux I__2183 (
            .O(N__12276),
            .I(N__12273));
    Odrv4 I__2182 (
            .O(N__12273),
            .I(\uu2.N_401 ));
    InMux I__2181 (
            .O(N__12270),
            .I(N__12267));
    LocalMux I__2180 (
            .O(N__12267),
            .I(\uu2.bitmapZ0Z_296 ));
    InMux I__2179 (
            .O(N__12264),
            .I(N__12259));
    CascadeMux I__2178 (
            .O(N__12263),
            .I(N__12254));
    InMux I__2177 (
            .O(N__12262),
            .I(N__12249));
    LocalMux I__2176 (
            .O(N__12259),
            .I(N__12246));
    InMux I__2175 (
            .O(N__12258),
            .I(N__12243));
    InMux I__2174 (
            .O(N__12257),
            .I(N__12234));
    InMux I__2173 (
            .O(N__12254),
            .I(N__12234));
    InMux I__2172 (
            .O(N__12253),
            .I(N__12234));
    InMux I__2171 (
            .O(N__12252),
            .I(N__12234));
    LocalMux I__2170 (
            .O(N__12249),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    Odrv4 I__2169 (
            .O(N__12246),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2168 (
            .O(N__12243),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    LocalMux I__2167 (
            .O(N__12234),
            .I(\uu2.w_addr_displaying_3_repZ0Z1 ));
    CascadeMux I__2166 (
            .O(N__12225),
            .I(N__12222));
    InMux I__2165 (
            .O(N__12222),
            .I(N__12219));
    LocalMux I__2164 (
            .O(N__12219),
            .I(N__12216));
    Odrv4 I__2163 (
            .O(N__12216),
            .I(\uu2.bitmapZ0Z_40 ));
    InMux I__2162 (
            .O(N__12213),
            .I(N__12210));
    LocalMux I__2161 (
            .O(N__12210),
            .I(\uu2.bitmap_pmux_15_i_m2_ns_1 ));
    InMux I__2160 (
            .O(N__12207),
            .I(N__12204));
    LocalMux I__2159 (
            .O(N__12204),
            .I(\uu2.N_123 ));
    CascadeMux I__2158 (
            .O(N__12201),
            .I(N__12196));
    InMux I__2157 (
            .O(N__12200),
            .I(N__12187));
    InMux I__2156 (
            .O(N__12199),
            .I(N__12184));
    InMux I__2155 (
            .O(N__12196),
            .I(N__12180));
    InMux I__2154 (
            .O(N__12195),
            .I(N__12177));
    InMux I__2153 (
            .O(N__12194),
            .I(N__12168));
    InMux I__2152 (
            .O(N__12193),
            .I(N__12168));
    InMux I__2151 (
            .O(N__12192),
            .I(N__12168));
    InMux I__2150 (
            .O(N__12191),
            .I(N__12168));
    InMux I__2149 (
            .O(N__12190),
            .I(N__12165));
    LocalMux I__2148 (
            .O(N__12187),
            .I(N__12160));
    LocalMux I__2147 (
            .O(N__12184),
            .I(N__12160));
    InMux I__2146 (
            .O(N__12183),
            .I(N__12157));
    LocalMux I__2145 (
            .O(N__12180),
            .I(N__12154));
    LocalMux I__2144 (
            .O(N__12177),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2143 (
            .O(N__12168),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2142 (
            .O(N__12165),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2141 (
            .O(N__12160),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    LocalMux I__2140 (
            .O(N__12157),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    Odrv4 I__2139 (
            .O(N__12154),
            .I(\uu2.w_addr_displayingZ0Z_8 ));
    InMux I__2138 (
            .O(N__12141),
            .I(N__12138));
    LocalMux I__2137 (
            .O(N__12138),
            .I(\uu2.bitmapZ0Z_308 ));
    InMux I__2136 (
            .O(N__12135),
            .I(N__12132));
    LocalMux I__2135 (
            .O(N__12132),
            .I(\uu2.bitmap_RNIU2ISZ0Z_52 ));
    InMux I__2134 (
            .O(N__12129),
            .I(N__12126));
    LocalMux I__2133 (
            .O(N__12126),
            .I(\uu2.bitmapZ0Z_168 ));
    InMux I__2132 (
            .O(N__12123),
            .I(N__12120));
    LocalMux I__2131 (
            .O(N__12120),
            .I(\uu2.bitmapZ0Z_75 ));
    CascadeMux I__2130 (
            .O(N__12117),
            .I(N__12114));
    InMux I__2129 (
            .O(N__12114),
            .I(N__12111));
    LocalMux I__2128 (
            .O(N__12111),
            .I(\uu2.bitmapZ0Z_203 ));
    InMux I__2127 (
            .O(N__12108),
            .I(N__12105));
    LocalMux I__2126 (
            .O(N__12105),
            .I(\uu2.bitmapZ0Z_162 ));
    InMux I__2125 (
            .O(N__12102),
            .I(N__12099));
    LocalMux I__2124 (
            .O(N__12099),
            .I(\uu2.bitmapZ0Z_34 ));
    InMux I__2123 (
            .O(N__12096),
            .I(N__12092));
    InMux I__2122 (
            .O(N__12095),
            .I(N__12086));
    LocalMux I__2121 (
            .O(N__12092),
            .I(N__12083));
    InMux I__2120 (
            .O(N__12091),
            .I(N__12080));
    InMux I__2119 (
            .O(N__12090),
            .I(N__12075));
    InMux I__2118 (
            .O(N__12089),
            .I(N__12075));
    LocalMux I__2117 (
            .O(N__12086),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    Odrv4 I__2116 (
            .O(N__12083),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2115 (
            .O(N__12080),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    LocalMux I__2114 (
            .O(N__12075),
            .I(\uu2.w_addr_displaying_fastZ0Z_3 ));
    InMux I__2113 (
            .O(N__12066),
            .I(N__12063));
    LocalMux I__2112 (
            .O(N__12063),
            .I(\uu2.bitmapZ0Z_290 ));
    CascadeMux I__2111 (
            .O(N__12060),
            .I(N__12054));
    InMux I__2110 (
            .O(N__12059),
            .I(N__12048));
    InMux I__2109 (
            .O(N__12058),
            .I(N__12048));
    InMux I__2108 (
            .O(N__12057),
            .I(N__12045));
    InMux I__2107 (
            .O(N__12054),
            .I(N__12040));
    InMux I__2106 (
            .O(N__12053),
            .I(N__12040));
    LocalMux I__2105 (
            .O(N__12048),
            .I(N__12037));
    LocalMux I__2104 (
            .O(N__12045),
            .I(\buart.Z_rx.N_27_0_i ));
    LocalMux I__2103 (
            .O(N__12040),
            .I(\buart.Z_rx.N_27_0_i ));
    Odrv4 I__2102 (
            .O(N__12037),
            .I(\buart.Z_rx.N_27_0_i ));
    CEMux I__2101 (
            .O(N__12030),
            .I(N__12027));
    LocalMux I__2100 (
            .O(N__12027),
            .I(N__12022));
    CEMux I__2099 (
            .O(N__12026),
            .I(N__12019));
    CEMux I__2098 (
            .O(N__12025),
            .I(N__12016));
    Span4Mux_h I__2097 (
            .O(N__12022),
            .I(N__12011));
    LocalMux I__2096 (
            .O(N__12019),
            .I(N__12011));
    LocalMux I__2095 (
            .O(N__12016),
            .I(N__12008));
    Span4Mux_h I__2094 (
            .O(N__12011),
            .I(N__12005));
    Sp12to4 I__2093 (
            .O(N__12008),
            .I(N__12002));
    Odrv4 I__2092 (
            .O(N__12005),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    Odrv12 I__2091 (
            .O(N__12002),
            .I(\buart.Z_rx.bitcounte_0_0 ));
    InMux I__2090 (
            .O(N__11997),
            .I(N__11994));
    LocalMux I__2089 (
            .O(N__11994),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ));
    CascadeMux I__2088 (
            .O(N__11991),
            .I(N__11988));
    InMux I__2087 (
            .O(N__11988),
            .I(N__11983));
    InMux I__2086 (
            .O(N__11987),
            .I(N__11980));
    InMux I__2085 (
            .O(N__11986),
            .I(N__11977));
    LocalMux I__2084 (
            .O(N__11983),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__2083 (
            .O(N__11980),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    LocalMux I__2082 (
            .O(N__11977),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ));
    InMux I__2081 (
            .O(N__11970),
            .I(N__11966));
    InMux I__2080 (
            .O(N__11969),
            .I(N__11963));
    LocalMux I__2079 (
            .O(N__11966),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    LocalMux I__2078 (
            .O(N__11963),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ));
    CascadeMux I__2077 (
            .O(N__11958),
            .I(N__11954));
    CascadeMux I__2076 (
            .O(N__11957),
            .I(N__11951));
    InMux I__2075 (
            .O(N__11954),
            .I(N__11948));
    InMux I__2074 (
            .O(N__11951),
            .I(N__11945));
    LocalMux I__2073 (
            .O(N__11948),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    LocalMux I__2072 (
            .O(N__11945),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ));
    InMux I__2071 (
            .O(N__11940),
            .I(N__11935));
    InMux I__2070 (
            .O(N__11939),
            .I(N__11930));
    InMux I__2069 (
            .O(N__11938),
            .I(N__11930));
    LocalMux I__2068 (
            .O(N__11935),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    LocalMux I__2067 (
            .O(N__11930),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ));
    CascadeMux I__2066 (
            .O(N__11925),
            .I(N__11922));
    InMux I__2065 (
            .O(N__11922),
            .I(N__11915));
    InMux I__2064 (
            .O(N__11921),
            .I(N__11915));
    InMux I__2063 (
            .O(N__11920),
            .I(N__11912));
    LocalMux I__2062 (
            .O(N__11915),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    LocalMux I__2061 (
            .O(N__11912),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ));
    CascadeMux I__2060 (
            .O(N__11907),
            .I(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ));
    CascadeMux I__2059 (
            .O(N__11904),
            .I(N__11901));
    InMux I__2058 (
            .O(N__11901),
            .I(N__11895));
    InMux I__2057 (
            .O(N__11900),
            .I(N__11892));
    InMux I__2056 (
            .O(N__11899),
            .I(N__11887));
    InMux I__2055 (
            .O(N__11898),
            .I(N__11887));
    LocalMux I__2054 (
            .O(N__11895),
            .I(N__11884));
    LocalMux I__2053 (
            .O(N__11892),
            .I(\buart.Z_rx.ser_clk ));
    LocalMux I__2052 (
            .O(N__11887),
            .I(\buart.Z_rx.ser_clk ));
    Odrv4 I__2051 (
            .O(N__11884),
            .I(\buart.Z_rx.ser_clk ));
    InMux I__2050 (
            .O(N__11877),
            .I(N__11874));
    LocalMux I__2049 (
            .O(N__11874),
            .I(\buart.Z_rx.un1_sample_0 ));
    CascadeMux I__2048 (
            .O(N__11871),
            .I(\buart.Z_rx.ser_clk_cascade_ ));
    InMux I__2047 (
            .O(N__11868),
            .I(N__11861));
    InMux I__2046 (
            .O(N__11867),
            .I(N__11858));
    InMux I__2045 (
            .O(N__11866),
            .I(N__11851));
    InMux I__2044 (
            .O(N__11865),
            .I(N__11851));
    InMux I__2043 (
            .O(N__11864),
            .I(N__11851));
    LocalMux I__2042 (
            .O(N__11861),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2041 (
            .O(N__11858),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    LocalMux I__2040 (
            .O(N__11851),
            .I(\buart.Z_rx.bitcountZ0Z_0 ));
    IoInMux I__2039 (
            .O(N__11844),
            .I(N__11841));
    LocalMux I__2038 (
            .O(N__11841),
            .I(N__11838));
    IoSpan4Mux I__2037 (
            .O(N__11838),
            .I(N__11835));
    Span4Mux_s1_v I__2036 (
            .O(N__11835),
            .I(N__11832));
    Odrv4 I__2035 (
            .O(N__11832),
            .I(\buart.Z_rx.sample ));
    InMux I__2034 (
            .O(N__11829),
            .I(N__11814));
    InMux I__2033 (
            .O(N__11828),
            .I(N__11814));
    InMux I__2032 (
            .O(N__11827),
            .I(N__11811));
    InMux I__2031 (
            .O(N__11826),
            .I(N__11804));
    InMux I__2030 (
            .O(N__11825),
            .I(N__11804));
    InMux I__2029 (
            .O(N__11824),
            .I(N__11804));
    InMux I__2028 (
            .O(N__11823),
            .I(N__11797));
    InMux I__2027 (
            .O(N__11822),
            .I(N__11797));
    InMux I__2026 (
            .O(N__11821),
            .I(N__11797));
    InMux I__2025 (
            .O(N__11820),
            .I(N__11791));
    InMux I__2024 (
            .O(N__11819),
            .I(N__11791));
    LocalMux I__2023 (
            .O(N__11814),
            .I(N__11782));
    LocalMux I__2022 (
            .O(N__11811),
            .I(N__11782));
    LocalMux I__2021 (
            .O(N__11804),
            .I(N__11782));
    LocalMux I__2020 (
            .O(N__11797),
            .I(N__11782));
    InMux I__2019 (
            .O(N__11796),
            .I(N__11779));
    LocalMux I__2018 (
            .O(N__11791),
            .I(\buart.Z_rx.startbit ));
    Odrv4 I__2017 (
            .O(N__11782),
            .I(\buart.Z_rx.startbit ));
    LocalMux I__2016 (
            .O(N__11779),
            .I(\buart.Z_rx.startbit ));
    CascadeMux I__2015 (
            .O(N__11772),
            .I(N__11768));
    CascadeMux I__2014 (
            .O(N__11771),
            .I(N__11765));
    InMux I__2013 (
            .O(N__11768),
            .I(N__11760));
    InMux I__2012 (
            .O(N__11765),
            .I(N__11753));
    InMux I__2011 (
            .O(N__11764),
            .I(N__11753));
    InMux I__2010 (
            .O(N__11763),
            .I(N__11753));
    LocalMux I__2009 (
            .O(N__11760),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    LocalMux I__2008 (
            .O(N__11753),
            .I(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ));
    CascadeMux I__2007 (
            .O(N__11748),
            .I(\buart.Z_rx.idle_0_cascade_ ));
    InMux I__2006 (
            .O(N__11745),
            .I(N__11740));
    InMux I__2005 (
            .O(N__11744),
            .I(N__11737));
    InMux I__2004 (
            .O(N__11743),
            .I(N__11734));
    LocalMux I__2003 (
            .O(N__11740),
            .I(N__11731));
    LocalMux I__2002 (
            .O(N__11737),
            .I(\buart.Z_rx.idle ));
    LocalMux I__2001 (
            .O(N__11734),
            .I(\buart.Z_rx.idle ));
    Odrv4 I__2000 (
            .O(N__11731),
            .I(\buart.Z_rx.idle ));
    CascadeMux I__1999 (
            .O(N__11724),
            .I(N__11721));
    InMux I__1998 (
            .O(N__11721),
            .I(N__11718));
    LocalMux I__1997 (
            .O(N__11718),
            .I(N__11715));
    Odrv4 I__1996 (
            .O(N__11715),
            .I(\buart.Z_rx.bitcount_cry_2_THRU_CO ));
    CascadeMux I__1995 (
            .O(N__11712),
            .I(N__11708));
    InMux I__1994 (
            .O(N__11711),
            .I(N__11702));
    InMux I__1993 (
            .O(N__11708),
            .I(N__11699));
    InMux I__1992 (
            .O(N__11707),
            .I(N__11692));
    InMux I__1991 (
            .O(N__11706),
            .I(N__11692));
    InMux I__1990 (
            .O(N__11705),
            .I(N__11692));
    LocalMux I__1989 (
            .O(N__11702),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1988 (
            .O(N__11699),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    LocalMux I__1987 (
            .O(N__11692),
            .I(\buart.Z_rx.bitcountZ0Z_3 ));
    CascadeMux I__1986 (
            .O(N__11685),
            .I(N__11682));
    InMux I__1985 (
            .O(N__11682),
            .I(N__11675));
    InMux I__1984 (
            .O(N__11681),
            .I(N__11672));
    InMux I__1983 (
            .O(N__11680),
            .I(N__11669));
    InMux I__1982 (
            .O(N__11679),
            .I(N__11664));
    InMux I__1981 (
            .O(N__11678),
            .I(N__11664));
    LocalMux I__1980 (
            .O(N__11675),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1979 (
            .O(N__11672),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1978 (
            .O(N__11669),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    LocalMux I__1977 (
            .O(N__11664),
            .I(\buart.Z_rx.bitcountZ0Z_1 ));
    CascadeMux I__1976 (
            .O(N__11655),
            .I(N__11652));
    InMux I__1975 (
            .O(N__11652),
            .I(N__11646));
    InMux I__1974 (
            .O(N__11651),
            .I(N__11643));
    InMux I__1973 (
            .O(N__11650),
            .I(N__11638));
    InMux I__1972 (
            .O(N__11649),
            .I(N__11638));
    LocalMux I__1971 (
            .O(N__11646),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1970 (
            .O(N__11643),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    LocalMux I__1969 (
            .O(N__11638),
            .I(\buart.Z_rx.bitcountZ0Z_4 ));
    CascadeMux I__1968 (
            .O(N__11631),
            .I(\buart.Z_rx.valid_1_cascade_ ));
    InMux I__1967 (
            .O(N__11628),
            .I(N__11621));
    InMux I__1966 (
            .O(N__11627),
            .I(N__11618));
    InMux I__1965 (
            .O(N__11626),
            .I(N__11611));
    InMux I__1964 (
            .O(N__11625),
            .I(N__11611));
    InMux I__1963 (
            .O(N__11624),
            .I(N__11611));
    LocalMux I__1962 (
            .O(N__11621),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1961 (
            .O(N__11618),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    LocalMux I__1960 (
            .O(N__11611),
            .I(\buart.Z_rx.bitcountZ0Z_2 ));
    CascadeMux I__1959 (
            .O(N__11604),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ));
    InMux I__1958 (
            .O(N__11601),
            .I(N__11597));
    InMux I__1957 (
            .O(N__11600),
            .I(N__11594));
    LocalMux I__1956 (
            .O(N__11597),
            .I(N__11589));
    LocalMux I__1955 (
            .O(N__11594),
            .I(N__11589));
    Odrv12 I__1954 (
            .O(N__11589),
            .I(\Lab_UT.dispString.N_191 ));
    InMux I__1953 (
            .O(N__11586),
            .I(N__11583));
    LocalMux I__1952 (
            .O(N__11583),
            .I(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ));
    InMux I__1951 (
            .O(N__11580),
            .I(N__11576));
    InMux I__1950 (
            .O(N__11579),
            .I(N__11573));
    LocalMux I__1949 (
            .O(N__11576),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    LocalMux I__1948 (
            .O(N__11573),
            .I(\buart.Z_tx.bitcountZ0Z_3 ));
    InMux I__1947 (
            .O(N__11568),
            .I(N__11565));
    LocalMux I__1946 (
            .O(N__11565),
            .I(\buart.Z_tx.uart_busy_0_0 ));
    InMux I__1945 (
            .O(N__11562),
            .I(N__11559));
    LocalMux I__1944 (
            .O(N__11559),
            .I(N__11555));
    InMux I__1943 (
            .O(N__11558),
            .I(N__11552));
    Span4Mux_h I__1942 (
            .O(N__11555),
            .I(N__11549));
    LocalMux I__1941 (
            .O(N__11552),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    Odrv4 I__1940 (
            .O(N__11549),
            .I(\buart.Z_rx.hhZ0Z_0 ));
    InMux I__1939 (
            .O(N__11544),
            .I(N__11533));
    InMux I__1938 (
            .O(N__11543),
            .I(N__11533));
    InMux I__1937 (
            .O(N__11542),
            .I(N__11533));
    InMux I__1936 (
            .O(N__11541),
            .I(N__11528));
    InMux I__1935 (
            .O(N__11540),
            .I(N__11528));
    LocalMux I__1934 (
            .O(N__11533),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    LocalMux I__1933 (
            .O(N__11528),
            .I(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ));
    CascadeMux I__1932 (
            .O(N__11523),
            .I(N__11520));
    InMux I__1931 (
            .O(N__11520),
            .I(N__11511));
    InMux I__1930 (
            .O(N__11519),
            .I(N__11511));
    InMux I__1929 (
            .O(N__11518),
            .I(N__11504));
    InMux I__1928 (
            .O(N__11517),
            .I(N__11504));
    InMux I__1927 (
            .O(N__11516),
            .I(N__11504));
    LocalMux I__1926 (
            .O(N__11511),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    LocalMux I__1925 (
            .O(N__11504),
            .I(\buart.Z_tx.bitcountZ0Z_0 ));
    CascadeMux I__1924 (
            .O(N__11499),
            .I(N__11495));
    CascadeMux I__1923 (
            .O(N__11498),
            .I(N__11491));
    InMux I__1922 (
            .O(N__11495),
            .I(N__11484));
    InMux I__1921 (
            .O(N__11494),
            .I(N__11484));
    InMux I__1920 (
            .O(N__11491),
            .I(N__11484));
    LocalMux I__1919 (
            .O(N__11484),
            .I(\buart.Z_tx.bitcountZ0Z_2 ));
    CascadeMux I__1918 (
            .O(N__11481),
            .I(N__11476));
    InMux I__1917 (
            .O(N__11480),
            .I(N__11472));
    InMux I__1916 (
            .O(N__11479),
            .I(N__11467));
    InMux I__1915 (
            .O(N__11476),
            .I(N__11467));
    InMux I__1914 (
            .O(N__11475),
            .I(N__11464));
    LocalMux I__1913 (
            .O(N__11472),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__1912 (
            .O(N__11467),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    LocalMux I__1911 (
            .O(N__11464),
            .I(\buart.Z_tx.bitcountZ0Z_1 ));
    InMux I__1910 (
            .O(N__11457),
            .I(N__11454));
    LocalMux I__1909 (
            .O(N__11454),
            .I(\buart.Z_tx.un1_bitcount_c3 ));
    InMux I__1908 (
            .O(N__11451),
            .I(N__11448));
    LocalMux I__1907 (
            .O(N__11448),
            .I(vbuf_tx_data_0));
    InMux I__1906 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__1905 (
            .O(N__11442),
            .I(\buart.Z_tx.shifterZ0Z_1 ));
    InMux I__1904 (
            .O(N__11439),
            .I(N__11436));
    LocalMux I__1903 (
            .O(N__11436),
            .I(\buart.Z_tx.shifterZ0Z_0 ));
    IoInMux I__1902 (
            .O(N__11433),
            .I(N__11430));
    LocalMux I__1901 (
            .O(N__11430),
            .I(N__11427));
    Span4Mux_s3_h I__1900 (
            .O(N__11427),
            .I(N__11424));
    Span4Mux_v I__1899 (
            .O(N__11424),
            .I(N__11421));
    Odrv4 I__1898 (
            .O(N__11421),
            .I(o_serial_data_c));
    InMux I__1897 (
            .O(N__11418),
            .I(N__11415));
    LocalMux I__1896 (
            .O(N__11415),
            .I(vbuf_tx_data_1));
    InMux I__1895 (
            .O(N__11412),
            .I(N__11409));
    LocalMux I__1894 (
            .O(N__11409),
            .I(\buart.Z_tx.shifterZ0Z_2 ));
    InMux I__1893 (
            .O(N__11406),
            .I(N__11403));
    LocalMux I__1892 (
            .O(N__11403),
            .I(vbuf_tx_data_2));
    InMux I__1891 (
            .O(N__11400),
            .I(N__11397));
    LocalMux I__1890 (
            .O(N__11397),
            .I(\buart.Z_tx.shifterZ0Z_3 ));
    InMux I__1889 (
            .O(N__11394),
            .I(N__11391));
    LocalMux I__1888 (
            .O(N__11391),
            .I(vbuf_tx_data_3));
    InMux I__1887 (
            .O(N__11388),
            .I(N__11385));
    LocalMux I__1886 (
            .O(N__11385),
            .I(\buart.Z_tx.shifterZ0Z_4 ));
    InMux I__1885 (
            .O(N__11382),
            .I(N__11379));
    LocalMux I__1884 (
            .O(N__11379),
            .I(vbuf_tx_data_4));
    InMux I__1883 (
            .O(N__11376),
            .I(N__11373));
    LocalMux I__1882 (
            .O(N__11373),
            .I(\buart.Z_tx.shifterZ0Z_5 ));
    InMux I__1881 (
            .O(N__11370),
            .I(N__11367));
    LocalMux I__1880 (
            .O(N__11367),
            .I(vbuf_tx_data_5));
    InMux I__1879 (
            .O(N__11364),
            .I(N__11361));
    LocalMux I__1878 (
            .O(N__11361),
            .I(\buart.Z_tx.shifterZ0Z_6 ));
    CascadeMux I__1877 (
            .O(N__11358),
            .I(\Lab_UT.dispString.N_211_cascade_ ));
    InMux I__1876 (
            .O(N__11355),
            .I(N__11352));
    LocalMux I__1875 (
            .O(N__11352),
            .I(\Lab_UT.dispString.dOutP_0_iv_0_2 ));
    InMux I__1874 (
            .O(N__11349),
            .I(N__11346));
    LocalMux I__1873 (
            .O(N__11346),
            .I(\Lab_UT.dispString.dOutP_0_iv_1_2 ));
    CEMux I__1872 (
            .O(N__11343),
            .I(N__11340));
    LocalMux I__1871 (
            .O(N__11340),
            .I(N__11337));
    Span4Mux_h I__1870 (
            .O(N__11337),
            .I(N__11334));
    Odrv4 I__1869 (
            .O(N__11334),
            .I(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ));
    CascadeMux I__1868 (
            .O(N__11331),
            .I(N__11328));
    InMux I__1867 (
            .O(N__11328),
            .I(N__11325));
    LocalMux I__1866 (
            .O(N__11325),
            .I(N__11322));
    Span4Mux_h I__1865 (
            .O(N__11322),
            .I(N__11317));
    InMux I__1864 (
            .O(N__11321),
            .I(N__11314));
    InMux I__1863 (
            .O(N__11320),
            .I(N__11311));
    Odrv4 I__1862 (
            .O(N__11317),
            .I(L3_tx_data_4));
    LocalMux I__1861 (
            .O(N__11314),
            .I(L3_tx_data_4));
    LocalMux I__1860 (
            .O(N__11311),
            .I(L3_tx_data_4));
    InMux I__1859 (
            .O(N__11304),
            .I(N__11299));
    InMux I__1858 (
            .O(N__11303),
            .I(N__11296));
    InMux I__1857 (
            .O(N__11302),
            .I(N__11293));
    LocalMux I__1856 (
            .O(N__11299),
            .I(L3_tx_data_2));
    LocalMux I__1855 (
            .O(N__11296),
            .I(L3_tx_data_2));
    LocalMux I__1854 (
            .O(N__11293),
            .I(L3_tx_data_2));
    CascadeMux I__1853 (
            .O(N__11286),
            .I(\uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_ ));
    InMux I__1852 (
            .O(N__11283),
            .I(N__11280));
    LocalMux I__1851 (
            .O(N__11280),
            .I(N__11277));
    Span4Mux_h I__1850 (
            .O(N__11277),
            .I(N__11272));
    InMux I__1849 (
            .O(N__11276),
            .I(N__11269));
    InMux I__1848 (
            .O(N__11275),
            .I(N__11266));
    Odrv4 I__1847 (
            .O(N__11272),
            .I(L3_tx_data_0));
    LocalMux I__1846 (
            .O(N__11269),
            .I(L3_tx_data_0));
    LocalMux I__1845 (
            .O(N__11266),
            .I(L3_tx_data_0));
    InMux I__1844 (
            .O(N__11259),
            .I(N__11241));
    InMux I__1843 (
            .O(N__11258),
            .I(N__11241));
    InMux I__1842 (
            .O(N__11257),
            .I(N__11241));
    InMux I__1841 (
            .O(N__11256),
            .I(N__11241));
    InMux I__1840 (
            .O(N__11255),
            .I(N__11236));
    InMux I__1839 (
            .O(N__11254),
            .I(N__11236));
    CascadeMux I__1838 (
            .O(N__11253),
            .I(N__11233));
    InMux I__1837 (
            .O(N__11252),
            .I(N__11230));
    InMux I__1836 (
            .O(N__11251),
            .I(N__11225));
    InMux I__1835 (
            .O(N__11250),
            .I(N__11225));
    LocalMux I__1834 (
            .O(N__11241),
            .I(N__11220));
    LocalMux I__1833 (
            .O(N__11236),
            .I(N__11220));
    InMux I__1832 (
            .O(N__11233),
            .I(N__11217));
    LocalMux I__1831 (
            .O(N__11230),
            .I(N__11214));
    LocalMux I__1830 (
            .O(N__11225),
            .I(N__11211));
    Span4Mux_s2_h I__1829 (
            .O(N__11220),
            .I(N__11208));
    LocalMux I__1828 (
            .O(N__11217),
            .I(N__11200));
    Span4Mux_h I__1827 (
            .O(N__11214),
            .I(N__11197));
    Span4Mux_h I__1826 (
            .O(N__11211),
            .I(N__11194));
    Span4Mux_v I__1825 (
            .O(N__11208),
            .I(N__11191));
    InMux I__1824 (
            .O(N__11207),
            .I(N__11186));
    InMux I__1823 (
            .O(N__11206),
            .I(N__11186));
    InMux I__1822 (
            .O(N__11205),
            .I(N__11179));
    InMux I__1821 (
            .O(N__11204),
            .I(N__11179));
    InMux I__1820 (
            .O(N__11203),
            .I(N__11179));
    Odrv12 I__1819 (
            .O(N__11200),
            .I(\uu2.un1_w_user_cr_0 ));
    Odrv4 I__1818 (
            .O(N__11197),
            .I(\uu2.un1_w_user_cr_0 ));
    Odrv4 I__1817 (
            .O(N__11194),
            .I(\uu2.un1_w_user_cr_0 ));
    Odrv4 I__1816 (
            .O(N__11191),
            .I(\uu2.un1_w_user_cr_0 ));
    LocalMux I__1815 (
            .O(N__11186),
            .I(\uu2.un1_w_user_cr_0 ));
    LocalMux I__1814 (
            .O(N__11179),
            .I(\uu2.un1_w_user_cr_0 ));
    CascadeMux I__1813 (
            .O(N__11166),
            .I(N__11163));
    InMux I__1812 (
            .O(N__11163),
            .I(N__11160));
    LocalMux I__1811 (
            .O(N__11160),
            .I(N__11157));
    Span12Mux_s6_v I__1810 (
            .O(N__11157),
            .I(N__11152));
    InMux I__1809 (
            .O(N__11156),
            .I(N__11149));
    InMux I__1808 (
            .O(N__11155),
            .I(N__11146));
    Odrv12 I__1807 (
            .O(N__11152),
            .I(L3_tx_data_5));
    LocalMux I__1806 (
            .O(N__11149),
            .I(L3_tx_data_5));
    LocalMux I__1805 (
            .O(N__11146),
            .I(L3_tx_data_5));
    CascadeMux I__1804 (
            .O(N__11139),
            .I(\Lab_UT.didp.countrce1.q_5_0_cascade_ ));
    CascadeMux I__1803 (
            .O(N__11136),
            .I(N__11133));
    InMux I__1802 (
            .O(N__11133),
            .I(N__11121));
    InMux I__1801 (
            .O(N__11132),
            .I(N__11121));
    InMux I__1800 (
            .O(N__11131),
            .I(N__11121));
    InMux I__1799 (
            .O(N__11130),
            .I(N__11121));
    LocalMux I__1798 (
            .O(N__11121),
            .I(N__11115));
    InMux I__1797 (
            .O(N__11120),
            .I(N__11108));
    InMux I__1796 (
            .O(N__11119),
            .I(N__11108));
    InMux I__1795 (
            .O(N__11118),
            .I(N__11108));
    Odrv4 I__1794 (
            .O(N__11115),
            .I(\Lab_UT.sec2_1 ));
    LocalMux I__1793 (
            .O(N__11108),
            .I(\Lab_UT.sec2_1 ));
    InMux I__1792 (
            .O(N__11103),
            .I(N__11091));
    InMux I__1791 (
            .O(N__11102),
            .I(N__11091));
    InMux I__1790 (
            .O(N__11101),
            .I(N__11091));
    InMux I__1789 (
            .O(N__11100),
            .I(N__11091));
    LocalMux I__1788 (
            .O(N__11091),
            .I(N__11086));
    CascadeMux I__1787 (
            .O(N__11090),
            .I(N__11083));
    CascadeMux I__1786 (
            .O(N__11089),
            .I(N__11080));
    Span4Mux_h I__1785 (
            .O(N__11086),
            .I(N__11076));
    InMux I__1784 (
            .O(N__11083),
            .I(N__11069));
    InMux I__1783 (
            .O(N__11080),
            .I(N__11069));
    InMux I__1782 (
            .O(N__11079),
            .I(N__11069));
    Odrv4 I__1781 (
            .O(N__11076),
            .I(\Lab_UT.sec2_2 ));
    LocalMux I__1780 (
            .O(N__11069),
            .I(\Lab_UT.sec2_2 ));
    CascadeMux I__1779 (
            .O(N__11064),
            .I(N__11057));
    CascadeMux I__1778 (
            .O(N__11063),
            .I(N__11054));
    CascadeMux I__1777 (
            .O(N__11062),
            .I(N__11051));
    CascadeMux I__1776 (
            .O(N__11061),
            .I(N__11046));
    InMux I__1775 (
            .O(N__11060),
            .I(N__11037));
    InMux I__1774 (
            .O(N__11057),
            .I(N__11037));
    InMux I__1773 (
            .O(N__11054),
            .I(N__11037));
    InMux I__1772 (
            .O(N__11051),
            .I(N__11037));
    InMux I__1771 (
            .O(N__11050),
            .I(N__11030));
    InMux I__1770 (
            .O(N__11049),
            .I(N__11030));
    InMux I__1769 (
            .O(N__11046),
            .I(N__11030));
    LocalMux I__1768 (
            .O(N__11037),
            .I(N__11027));
    LocalMux I__1767 (
            .O(N__11030),
            .I(N__11024));
    Odrv4 I__1766 (
            .O(N__11027),
            .I(\Lab_UT.sec2_3 ));
    Odrv4 I__1765 (
            .O(N__11024),
            .I(\Lab_UT.sec2_3 ));
    CascadeMux I__1764 (
            .O(N__11019),
            .I(N__11016));
    InMux I__1763 (
            .O(N__11016),
            .I(N__11013));
    LocalMux I__1762 (
            .O(N__11013),
            .I(\uu2.un28_w_addr_user_i_0_a2_0Z0Z_4 ));
    CascadeMux I__1761 (
            .O(N__11010),
            .I(\Lab_UT.dispString.un42_dOutP_cascade_ ));
    InMux I__1760 (
            .O(N__11007),
            .I(N__11004));
    LocalMux I__1759 (
            .O(N__11004),
            .I(\uu2.un28_w_addr_user_i_0_a2_0Z0Z_0 ));
    CascadeMux I__1758 (
            .O(N__11001),
            .I(N__10998));
    InMux I__1757 (
            .O(N__10998),
            .I(N__10995));
    LocalMux I__1756 (
            .O(N__10995),
            .I(\uu2.bitmapZ0Z_218 ));
    InMux I__1755 (
            .O(N__10992),
            .I(N__10989));
    LocalMux I__1754 (
            .O(N__10989),
            .I(\uu2.bitmapZ0Z_90 ));
    InMux I__1753 (
            .O(N__10986),
            .I(N__10983));
    LocalMux I__1752 (
            .O(N__10983),
            .I(\uu2.bitmap_pmux_25_i_m2_bm_1 ));
    InMux I__1751 (
            .O(N__10980),
            .I(N__10974));
    InMux I__1750 (
            .O(N__10979),
            .I(N__10971));
    InMux I__1749 (
            .O(N__10978),
            .I(N__10965));
    InMux I__1748 (
            .O(N__10977),
            .I(N__10965));
    LocalMux I__1747 (
            .O(N__10974),
            .I(N__10960));
    LocalMux I__1746 (
            .O(N__10971),
            .I(N__10960));
    InMux I__1745 (
            .O(N__10970),
            .I(N__10957));
    LocalMux I__1744 (
            .O(N__10965),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    Odrv4 I__1743 (
            .O(N__10960),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    LocalMux I__1742 (
            .O(N__10957),
            .I(\uu2.w_addr_displaying_fastZ0Z_7 ));
    CascadeMux I__1741 (
            .O(N__10950),
            .I(\uu2.bitmap_pmux_21_ns_1_cascade_ ));
    InMux I__1740 (
            .O(N__10947),
            .I(N__10944));
    LocalMux I__1739 (
            .O(N__10944),
            .I(N__10941));
    Span4Mux_h I__1738 (
            .O(N__10941),
            .I(N__10938));
    Odrv4 I__1737 (
            .O(N__10938),
            .I(\uu2.bitmap_pmux_sn_N_11 ));
    CascadeMux I__1736 (
            .O(N__10935),
            .I(\uu2.N_393_cascade_ ));
    InMux I__1735 (
            .O(N__10932),
            .I(N__10929));
    LocalMux I__1734 (
            .O(N__10929),
            .I(\uu2.N_397 ));
    InMux I__1733 (
            .O(N__10926),
            .I(N__10920));
    InMux I__1732 (
            .O(N__10925),
            .I(N__10920));
    LocalMux I__1731 (
            .O(N__10920),
            .I(\uu2.bitmapZ0Z_314 ));
    InMux I__1730 (
            .O(N__10917),
            .I(N__10914));
    LocalMux I__1729 (
            .O(N__10914),
            .I(\uu2.N_128 ));
    InMux I__1728 (
            .O(N__10911),
            .I(N__10908));
    LocalMux I__1727 (
            .O(N__10908),
            .I(\uu2.N_131 ));
    InMux I__1726 (
            .O(N__10905),
            .I(N__10902));
    LocalMux I__1725 (
            .O(N__10902),
            .I(N__10899));
    Span4Mux_h I__1724 (
            .O(N__10899),
            .I(N__10895));
    InMux I__1723 (
            .O(N__10898),
            .I(N__10892));
    Span4Mux_v I__1722 (
            .O(N__10895),
            .I(N__10887));
    LocalMux I__1721 (
            .O(N__10892),
            .I(N__10887));
    Odrv4 I__1720 (
            .O(N__10887),
            .I(\uu2.un1_l_count_1_0 ));
    InMux I__1719 (
            .O(N__10884),
            .I(N__10881));
    LocalMux I__1718 (
            .O(N__10881),
            .I(\uu2.bitmap_RNIFJI02Z0Z_212 ));
    InMux I__1717 (
            .O(N__10878),
            .I(N__10871));
    InMux I__1716 (
            .O(N__10877),
            .I(N__10871));
    InMux I__1715 (
            .O(N__10876),
            .I(N__10868));
    LocalMux I__1714 (
            .O(N__10871),
            .I(N__10865));
    LocalMux I__1713 (
            .O(N__10868),
            .I(N__10862));
    Odrv4 I__1712 (
            .O(N__10865),
            .I(\uu2.N_65 ));
    Odrv4 I__1711 (
            .O(N__10862),
            .I(\uu2.N_65 ));
    InMux I__1710 (
            .O(N__10857),
            .I(N__10854));
    LocalMux I__1709 (
            .O(N__10854),
            .I(N__10851));
    Odrv12 I__1708 (
            .O(N__10851),
            .I(\uu2.bitmap_pmux_u_0_83_0 ));
    InMux I__1707 (
            .O(N__10848),
            .I(N__10832));
    InMux I__1706 (
            .O(N__10847),
            .I(N__10832));
    InMux I__1705 (
            .O(N__10846),
            .I(N__10832));
    InMux I__1704 (
            .O(N__10845),
            .I(N__10832));
    InMux I__1703 (
            .O(N__10844),
            .I(N__10832));
    InMux I__1702 (
            .O(N__10843),
            .I(N__10824));
    LocalMux I__1701 (
            .O(N__10832),
            .I(N__10821));
    InMux I__1700 (
            .O(N__10831),
            .I(N__10818));
    InMux I__1699 (
            .O(N__10830),
            .I(N__10809));
    InMux I__1698 (
            .O(N__10829),
            .I(N__10809));
    InMux I__1697 (
            .O(N__10828),
            .I(N__10809));
    InMux I__1696 (
            .O(N__10827),
            .I(N__10809));
    LocalMux I__1695 (
            .O(N__10824),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    Odrv4 I__1694 (
            .O(N__10821),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__1693 (
            .O(N__10818),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    LocalMux I__1692 (
            .O(N__10809),
            .I(\uu2.w_addr_displayingZ0Z_5 ));
    CascadeMux I__1691 (
            .O(N__10800),
            .I(N__10794));
    CascadeMux I__1690 (
            .O(N__10799),
            .I(N__10790));
    CascadeMux I__1689 (
            .O(N__10798),
            .I(N__10784));
    InMux I__1688 (
            .O(N__10797),
            .I(N__10780));
    InMux I__1687 (
            .O(N__10794),
            .I(N__10771));
    InMux I__1686 (
            .O(N__10793),
            .I(N__10771));
    InMux I__1685 (
            .O(N__10790),
            .I(N__10771));
    InMux I__1684 (
            .O(N__10789),
            .I(N__10771));
    InMux I__1683 (
            .O(N__10788),
            .I(N__10764));
    InMux I__1682 (
            .O(N__10787),
            .I(N__10764));
    InMux I__1681 (
            .O(N__10784),
            .I(N__10764));
    InMux I__1680 (
            .O(N__10783),
            .I(N__10761));
    LocalMux I__1679 (
            .O(N__10780),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__1678 (
            .O(N__10771),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__1677 (
            .O(N__10764),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    LocalMux I__1676 (
            .O(N__10761),
            .I(\uu2.w_addr_displayingZ0Z_6 ));
    InMux I__1675 (
            .O(N__10752),
            .I(N__10749));
    LocalMux I__1674 (
            .O(N__10749),
            .I(\uu2.bitmap_pmux_sn_N_42 ));
    InMux I__1673 (
            .O(N__10746),
            .I(N__10743));
    LocalMux I__1672 (
            .O(N__10743),
            .I(\uu2.N_112_i ));
    CascadeMux I__1671 (
            .O(N__10740),
            .I(\uu2.N_100_cascade_ ));
    InMux I__1670 (
            .O(N__10737),
            .I(N__10734));
    LocalMux I__1669 (
            .O(N__10734),
            .I(\uu2.N_921_tz_tz ));
    InMux I__1668 (
            .O(N__10731),
            .I(N__10728));
    LocalMux I__1667 (
            .O(N__10728),
            .I(N__10725));
    Odrv4 I__1666 (
            .O(N__10725),
            .I(\uu2.bitmap_pmux_sn_N_20 ));
    CascadeMux I__1665 (
            .O(N__10722),
            .I(\uu2.N_923_tz_cascade_ ));
    InMux I__1664 (
            .O(N__10719),
            .I(N__10716));
    LocalMux I__1663 (
            .O(N__10716),
            .I(N__10713));
    Odrv4 I__1662 (
            .O(N__10713),
            .I(\uu2.w_addr_displaying_RNI8ND5GZ0Z_3 ));
    CascadeMux I__1661 (
            .O(N__10710),
            .I(N__10707));
    InMux I__1660 (
            .O(N__10707),
            .I(N__10701));
    InMux I__1659 (
            .O(N__10706),
            .I(N__10701));
    LocalMux I__1658 (
            .O(N__10701),
            .I(N__10692));
    InMux I__1657 (
            .O(N__10700),
            .I(N__10687));
    InMux I__1656 (
            .O(N__10699),
            .I(N__10687));
    InMux I__1655 (
            .O(N__10698),
            .I(N__10675));
    InMux I__1654 (
            .O(N__10697),
            .I(N__10675));
    InMux I__1653 (
            .O(N__10696),
            .I(N__10675));
    InMux I__1652 (
            .O(N__10695),
            .I(N__10675));
    Span12Mux_s4_h I__1651 (
            .O(N__10692),
            .I(N__10672));
    LocalMux I__1650 (
            .O(N__10687),
            .I(N__10669));
    InMux I__1649 (
            .O(N__10686),
            .I(N__10662));
    InMux I__1648 (
            .O(N__10685),
            .I(N__10662));
    InMux I__1647 (
            .O(N__10684),
            .I(N__10662));
    LocalMux I__1646 (
            .O(N__10675),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__1645 (
            .O(N__10672),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    Odrv12 I__1644 (
            .O(N__10669),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    LocalMux I__1643 (
            .O(N__10662),
            .I(\uu2.w_addr_displayingZ0Z_2 ));
    CascadeMux I__1642 (
            .O(N__10653),
            .I(N__10650));
    InMux I__1641 (
            .O(N__10650),
            .I(N__10645));
    CascadeMux I__1640 (
            .O(N__10649),
            .I(N__10642));
    CascadeMux I__1639 (
            .O(N__10648),
            .I(N__10639));
    LocalMux I__1638 (
            .O(N__10645),
            .I(N__10633));
    InMux I__1637 (
            .O(N__10642),
            .I(N__10624));
    InMux I__1636 (
            .O(N__10639),
            .I(N__10624));
    InMux I__1635 (
            .O(N__10638),
            .I(N__10624));
    InMux I__1634 (
            .O(N__10637),
            .I(N__10624));
    InMux I__1633 (
            .O(N__10636),
            .I(N__10621));
    Span4Mux_s1_v I__1632 (
            .O(N__10633),
            .I(N__10618));
    LocalMux I__1631 (
            .O(N__10624),
            .I(N__10615));
    LocalMux I__1630 (
            .O(N__10621),
            .I(N__10612));
    Odrv4 I__1629 (
            .O(N__10618),
            .I(\uu2.N_34 ));
    Odrv4 I__1628 (
            .O(N__10615),
            .I(\uu2.N_34 ));
    Odrv12 I__1627 (
            .O(N__10612),
            .I(\uu2.N_34 ));
    InMux I__1626 (
            .O(N__10605),
            .I(N__10601));
    CascadeMux I__1625 (
            .O(N__10604),
            .I(N__10597));
    LocalMux I__1624 (
            .O(N__10601),
            .I(N__10592));
    InMux I__1623 (
            .O(N__10600),
            .I(N__10587));
    InMux I__1622 (
            .O(N__10597),
            .I(N__10587));
    CascadeMux I__1621 (
            .O(N__10596),
            .I(N__10583));
    InMux I__1620 (
            .O(N__10595),
            .I(N__10580));
    Span4Mux_v I__1619 (
            .O(N__10592),
            .I(N__10574));
    LocalMux I__1618 (
            .O(N__10587),
            .I(N__10574));
    InMux I__1617 (
            .O(N__10586),
            .I(N__10569));
    InMux I__1616 (
            .O(N__10583),
            .I(N__10566));
    LocalMux I__1615 (
            .O(N__10580),
            .I(N__10563));
    InMux I__1614 (
            .O(N__10579),
            .I(N__10560));
    Span4Mux_h I__1613 (
            .O(N__10574),
            .I(N__10557));
    InMux I__1612 (
            .O(N__10573),
            .I(N__10552));
    InMux I__1611 (
            .O(N__10572),
            .I(N__10552));
    LocalMux I__1610 (
            .O(N__10569),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__1609 (
            .O(N__10566),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__1608 (
            .O(N__10563),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__1607 (
            .O(N__10560),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    Odrv4 I__1606 (
            .O(N__10557),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    LocalMux I__1605 (
            .O(N__10552),
            .I(\uu2.w_addr_displayingZ0Z_3 ));
    InMux I__1604 (
            .O(N__10539),
            .I(N__10536));
    LocalMux I__1603 (
            .O(N__10536),
            .I(N__10533));
    Span4Mux_h I__1602 (
            .O(N__10533),
            .I(N__10530));
    Odrv4 I__1601 (
            .O(N__10530),
            .I(\uu2.N_47 ));
    CascadeMux I__1600 (
            .O(N__10527),
            .I(N__10521));
    CascadeMux I__1599 (
            .O(N__10526),
            .I(N__10518));
    CascadeMux I__1598 (
            .O(N__10525),
            .I(N__10514));
    InMux I__1597 (
            .O(N__10524),
            .I(N__10502));
    InMux I__1596 (
            .O(N__10521),
            .I(N__10502));
    InMux I__1595 (
            .O(N__10518),
            .I(N__10502));
    InMux I__1594 (
            .O(N__10517),
            .I(N__10502));
    InMux I__1593 (
            .O(N__10514),
            .I(N__10502));
    InMux I__1592 (
            .O(N__10513),
            .I(N__10499));
    LocalMux I__1591 (
            .O(N__10502),
            .I(N__10496));
    LocalMux I__1590 (
            .O(N__10499),
            .I(N__10493));
    Span4Mux_h I__1589 (
            .O(N__10496),
            .I(N__10490));
    Odrv12 I__1588 (
            .O(N__10493),
            .I(\uu2.N_38 ));
    Odrv4 I__1587 (
            .O(N__10490),
            .I(\uu2.N_38 ));
    InMux I__1586 (
            .O(N__10485),
            .I(N__10473));
    InMux I__1585 (
            .O(N__10484),
            .I(N__10456));
    InMux I__1584 (
            .O(N__10483),
            .I(N__10456));
    InMux I__1583 (
            .O(N__10482),
            .I(N__10456));
    InMux I__1582 (
            .O(N__10481),
            .I(N__10456));
    InMux I__1581 (
            .O(N__10480),
            .I(N__10456));
    InMux I__1580 (
            .O(N__10479),
            .I(N__10456));
    InMux I__1579 (
            .O(N__10478),
            .I(N__10456));
    InMux I__1578 (
            .O(N__10477),
            .I(N__10456));
    InMux I__1577 (
            .O(N__10476),
            .I(N__10453));
    LocalMux I__1576 (
            .O(N__10473),
            .I(N__10448));
    LocalMux I__1575 (
            .O(N__10456),
            .I(N__10448));
    LocalMux I__1574 (
            .O(N__10453),
            .I(N__10445));
    Span4Mux_s1_v I__1573 (
            .O(N__10448),
            .I(N__10442));
    Odrv12 I__1572 (
            .O(N__10445),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_5 ));
    Odrv4 I__1571 (
            .O(N__10442),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_5 ));
    InMux I__1570 (
            .O(N__10437),
            .I(N__10428));
    InMux I__1569 (
            .O(N__10436),
            .I(N__10428));
    InMux I__1568 (
            .O(N__10435),
            .I(N__10428));
    LocalMux I__1567 (
            .O(N__10428),
            .I(N__10422));
    InMux I__1566 (
            .O(N__10427),
            .I(N__10417));
    InMux I__1565 (
            .O(N__10426),
            .I(N__10417));
    InMux I__1564 (
            .O(N__10425),
            .I(N__10414));
    Span4Mux_s3_h I__1563 (
            .O(N__10422),
            .I(N__10409));
    LocalMux I__1562 (
            .O(N__10417),
            .I(N__10409));
    LocalMux I__1561 (
            .O(N__10414),
            .I(\uu2.N_33 ));
    Odrv4 I__1560 (
            .O(N__10409),
            .I(\uu2.N_33 ));
    InMux I__1559 (
            .O(N__10404),
            .I(N__10392));
    InMux I__1558 (
            .O(N__10403),
            .I(N__10392));
    InMux I__1557 (
            .O(N__10402),
            .I(N__10392));
    InMux I__1556 (
            .O(N__10401),
            .I(N__10384));
    InMux I__1555 (
            .O(N__10400),
            .I(N__10384));
    InMux I__1554 (
            .O(N__10399),
            .I(N__10384));
    LocalMux I__1553 (
            .O(N__10392),
            .I(N__10381));
    InMux I__1552 (
            .O(N__10391),
            .I(N__10371));
    LocalMux I__1551 (
            .O(N__10384),
            .I(N__10368));
    Span4Mux_h I__1550 (
            .O(N__10381),
            .I(N__10365));
    InMux I__1549 (
            .O(N__10380),
            .I(N__10362));
    InMux I__1548 (
            .O(N__10379),
            .I(N__10357));
    InMux I__1547 (
            .O(N__10378),
            .I(N__10357));
    InMux I__1546 (
            .O(N__10377),
            .I(N__10348));
    InMux I__1545 (
            .O(N__10376),
            .I(N__10348));
    InMux I__1544 (
            .O(N__10375),
            .I(N__10348));
    InMux I__1543 (
            .O(N__10374),
            .I(N__10348));
    LocalMux I__1542 (
            .O(N__10371),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1541 (
            .O(N__10368),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    Odrv4 I__1540 (
            .O(N__10365),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1539 (
            .O(N__10362),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1538 (
            .O(N__10357),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    LocalMux I__1537 (
            .O(N__10348),
            .I(\uu2.w_addr_displayingZ0Z_1 ));
    CascadeMux I__1536 (
            .O(N__10335),
            .I(N__10325));
    CascadeMux I__1535 (
            .O(N__10334),
            .I(N__10321));
    CascadeMux I__1534 (
            .O(N__10333),
            .I(N__10318));
    InMux I__1533 (
            .O(N__10332),
            .I(N__10313));
    InMux I__1532 (
            .O(N__10331),
            .I(N__10310));
    InMux I__1531 (
            .O(N__10330),
            .I(N__10303));
    InMux I__1530 (
            .O(N__10329),
            .I(N__10303));
    InMux I__1529 (
            .O(N__10328),
            .I(N__10303));
    InMux I__1528 (
            .O(N__10325),
            .I(N__10298));
    InMux I__1527 (
            .O(N__10324),
            .I(N__10298));
    InMux I__1526 (
            .O(N__10321),
            .I(N__10294));
    InMux I__1525 (
            .O(N__10318),
            .I(N__10291));
    InMux I__1524 (
            .O(N__10317),
            .I(N__10286));
    InMux I__1523 (
            .O(N__10316),
            .I(N__10286));
    LocalMux I__1522 (
            .O(N__10313),
            .I(N__10283));
    LocalMux I__1521 (
            .O(N__10310),
            .I(N__10276));
    LocalMux I__1520 (
            .O(N__10303),
            .I(N__10276));
    LocalMux I__1519 (
            .O(N__10298),
            .I(N__10276));
    InMux I__1518 (
            .O(N__10297),
            .I(N__10270));
    LocalMux I__1517 (
            .O(N__10294),
            .I(N__10265));
    LocalMux I__1516 (
            .O(N__10291),
            .I(N__10265));
    LocalMux I__1515 (
            .O(N__10286),
            .I(N__10258));
    Span4Mux_h I__1514 (
            .O(N__10283),
            .I(N__10258));
    Span4Mux_s3_h I__1513 (
            .O(N__10276),
            .I(N__10258));
    InMux I__1512 (
            .O(N__10275),
            .I(N__10255));
    InMux I__1511 (
            .O(N__10274),
            .I(N__10250));
    InMux I__1510 (
            .O(N__10273),
            .I(N__10250));
    LocalMux I__1509 (
            .O(N__10270),
            .I(L3_tx_data_rdy));
    Odrv12 I__1508 (
            .O(N__10265),
            .I(L3_tx_data_rdy));
    Odrv4 I__1507 (
            .O(N__10258),
            .I(L3_tx_data_rdy));
    LocalMux I__1506 (
            .O(N__10255),
            .I(L3_tx_data_rdy));
    LocalMux I__1505 (
            .O(N__10250),
            .I(L3_tx_data_rdy));
    CascadeMux I__1504 (
            .O(N__10239),
            .I(N__10236));
    InMux I__1503 (
            .O(N__10236),
            .I(N__10233));
    LocalMux I__1502 (
            .O(N__10233),
            .I(N__10230));
    Odrv4 I__1501 (
            .O(N__10230),
            .I(\uu2.mem0.N_136 ));
    InMux I__1500 (
            .O(N__10227),
            .I(N__10224));
    LocalMux I__1499 (
            .O(N__10224),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ));
    InMux I__1498 (
            .O(N__10221),
            .I(N__10218));
    LocalMux I__1497 (
            .O(N__10218),
            .I(\uu2.bitmapZ0Z_194 ));
    CascadeMux I__1496 (
            .O(N__10215),
            .I(\uu2.bitmap_pmux_25_i_m2_am_1_cascade_ ));
    InMux I__1495 (
            .O(N__10212),
            .I(N__10209));
    LocalMux I__1494 (
            .O(N__10209),
            .I(N__10206));
    Odrv4 I__1493 (
            .O(N__10206),
            .I(\uu2.bitmap_RNIG91I1Z0Z_66 ));
    CascadeMux I__1492 (
            .O(N__10203),
            .I(N__10200));
    InMux I__1491 (
            .O(N__10200),
            .I(N__10197));
    LocalMux I__1490 (
            .O(N__10197),
            .I(\uu2.bitmapZ0Z_69 ));
    InMux I__1489 (
            .O(N__10194),
            .I(N__10191));
    LocalMux I__1488 (
            .O(N__10191),
            .I(\uu2.bitmapZ0Z_66 ));
    InMux I__1487 (
            .O(N__10188),
            .I(N__10185));
    LocalMux I__1486 (
            .O(N__10185),
            .I(\uu2.bitmapZ0Z_197 ));
    InMux I__1485 (
            .O(N__10182),
            .I(N__10179));
    LocalMux I__1484 (
            .O(N__10179),
            .I(\buart.Z_rx.bitcount_cry_0_THRU_CO ));
    InMux I__1483 (
            .O(N__10176),
            .I(\buart.Z_rx.bitcount_cry_0 ));
    InMux I__1482 (
            .O(N__10173),
            .I(N__10170));
    LocalMux I__1481 (
            .O(N__10170),
            .I(\buart.Z_rx.bitcount_cry_1_THRU_CO ));
    InMux I__1480 (
            .O(N__10167),
            .I(\buart.Z_rx.bitcount_cry_1 ));
    InMux I__1479 (
            .O(N__10164),
            .I(\buart.Z_rx.bitcount_cry_2 ));
    InMux I__1478 (
            .O(N__10161),
            .I(\buart.Z_rx.bitcount_cry_3 ));
    InMux I__1477 (
            .O(N__10158),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ));
    InMux I__1476 (
            .O(N__10155),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ));
    InMux I__1475 (
            .O(N__10152),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ));
    InMux I__1474 (
            .O(N__10149),
            .I(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ));
    InMux I__1473 (
            .O(N__10146),
            .I(N__10143));
    LocalMux I__1472 (
            .O(N__10143),
            .I(N__10140));
    Odrv4 I__1471 (
            .O(N__10140),
            .I(\uu2.trig_rd_detZ0Z_1 ));
    InMux I__1470 (
            .O(N__10137),
            .I(N__10133));
    InMux I__1469 (
            .O(N__10136),
            .I(N__10130));
    LocalMux I__1468 (
            .O(N__10133),
            .I(N__10127));
    LocalMux I__1467 (
            .O(N__10130),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    Odrv4 I__1466 (
            .O(N__10127),
            .I(\uu2.trig_rd_detZ0Z_0 ));
    CascadeMux I__1465 (
            .O(N__10122),
            .I(N__10118));
    InMux I__1464 (
            .O(N__10121),
            .I(N__10111));
    InMux I__1463 (
            .O(N__10118),
            .I(N__10108));
    InMux I__1462 (
            .O(N__10117),
            .I(N__10103));
    InMux I__1461 (
            .O(N__10116),
            .I(N__10103));
    InMux I__1460 (
            .O(N__10115),
            .I(N__10098));
    InMux I__1459 (
            .O(N__10114),
            .I(N__10098));
    LocalMux I__1458 (
            .O(N__10111),
            .I(N__10095));
    LocalMux I__1457 (
            .O(N__10108),
            .I(N__10092));
    LocalMux I__1456 (
            .O(N__10103),
            .I(N__10089));
    LocalMux I__1455 (
            .O(N__10098),
            .I(N__10086));
    Span4Mux_s3_h I__1454 (
            .O(N__10095),
            .I(N__10083));
    Span4Mux_s2_h I__1453 (
            .O(N__10092),
            .I(N__10080));
    Span12Mux_s3_h I__1452 (
            .O(N__10089),
            .I(N__10077));
    Span4Mux_s3_h I__1451 (
            .O(N__10086),
            .I(N__10074));
    Span4Mux_v I__1450 (
            .O(N__10083),
            .I(N__10071));
    Odrv4 I__1449 (
            .O(N__10080),
            .I(\uu2.trig_rd_is_det ));
    Odrv12 I__1448 (
            .O(N__10077),
            .I(\uu2.trig_rd_is_det ));
    Odrv4 I__1447 (
            .O(N__10074),
            .I(\uu2.trig_rd_is_det ));
    Odrv4 I__1446 (
            .O(N__10071),
            .I(\uu2.trig_rd_is_det ));
    InMux I__1445 (
            .O(N__10062),
            .I(N__10058));
    InMux I__1444 (
            .O(N__10061),
            .I(N__10055));
    LocalMux I__1443 (
            .O(N__10058),
            .I(N__10052));
    LocalMux I__1442 (
            .O(N__10055),
            .I(N__10046));
    Span4Mux_v I__1441 (
            .O(N__10052),
            .I(N__10043));
    InMux I__1440 (
            .O(N__10051),
            .I(N__10036));
    InMux I__1439 (
            .O(N__10050),
            .I(N__10036));
    InMux I__1438 (
            .O(N__10049),
            .I(N__10036));
    Odrv4 I__1437 (
            .O(N__10046),
            .I(\uu2.l_countZ0Z_4 ));
    Odrv4 I__1436 (
            .O(N__10043),
            .I(\uu2.l_countZ0Z_4 ));
    LocalMux I__1435 (
            .O(N__10036),
            .I(\uu2.l_countZ0Z_4 ));
    InMux I__1434 (
            .O(N__10029),
            .I(N__10024));
    InMux I__1433 (
            .O(N__10028),
            .I(N__10021));
    InMux I__1432 (
            .O(N__10027),
            .I(N__10018));
    LocalMux I__1431 (
            .O(N__10024),
            .I(N__10015));
    LocalMux I__1430 (
            .O(N__10021),
            .I(N__10012));
    LocalMux I__1429 (
            .O(N__10018),
            .I(\uu2.l_countZ0Z_5 ));
    Odrv4 I__1428 (
            .O(N__10015),
            .I(\uu2.l_countZ0Z_5 ));
    Odrv4 I__1427 (
            .O(N__10012),
            .I(\uu2.l_countZ0Z_5 ));
    InMux I__1426 (
            .O(N__10005),
            .I(N__9998));
    InMux I__1425 (
            .O(N__10004),
            .I(N__9998));
    InMux I__1424 (
            .O(N__10003),
            .I(N__9995));
    LocalMux I__1423 (
            .O(N__9998),
            .I(N__9992));
    LocalMux I__1422 (
            .O(N__9995),
            .I(N__9989));
    Span4Mux_s3_h I__1421 (
            .O(N__9992),
            .I(N__9986));
    Odrv4 I__1420 (
            .O(N__9989),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    Odrv4 I__1419 (
            .O(N__9986),
            .I(\uu2.vbuf_count.un328_ci_3 ));
    InMux I__1418 (
            .O(N__9981),
            .I(N__9978));
    LocalMux I__1417 (
            .O(N__9978),
            .I(N__9975));
    Span4Mux_v I__1416 (
            .O(N__9975),
            .I(N__9972));
    Odrv4 I__1415 (
            .O(N__9972),
            .I(\uu2.mem0.N_54_i ));
    InMux I__1414 (
            .O(N__9969),
            .I(N__9966));
    LocalMux I__1413 (
            .O(N__9966),
            .I(N__9963));
    Span4Mux_v I__1412 (
            .O(N__9963),
            .I(N__9960));
    Odrv4 I__1411 (
            .O(N__9960),
            .I(\uu2.r_data_wire_0 ));
    InMux I__1410 (
            .O(N__9957),
            .I(N__9954));
    LocalMux I__1409 (
            .O(N__9954),
            .I(N__9951));
    Span4Mux_v I__1408 (
            .O(N__9951),
            .I(N__9948));
    Odrv4 I__1407 (
            .O(N__9948),
            .I(\uu2.r_data_wire_1 ));
    InMux I__1406 (
            .O(N__9945),
            .I(N__9942));
    LocalMux I__1405 (
            .O(N__9942),
            .I(N__9939));
    Span4Mux_v I__1404 (
            .O(N__9939),
            .I(N__9936));
    Odrv4 I__1403 (
            .O(N__9936),
            .I(\uu2.r_data_wire_2 ));
    InMux I__1402 (
            .O(N__9933),
            .I(N__9930));
    LocalMux I__1401 (
            .O(N__9930),
            .I(N__9927));
    Span4Mux_v I__1400 (
            .O(N__9927),
            .I(N__9924));
    Odrv4 I__1399 (
            .O(N__9924),
            .I(\uu2.r_data_wire_3 ));
    InMux I__1398 (
            .O(N__9921),
            .I(N__9918));
    LocalMux I__1397 (
            .O(N__9918),
            .I(N__9915));
    Span4Mux_v I__1396 (
            .O(N__9915),
            .I(N__9912));
    Odrv4 I__1395 (
            .O(N__9912),
            .I(\uu2.r_data_wire_4 ));
    InMux I__1394 (
            .O(N__9909),
            .I(N__9906));
    LocalMux I__1393 (
            .O(N__9906),
            .I(N__9903));
    Span4Mux_v I__1392 (
            .O(N__9903),
            .I(N__9900));
    Odrv4 I__1391 (
            .O(N__9900),
            .I(\uu2.r_data_wire_5 ));
    InMux I__1390 (
            .O(N__9897),
            .I(N__9894));
    LocalMux I__1389 (
            .O(N__9894),
            .I(N__9891));
    Span4Mux_v I__1388 (
            .O(N__9891),
            .I(N__9888));
    Odrv4 I__1387 (
            .O(N__9888),
            .I(\uu2.r_data_wire_6 ));
    InMux I__1386 (
            .O(N__9885),
            .I(N__9882));
    LocalMux I__1385 (
            .O(N__9882),
            .I(N__9879));
    Span4Mux_v I__1384 (
            .O(N__9879),
            .I(N__9876));
    Odrv4 I__1383 (
            .O(N__9876),
            .I(\uu2.r_data_wire_7 ));
    CascadeMux I__1382 (
            .O(N__9873),
            .I(\uu2.N_106_cascade_ ));
    CascadeMux I__1381 (
            .O(N__9870),
            .I(N__9867));
    InMux I__1380 (
            .O(N__9867),
            .I(N__9864));
    LocalMux I__1379 (
            .O(N__9864),
            .I(N__9861));
    Odrv4 I__1378 (
            .O(N__9861),
            .I(\uu2.N_164 ));
    InMux I__1377 (
            .O(N__9858),
            .I(N__9854));
    CascadeMux I__1376 (
            .O(N__9857),
            .I(N__9851));
    LocalMux I__1375 (
            .O(N__9854),
            .I(N__9847));
    InMux I__1374 (
            .O(N__9851),
            .I(N__9840));
    InMux I__1373 (
            .O(N__9850),
            .I(N__9840));
    Span4Mux_v I__1372 (
            .O(N__9847),
            .I(N__9837));
    InMux I__1371 (
            .O(N__9846),
            .I(N__9832));
    InMux I__1370 (
            .O(N__9845),
            .I(N__9832));
    LocalMux I__1369 (
            .O(N__9840),
            .I(\uu2.w_addr_userZ0Z_2 ));
    Odrv4 I__1368 (
            .O(N__9837),
            .I(\uu2.w_addr_userZ0Z_2 ));
    LocalMux I__1367 (
            .O(N__9832),
            .I(\uu2.w_addr_userZ0Z_2 ));
    InMux I__1366 (
            .O(N__9825),
            .I(N__9822));
    LocalMux I__1365 (
            .O(N__9822),
            .I(\uu2.w_addr_user_3_i_a2_3_6 ));
    CascadeMux I__1364 (
            .O(N__9819),
            .I(\uu2.w_addr_user_3_i_a2_2_6_cascade_ ));
    InMux I__1363 (
            .O(N__9816),
            .I(N__9811));
    InMux I__1362 (
            .O(N__9815),
            .I(N__9808));
    InMux I__1361 (
            .O(N__9814),
            .I(N__9805));
    LocalMux I__1360 (
            .O(N__9811),
            .I(\uu2.N_230 ));
    LocalMux I__1359 (
            .O(N__9808),
            .I(\uu2.N_230 ));
    LocalMux I__1358 (
            .O(N__9805),
            .I(\uu2.N_230 ));
    InMux I__1357 (
            .O(N__9798),
            .I(N__9792));
    InMux I__1356 (
            .O(N__9797),
            .I(N__9789));
    InMux I__1355 (
            .O(N__9796),
            .I(N__9784));
    InMux I__1354 (
            .O(N__9795),
            .I(N__9784));
    LocalMux I__1353 (
            .O(N__9792),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1352 (
            .O(N__9789),
            .I(\uu2.w_addr_userZ0Z_3 ));
    LocalMux I__1351 (
            .O(N__9784),
            .I(\uu2.w_addr_userZ0Z_3 ));
    CascadeMux I__1350 (
            .O(N__9777),
            .I(N__9774));
    InMux I__1349 (
            .O(N__9774),
            .I(N__9771));
    LocalMux I__1348 (
            .O(N__9771),
            .I(N__9768));
    Span4Mux_s3_h I__1347 (
            .O(N__9768),
            .I(N__9765));
    Odrv4 I__1346 (
            .O(N__9765),
            .I(\uu2.mem0.N_138 ));
    CascadeMux I__1345 (
            .O(N__9762),
            .I(oneSecStrb_cascade_));
    IoInMux I__1344 (
            .O(N__9759),
            .I(N__9755));
    InMux I__1343 (
            .O(N__9758),
            .I(N__9752));
    LocalMux I__1342 (
            .O(N__9755),
            .I(N__9749));
    LocalMux I__1341 (
            .O(N__9752),
            .I(N__9746));
    Span12Mux_s9_v I__1340 (
            .O(N__9749),
            .I(N__9741));
    Span12Mux_s5_h I__1339 (
            .O(N__9746),
            .I(N__9741));
    Odrv12 I__1338 (
            .O(N__9741),
            .I(clk));
    SRMux I__1337 (
            .O(N__9738),
            .I(N__9734));
    CEMux I__1336 (
            .O(N__9737),
            .I(N__9731));
    LocalMux I__1335 (
            .O(N__9734),
            .I(N__9728));
    LocalMux I__1334 (
            .O(N__9731),
            .I(N__9725));
    Span4Mux_h I__1333 (
            .O(N__9728),
            .I(N__9720));
    Span4Mux_h I__1332 (
            .O(N__9725),
            .I(N__9720));
    Odrv4 I__1331 (
            .O(N__9720),
            .I(\uu2.vram_wr_en_0_iZ0 ));
    CascadeMux I__1330 (
            .O(N__9717),
            .I(N__9711));
    InMux I__1329 (
            .O(N__9716),
            .I(N__9706));
    InMux I__1328 (
            .O(N__9715),
            .I(N__9701));
    InMux I__1327 (
            .O(N__9714),
            .I(N__9701));
    InMux I__1326 (
            .O(N__9711),
            .I(N__9694));
    InMux I__1325 (
            .O(N__9710),
            .I(N__9694));
    InMux I__1324 (
            .O(N__9709),
            .I(N__9694));
    LocalMux I__1323 (
            .O(N__9706),
            .I(N__9691));
    LocalMux I__1322 (
            .O(N__9701),
            .I(N__9686));
    LocalMux I__1321 (
            .O(N__9694),
            .I(N__9686));
    Span4Mux_s3_h I__1320 (
            .O(N__9691),
            .I(N__9682));
    Span4Mux_h I__1319 (
            .O(N__9686),
            .I(N__9679));
    InMux I__1318 (
            .O(N__9685),
            .I(N__9676));
    Span4Mux_v I__1317 (
            .O(N__9682),
            .I(N__9673));
    Span4Mux_s2_v I__1316 (
            .O(N__9679),
            .I(N__9668));
    LocalMux I__1315 (
            .O(N__9676),
            .I(N__9668));
    Odrv4 I__1314 (
            .O(N__9673),
            .I(\uu2.N_102 ));
    Odrv4 I__1313 (
            .O(N__9668),
            .I(\uu2.N_102 ));
    CascadeMux I__1312 (
            .O(N__9663),
            .I(N__9658));
    InMux I__1311 (
            .O(N__9662),
            .I(N__9655));
    InMux I__1310 (
            .O(N__9661),
            .I(N__9650));
    InMux I__1309 (
            .O(N__9658),
            .I(N__9650));
    LocalMux I__1308 (
            .O(N__9655),
            .I(\uu2.w_addr_userZ0Z_8 ));
    LocalMux I__1307 (
            .O(N__9650),
            .I(\uu2.w_addr_userZ0Z_8 ));
    CascadeMux I__1306 (
            .O(N__9645),
            .I(\uu2.N_161_cascade_ ));
    CascadeMux I__1305 (
            .O(N__9642),
            .I(\uu2.N_101_cascade_ ));
    CascadeMux I__1304 (
            .O(N__9639),
            .I(N__9633));
    CascadeMux I__1303 (
            .O(N__9638),
            .I(N__9628));
    CascadeMux I__1302 (
            .O(N__9637),
            .I(N__9625));
    InMux I__1301 (
            .O(N__9636),
            .I(N__9618));
    InMux I__1300 (
            .O(N__9633),
            .I(N__9618));
    InMux I__1299 (
            .O(N__9632),
            .I(N__9618));
    CascadeMux I__1298 (
            .O(N__9631),
            .I(N__9615));
    InMux I__1297 (
            .O(N__9628),
            .I(N__9612));
    InMux I__1296 (
            .O(N__9625),
            .I(N__9609));
    LocalMux I__1295 (
            .O(N__9618),
            .I(N__9606));
    InMux I__1294 (
            .O(N__9615),
            .I(N__9603));
    LocalMux I__1293 (
            .O(N__9612),
            .I(N__9600));
    LocalMux I__1292 (
            .O(N__9609),
            .I(N__9597));
    Span4Mux_h I__1291 (
            .O(N__9606),
            .I(N__9594));
    LocalMux I__1290 (
            .O(N__9603),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv12 I__1289 (
            .O(N__9600),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv12 I__1288 (
            .O(N__9597),
            .I(\uu2.w_addr_userZ0Z_1 ));
    Odrv4 I__1287 (
            .O(N__9594),
            .I(\uu2.w_addr_userZ0Z_1 ));
    CascadeMux I__1286 (
            .O(N__9585),
            .I(N__9581));
    InMux I__1285 (
            .O(N__9584),
            .I(N__9578));
    InMux I__1284 (
            .O(N__9581),
            .I(N__9575));
    LocalMux I__1283 (
            .O(N__9578),
            .I(N__9571));
    LocalMux I__1282 (
            .O(N__9575),
            .I(N__9568));
    InMux I__1281 (
            .O(N__9574),
            .I(N__9561));
    Span4Mux_v I__1280 (
            .O(N__9571),
            .I(N__9556));
    Span4Mux_v I__1279 (
            .O(N__9568),
            .I(N__9556));
    InMux I__1278 (
            .O(N__9567),
            .I(N__9547));
    InMux I__1277 (
            .O(N__9566),
            .I(N__9547));
    InMux I__1276 (
            .O(N__9565),
            .I(N__9547));
    InMux I__1275 (
            .O(N__9564),
            .I(N__9547));
    LocalMux I__1274 (
            .O(N__9561),
            .I(\uu2.w_addr_userZ0Z_0 ));
    Odrv4 I__1273 (
            .O(N__9556),
            .I(\uu2.w_addr_userZ0Z_0 ));
    LocalMux I__1272 (
            .O(N__9547),
            .I(\uu2.w_addr_userZ0Z_0 ));
    CascadeMux I__1271 (
            .O(N__9540),
            .I(N__9537));
    InMux I__1270 (
            .O(N__9537),
            .I(N__9534));
    LocalMux I__1269 (
            .O(N__9534),
            .I(N__9531));
    Odrv4 I__1268 (
            .O(N__9531),
            .I(\uu2.mem0.N_135 ));
    CascadeMux I__1267 (
            .O(N__9528),
            .I(N__9525));
    InMux I__1266 (
            .O(N__9525),
            .I(N__9522));
    LocalMux I__1265 (
            .O(N__9522),
            .I(\uu2.mem0.N_134 ));
    CascadeMux I__1264 (
            .O(N__9519),
            .I(\uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_ ));
    CEMux I__1263 (
            .O(N__9516),
            .I(N__9512));
    CEMux I__1262 (
            .O(N__9515),
            .I(N__9509));
    LocalMux I__1261 (
            .O(N__9512),
            .I(N__9506));
    LocalMux I__1260 (
            .O(N__9509),
            .I(N__9503));
    Span4Mux_h I__1259 (
            .O(N__9506),
            .I(N__9500));
    Span4Mux_s0_v I__1258 (
            .O(N__9503),
            .I(N__9497));
    Span4Mux_s0_h I__1257 (
            .O(N__9500),
            .I(N__9494));
    Odrv4 I__1256 (
            .O(N__9497),
            .I(\uu2.N_32_0 ));
    Odrv4 I__1255 (
            .O(N__9494),
            .I(\uu2.N_32_0 ));
    CascadeMux I__1254 (
            .O(N__9489),
            .I(N__9486));
    InMux I__1253 (
            .O(N__9486),
            .I(N__9483));
    LocalMux I__1252 (
            .O(N__9483),
            .I(N__9480));
    Odrv4 I__1251 (
            .O(N__9480),
            .I(\uu2.mem0.N_133 ));
    CascadeMux I__1250 (
            .O(N__9477),
            .I(N__9471));
    InMux I__1249 (
            .O(N__9476),
            .I(N__9459));
    InMux I__1248 (
            .O(N__9475),
            .I(N__9459));
    InMux I__1247 (
            .O(N__9474),
            .I(N__9459));
    InMux I__1246 (
            .O(N__9471),
            .I(N__9459));
    InMux I__1245 (
            .O(N__9470),
            .I(N__9459));
    LocalMux I__1244 (
            .O(N__9459),
            .I(\uu2.w_addr_displaying_fastZ0Z_2 ));
    InMux I__1243 (
            .O(N__9456),
            .I(N__9453));
    LocalMux I__1242 (
            .O(N__9453),
            .I(\uu2.bitmapZ0Z_186 ));
    InMux I__1241 (
            .O(N__9450),
            .I(N__9447));
    LocalMux I__1240 (
            .O(N__9447),
            .I(\uu2.bitmapZ0Z_58 ));
    InMux I__1239 (
            .O(N__9444),
            .I(N__9441));
    LocalMux I__1238 (
            .O(N__9441),
            .I(\uu2.bitmapZ0Z_93 ));
    CascadeMux I__1237 (
            .O(N__9438),
            .I(N__9435));
    InMux I__1236 (
            .O(N__9435),
            .I(N__9432));
    LocalMux I__1235 (
            .O(N__9432),
            .I(\uu2.bitmapZ0Z_221 ));
    CascadeMux I__1234 (
            .O(N__9429),
            .I(\uu2.bitmap_RNIRETJ1Z0Z_93_cascade_ ));
    CascadeMux I__1233 (
            .O(N__9426),
            .I(\uu2.bitmap_pmux_27_ns_1_cascade_ ));
    CascadeMux I__1232 (
            .O(N__9423),
            .I(N__9420));
    InMux I__1231 (
            .O(N__9420),
            .I(N__9417));
    LocalMux I__1230 (
            .O(N__9417),
            .I(N__9414));
    Odrv4 I__1229 (
            .O(N__9414),
            .I(\uu2.N_404 ));
    InMux I__1228 (
            .O(N__9411),
            .I(N__9408));
    LocalMux I__1227 (
            .O(N__9408),
            .I(N__9405));
    Span4Mux_s3_h I__1226 (
            .O(N__9405),
            .I(N__9402));
    Odrv4 I__1225 (
            .O(N__9402),
            .I(\uu2.bitmap_pmux_u_0_a2_0_2_0 ));
    InMux I__1224 (
            .O(N__9399),
            .I(N__9394));
    InMux I__1223 (
            .O(N__9398),
            .I(N__9389));
    InMux I__1222 (
            .O(N__9397),
            .I(N__9389));
    LocalMux I__1221 (
            .O(N__9394),
            .I(N__9385));
    LocalMux I__1220 (
            .O(N__9389),
            .I(N__9382));
    CascadeMux I__1219 (
            .O(N__9388),
            .I(N__9377));
    Span4Mux_v I__1218 (
            .O(N__9385),
            .I(N__9371));
    Span4Mux_s3_h I__1217 (
            .O(N__9382),
            .I(N__9368));
    InMux I__1216 (
            .O(N__9381),
            .I(N__9359));
    InMux I__1215 (
            .O(N__9380),
            .I(N__9359));
    InMux I__1214 (
            .O(N__9377),
            .I(N__9359));
    InMux I__1213 (
            .O(N__9376),
            .I(N__9359));
    InMux I__1212 (
            .O(N__9375),
            .I(N__9354));
    InMux I__1211 (
            .O(N__9374),
            .I(N__9354));
    Odrv4 I__1210 (
            .O(N__9371),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    Odrv4 I__1209 (
            .O(N__9368),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__1208 (
            .O(N__9359),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    LocalMux I__1207 (
            .O(N__9354),
            .I(\uu2.w_addr_displayingZ0Z_4 ));
    CascadeMux I__1206 (
            .O(N__9345),
            .I(\uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_ ));
    InMux I__1205 (
            .O(N__9342),
            .I(N__9335));
    InMux I__1204 (
            .O(N__9341),
            .I(N__9328));
    InMux I__1203 (
            .O(N__9340),
            .I(N__9328));
    InMux I__1202 (
            .O(N__9339),
            .I(N__9328));
    InMux I__1201 (
            .O(N__9338),
            .I(N__9325));
    LocalMux I__1200 (
            .O(N__9335),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1199 (
            .O(N__9328),
            .I(\uu2.l_countZ0Z_1 ));
    LocalMux I__1198 (
            .O(N__9325),
            .I(\uu2.l_countZ0Z_1 ));
    InMux I__1197 (
            .O(N__9318),
            .I(N__9304));
    InMux I__1196 (
            .O(N__9317),
            .I(N__9304));
    InMux I__1195 (
            .O(N__9316),
            .I(N__9304));
    InMux I__1194 (
            .O(N__9315),
            .I(N__9304));
    InMux I__1193 (
            .O(N__9314),
            .I(N__9299));
    InMux I__1192 (
            .O(N__9313),
            .I(N__9299));
    LocalMux I__1191 (
            .O(N__9304),
            .I(\uu2.l_countZ0Z_0 ));
    LocalMux I__1190 (
            .O(N__9299),
            .I(\uu2.l_countZ0Z_0 ));
    CascadeMux I__1189 (
            .O(N__9294),
            .I(N__9290));
    CascadeMux I__1188 (
            .O(N__9293),
            .I(N__9287));
    InMux I__1187 (
            .O(N__9290),
            .I(N__9283));
    InMux I__1186 (
            .O(N__9287),
            .I(N__9280));
    InMux I__1185 (
            .O(N__9286),
            .I(N__9277));
    LocalMux I__1184 (
            .O(N__9283),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__1183 (
            .O(N__9280),
            .I(\uu2.l_countZ0Z_3 ));
    LocalMux I__1182 (
            .O(N__9277),
            .I(\uu2.l_countZ0Z_3 ));
    CascadeMux I__1181 (
            .O(N__9270),
            .I(N__9264));
    InMux I__1180 (
            .O(N__9269),
            .I(N__9259));
    InMux I__1179 (
            .O(N__9268),
            .I(N__9259));
    InMux I__1178 (
            .O(N__9267),
            .I(N__9256));
    InMux I__1177 (
            .O(N__9264),
            .I(N__9253));
    LocalMux I__1176 (
            .O(N__9259),
            .I(N__9250));
    LocalMux I__1175 (
            .O(N__9256),
            .I(\uu2.un306_ci ));
    LocalMux I__1174 (
            .O(N__9253),
            .I(\uu2.un306_ci ));
    Odrv4 I__1173 (
            .O(N__9250),
            .I(\uu2.un306_ci ));
    InMux I__1172 (
            .O(N__9243),
            .I(N__9236));
    InMux I__1171 (
            .O(N__9242),
            .I(N__9236));
    InMux I__1170 (
            .O(N__9241),
            .I(N__9233));
    LocalMux I__1169 (
            .O(N__9236),
            .I(\uu2.l_countZ0Z_7 ));
    LocalMux I__1168 (
            .O(N__9233),
            .I(\uu2.l_countZ0Z_7 ));
    CascadeMux I__1167 (
            .O(N__9228),
            .I(\uu2.un306_ci_cascade_ ));
    InMux I__1166 (
            .O(N__9225),
            .I(N__9216));
    InMux I__1165 (
            .O(N__9224),
            .I(N__9216));
    InMux I__1164 (
            .O(N__9223),
            .I(N__9211));
    InMux I__1163 (
            .O(N__9222),
            .I(N__9211));
    InMux I__1162 (
            .O(N__9221),
            .I(N__9208));
    LocalMux I__1161 (
            .O(N__9216),
            .I(N__9203));
    LocalMux I__1160 (
            .O(N__9211),
            .I(N__9203));
    LocalMux I__1159 (
            .O(N__9208),
            .I(\uu2.l_countZ0Z_6 ));
    Odrv4 I__1158 (
            .O(N__9203),
            .I(\uu2.l_countZ0Z_6 ));
    InMux I__1157 (
            .O(N__9198),
            .I(N__9194));
    InMux I__1156 (
            .O(N__9197),
            .I(N__9191));
    LocalMux I__1155 (
            .O(N__9194),
            .I(\uu2.un284_ci ));
    LocalMux I__1154 (
            .O(N__9191),
            .I(\uu2.un284_ci ));
    CascadeMux I__1153 (
            .O(N__9186),
            .I(N__9181));
    InMux I__1152 (
            .O(N__9185),
            .I(N__9172));
    InMux I__1151 (
            .O(N__9184),
            .I(N__9172));
    InMux I__1150 (
            .O(N__9181),
            .I(N__9172));
    InMux I__1149 (
            .O(N__9180),
            .I(N__9169));
    InMux I__1148 (
            .O(N__9179),
            .I(N__9166));
    LocalMux I__1147 (
            .O(N__9172),
            .I(N__9163));
    LocalMux I__1146 (
            .O(N__9169),
            .I(\uu2.l_countZ0Z_2 ));
    LocalMux I__1145 (
            .O(N__9166),
            .I(\uu2.l_countZ0Z_2 ));
    Odrv4 I__1144 (
            .O(N__9163),
            .I(\uu2.l_countZ0Z_2 ));
    InMux I__1143 (
            .O(N__9156),
            .I(N__9152));
    InMux I__1142 (
            .O(N__9155),
            .I(N__9149));
    LocalMux I__1141 (
            .O(N__9152),
            .I(\uu2.un350_ci ));
    LocalMux I__1140 (
            .O(N__9149),
            .I(\uu2.un350_ci ));
    CascadeMux I__1139 (
            .O(N__9144),
            .I(N__9140));
    InMux I__1138 (
            .O(N__9143),
            .I(N__9134));
    InMux I__1137 (
            .O(N__9140),
            .I(N__9134));
    InMux I__1136 (
            .O(N__9139),
            .I(N__9131));
    LocalMux I__1135 (
            .O(N__9134),
            .I(N__9128));
    LocalMux I__1134 (
            .O(N__9131),
            .I(\uu2.l_countZ0Z_8 ));
    Odrv4 I__1133 (
            .O(N__9128),
            .I(\uu2.l_countZ0Z_8 ));
    CascadeMux I__1132 (
            .O(N__9123),
            .I(N__9119));
    CascadeMux I__1131 (
            .O(N__9122),
            .I(N__9116));
    InMux I__1130 (
            .O(N__9119),
            .I(N__9113));
    InMux I__1129 (
            .O(N__9116),
            .I(N__9110));
    LocalMux I__1128 (
            .O(N__9113),
            .I(N__9106));
    LocalMux I__1127 (
            .O(N__9110),
            .I(N__9103));
    InMux I__1126 (
            .O(N__9109),
            .I(N__9100));
    Span4Mux_v I__1125 (
            .O(N__9106),
            .I(N__9095));
    Span4Mux_h I__1124 (
            .O(N__9103),
            .I(N__9095));
    LocalMux I__1123 (
            .O(N__9100),
            .I(\uu0.un88_ci_3 ));
    Odrv4 I__1122 (
            .O(N__9095),
            .I(\uu0.un88_ci_3 ));
    InMux I__1121 (
            .O(N__9090),
            .I(N__9087));
    LocalMux I__1120 (
            .O(N__9087),
            .I(N__9081));
    InMux I__1119 (
            .O(N__9086),
            .I(N__9078));
    InMux I__1118 (
            .O(N__9085),
            .I(N__9075));
    InMux I__1117 (
            .O(N__9084),
            .I(N__9072));
    Span4Mux_v I__1116 (
            .O(N__9081),
            .I(N__9067));
    LocalMux I__1115 (
            .O(N__9078),
            .I(N__9067));
    LocalMux I__1114 (
            .O(N__9075),
            .I(N__9064));
    LocalMux I__1113 (
            .O(N__9072),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1112 (
            .O(N__9067),
            .I(\uu0.l_countZ0Z_6 ));
    Odrv4 I__1111 (
            .O(N__9064),
            .I(\uu0.l_countZ0Z_6 ));
    CascadeMux I__1110 (
            .O(N__9057),
            .I(N__9054));
    InMux I__1109 (
            .O(N__9054),
            .I(N__9051));
    LocalMux I__1108 (
            .O(N__9051),
            .I(N__9048));
    Odrv12 I__1107 (
            .O(N__9048),
            .I(\uu0.un99_ci_0 ));
    CascadeMux I__1106 (
            .O(N__9045),
            .I(\uu2.w_data_0_a2_0_6_cascade_ ));
    InMux I__1105 (
            .O(N__9042),
            .I(N__9034));
    InMux I__1104 (
            .O(N__9041),
            .I(N__9023));
    InMux I__1103 (
            .O(N__9040),
            .I(N__9023));
    InMux I__1102 (
            .O(N__9039),
            .I(N__9023));
    InMux I__1101 (
            .O(N__9038),
            .I(N__9023));
    InMux I__1100 (
            .O(N__9037),
            .I(N__9023));
    LocalMux I__1099 (
            .O(N__9034),
            .I(N__9018));
    LocalMux I__1098 (
            .O(N__9023),
            .I(N__9018));
    Span4Mux_v I__1097 (
            .O(N__9018),
            .I(N__9015));
    Odrv4 I__1096 (
            .O(N__9015),
            .I(\uu2.w_data_0_a2_2_6 ));
    CascadeMux I__1095 (
            .O(N__9012),
            .I(\uu2.un1_l_count_2_2_cascade_ ));
    CascadeMux I__1094 (
            .O(N__9009),
            .I(\uu2.un1_l_count_2_0_cascade_ ));
    InMux I__1093 (
            .O(N__9006),
            .I(N__9000));
    InMux I__1092 (
            .O(N__9005),
            .I(N__9000));
    LocalMux I__1091 (
            .O(N__9000),
            .I(\uu2.un1_l_count_1_3 ));
    InMux I__1090 (
            .O(N__8997),
            .I(N__8992));
    InMux I__1089 (
            .O(N__8996),
            .I(N__8987));
    InMux I__1088 (
            .O(N__8995),
            .I(N__8987));
    LocalMux I__1087 (
            .O(N__8992),
            .I(N__8984));
    LocalMux I__1086 (
            .O(N__8987),
            .I(\uu2.un1_l_count_2_0 ));
    Odrv4 I__1085 (
            .O(N__8984),
            .I(\uu2.un1_l_count_2_0 ));
    CascadeMux I__1084 (
            .O(N__8979),
            .I(N__8974));
    CascadeMux I__1083 (
            .O(N__8978),
            .I(N__8971));
    CascadeMux I__1082 (
            .O(N__8977),
            .I(N__8968));
    InMux I__1081 (
            .O(N__8974),
            .I(N__8961));
    InMux I__1080 (
            .O(N__8971),
            .I(N__8961));
    InMux I__1079 (
            .O(N__8968),
            .I(N__8961));
    LocalMux I__1078 (
            .O(N__8961),
            .I(\uu2.l_countZ0Z_9 ));
    InMux I__1077 (
            .O(N__8958),
            .I(N__8955));
    LocalMux I__1076 (
            .O(N__8955),
            .I(\uu2.un1_l_count_1_2_0 ));
    InMux I__1075 (
            .O(N__8952),
            .I(N__8946));
    InMux I__1074 (
            .O(N__8951),
            .I(N__8943));
    InMux I__1073 (
            .O(N__8950),
            .I(N__8940));
    InMux I__1072 (
            .O(N__8949),
            .I(N__8937));
    LocalMux I__1071 (
            .O(N__8946),
            .I(N__8933));
    LocalMux I__1070 (
            .O(N__8943),
            .I(N__8930));
    LocalMux I__1069 (
            .O(N__8940),
            .I(N__8927));
    LocalMux I__1068 (
            .O(N__8937),
            .I(N__8924));
    InMux I__1067 (
            .O(N__8936),
            .I(N__8921));
    Odrv4 I__1066 (
            .O(N__8933),
            .I(\uu0.un66_ci ));
    Odrv4 I__1065 (
            .O(N__8930),
            .I(\uu0.un66_ci ));
    Odrv12 I__1064 (
            .O(N__8927),
            .I(\uu0.un66_ci ));
    Odrv4 I__1063 (
            .O(N__8924),
            .I(\uu0.un66_ci ));
    LocalMux I__1062 (
            .O(N__8921),
            .I(\uu0.un66_ci ));
    InMux I__1061 (
            .O(N__8910),
            .I(N__8905));
    InMux I__1060 (
            .O(N__8909),
            .I(N__8900));
    InMux I__1059 (
            .O(N__8908),
            .I(N__8900));
    LocalMux I__1058 (
            .O(N__8905),
            .I(N__8893));
    LocalMux I__1057 (
            .O(N__8900),
            .I(N__8893));
    CascadeMux I__1056 (
            .O(N__8899),
            .I(N__8890));
    CascadeMux I__1055 (
            .O(N__8898),
            .I(N__8886));
    Span4Mux_v I__1054 (
            .O(N__8893),
            .I(N__8879));
    InMux I__1053 (
            .O(N__8890),
            .I(N__8876));
    InMux I__1052 (
            .O(N__8889),
            .I(N__8871));
    InMux I__1051 (
            .O(N__8886),
            .I(N__8871));
    InMux I__1050 (
            .O(N__8885),
            .I(N__8862));
    InMux I__1049 (
            .O(N__8884),
            .I(N__8862));
    InMux I__1048 (
            .O(N__8883),
            .I(N__8862));
    InMux I__1047 (
            .O(N__8882),
            .I(N__8862));
    Odrv4 I__1046 (
            .O(N__8879),
            .I(\uu0.un110_ci ));
    LocalMux I__1045 (
            .O(N__8876),
            .I(\uu0.un110_ci ));
    LocalMux I__1044 (
            .O(N__8871),
            .I(\uu0.un110_ci ));
    LocalMux I__1043 (
            .O(N__8862),
            .I(\uu0.un110_ci ));
    InMux I__1042 (
            .O(N__8853),
            .I(N__8844));
    InMux I__1041 (
            .O(N__8852),
            .I(N__8844));
    InMux I__1040 (
            .O(N__8851),
            .I(N__8844));
    LocalMux I__1039 (
            .O(N__8844),
            .I(N__8841));
    Odrv4 I__1038 (
            .O(N__8841),
            .I(\uu0.un198_ci_2 ));
    CascadeMux I__1037 (
            .O(N__8838),
            .I(\uu0.un110_ci_cascade_ ));
    InMux I__1036 (
            .O(N__8835),
            .I(N__8825));
    InMux I__1035 (
            .O(N__8834),
            .I(N__8825));
    InMux I__1034 (
            .O(N__8833),
            .I(N__8825));
    InMux I__1033 (
            .O(N__8832),
            .I(N__8822));
    LocalMux I__1032 (
            .O(N__8825),
            .I(\uu0.l_countZ0Z_16 ));
    LocalMux I__1031 (
            .O(N__8822),
            .I(\uu0.l_countZ0Z_16 ));
    CascadeMux I__1030 (
            .O(N__8817),
            .I(N__8810));
    InMux I__1029 (
            .O(N__8816),
            .I(N__8806));
    InMux I__1028 (
            .O(N__8815),
            .I(N__8797));
    InMux I__1027 (
            .O(N__8814),
            .I(N__8790));
    InMux I__1026 (
            .O(N__8813),
            .I(N__8790));
    InMux I__1025 (
            .O(N__8810),
            .I(N__8790));
    InMux I__1024 (
            .O(N__8809),
            .I(N__8787));
    LocalMux I__1023 (
            .O(N__8806),
            .I(N__8784));
    InMux I__1022 (
            .O(N__8805),
            .I(N__8777));
    InMux I__1021 (
            .O(N__8804),
            .I(N__8777));
    InMux I__1020 (
            .O(N__8803),
            .I(N__8777));
    InMux I__1019 (
            .O(N__8802),
            .I(N__8774));
    InMux I__1018 (
            .O(N__8801),
            .I(N__8771));
    InMux I__1017 (
            .O(N__8800),
            .I(N__8768));
    LocalMux I__1016 (
            .O(N__8797),
            .I(N__8763));
    LocalMux I__1015 (
            .O(N__8790),
            .I(N__8763));
    LocalMux I__1014 (
            .O(N__8787),
            .I(N__8758));
    Span4Mux_h I__1013 (
            .O(N__8784),
            .I(N__8758));
    LocalMux I__1012 (
            .O(N__8777),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1011 (
            .O(N__8774),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1010 (
            .O(N__8771),
            .I(\uu0.un4_l_count_0 ));
    LocalMux I__1009 (
            .O(N__8768),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1008 (
            .O(N__8763),
            .I(\uu0.un4_l_count_0 ));
    Odrv4 I__1007 (
            .O(N__8758),
            .I(\uu0.un4_l_count_0 ));
    CascadeMux I__1006 (
            .O(N__8745),
            .I(\uu0.un220_ci_cascade_ ));
    InMux I__1005 (
            .O(N__8742),
            .I(N__8738));
    InMux I__1004 (
            .O(N__8741),
            .I(N__8735));
    LocalMux I__1003 (
            .O(N__8738),
            .I(\uu0.l_countZ0Z_18 ));
    LocalMux I__1002 (
            .O(N__8735),
            .I(\uu0.l_countZ0Z_18 ));
    CEMux I__1001 (
            .O(N__8730),
            .I(N__8709));
    CEMux I__1000 (
            .O(N__8729),
            .I(N__8709));
    CEMux I__999 (
            .O(N__8728),
            .I(N__8709));
    CEMux I__998 (
            .O(N__8727),
            .I(N__8709));
    CEMux I__997 (
            .O(N__8726),
            .I(N__8709));
    CEMux I__996 (
            .O(N__8725),
            .I(N__8709));
    CEMux I__995 (
            .O(N__8724),
            .I(N__8709));
    GlobalMux I__994 (
            .O(N__8709),
            .I(N__8706));
    gio2CtrlBuf I__993 (
            .O(N__8706),
            .I(\uu0.un11_l_count_i_g ));
    CascadeMux I__992 (
            .O(N__8703),
            .I(N__8697));
    CascadeMux I__991 (
            .O(N__8702),
            .I(N__8694));
    InMux I__990 (
            .O(N__8701),
            .I(N__8684));
    InMux I__989 (
            .O(N__8700),
            .I(N__8684));
    InMux I__988 (
            .O(N__8697),
            .I(N__8684));
    InMux I__987 (
            .O(N__8694),
            .I(N__8684));
    InMux I__986 (
            .O(N__8693),
            .I(N__8681));
    LocalMux I__985 (
            .O(N__8684),
            .I(\uu0.l_countZ0Z_9 ));
    LocalMux I__984 (
            .O(N__8681),
            .I(\uu0.l_countZ0Z_9 ));
    InMux I__983 (
            .O(N__8676),
            .I(N__8669));
    InMux I__982 (
            .O(N__8675),
            .I(N__8669));
    InMux I__981 (
            .O(N__8674),
            .I(N__8666));
    LocalMux I__980 (
            .O(N__8669),
            .I(N__8663));
    LocalMux I__979 (
            .O(N__8666),
            .I(\uu0.l_countZ0Z_7 ));
    Odrv4 I__978 (
            .O(N__8663),
            .I(\uu0.l_countZ0Z_7 ));
    CascadeMux I__977 (
            .O(N__8658),
            .I(N__8654));
    CascadeMux I__976 (
            .O(N__8657),
            .I(N__8650));
    InMux I__975 (
            .O(N__8654),
            .I(N__8643));
    InMux I__974 (
            .O(N__8653),
            .I(N__8643));
    InMux I__973 (
            .O(N__8650),
            .I(N__8643));
    LocalMux I__972 (
            .O(N__8643),
            .I(\uu0.l_countZ0Z_17 ));
    InMux I__971 (
            .O(N__8640),
            .I(N__8633));
    InMux I__970 (
            .O(N__8639),
            .I(N__8633));
    InMux I__969 (
            .O(N__8638),
            .I(N__8630));
    LocalMux I__968 (
            .O(N__8633),
            .I(\uu0.l_countZ0Z_3 ));
    LocalMux I__967 (
            .O(N__8630),
            .I(\uu0.l_countZ0Z_3 ));
    InMux I__966 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__965 (
            .O(N__8622),
            .I(\uu0.un4_l_count_12 ));
    CascadeMux I__964 (
            .O(N__8619),
            .I(N__8616));
    InMux I__963 (
            .O(N__8616),
            .I(N__8613));
    LocalMux I__962 (
            .O(N__8613),
            .I(N__8608));
    InMux I__961 (
            .O(N__8612),
            .I(N__8600));
    InMux I__960 (
            .O(N__8611),
            .I(N__8600));
    Span4Mux_h I__959 (
            .O(N__8608),
            .I(N__8597));
    InMux I__958 (
            .O(N__8607),
            .I(N__8594));
    InMux I__957 (
            .O(N__8606),
            .I(N__8589));
    InMux I__956 (
            .O(N__8605),
            .I(N__8589));
    LocalMux I__955 (
            .O(N__8600),
            .I(N__8586));
    Odrv4 I__954 (
            .O(N__8597),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__953 (
            .O(N__8594),
            .I(\uu2.r_addrZ0Z_0 ));
    LocalMux I__952 (
            .O(N__8589),
            .I(\uu2.r_addrZ0Z_0 ));
    Odrv12 I__951 (
            .O(N__8586),
            .I(\uu2.r_addrZ0Z_0 ));
    CascadeMux I__950 (
            .O(N__8577),
            .I(N__8574));
    InMux I__949 (
            .O(N__8574),
            .I(N__8571));
    LocalMux I__948 (
            .O(N__8571),
            .I(N__8566));
    InMux I__947 (
            .O(N__8570),
            .I(N__8559));
    InMux I__946 (
            .O(N__8569),
            .I(N__8559));
    Span4Mux_h I__945 (
            .O(N__8566),
            .I(N__8556));
    InMux I__944 (
            .O(N__8565),
            .I(N__8553));
    InMux I__943 (
            .O(N__8564),
            .I(N__8550));
    LocalMux I__942 (
            .O(N__8559),
            .I(N__8547));
    Odrv4 I__941 (
            .O(N__8556),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__940 (
            .O(N__8553),
            .I(\uu2.r_addrZ0Z_1 ));
    LocalMux I__939 (
            .O(N__8550),
            .I(\uu2.r_addrZ0Z_1 ));
    Odrv12 I__938 (
            .O(N__8547),
            .I(\uu2.r_addrZ0Z_1 ));
    CascadeMux I__937 (
            .O(N__8538),
            .I(N__8535));
    InMux I__936 (
            .O(N__8535),
            .I(N__8529));
    InMux I__935 (
            .O(N__8534),
            .I(N__8526));
    InMux I__934 (
            .O(N__8533),
            .I(N__8520));
    InMux I__933 (
            .O(N__8532),
            .I(N__8520));
    LocalMux I__932 (
            .O(N__8529),
            .I(N__8517));
    LocalMux I__931 (
            .O(N__8526),
            .I(N__8514));
    InMux I__930 (
            .O(N__8525),
            .I(N__8511));
    LocalMux I__929 (
            .O(N__8520),
            .I(N__8508));
    Odrv4 I__928 (
            .O(N__8517),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__927 (
            .O(N__8514),
            .I(\uu2.r_addrZ0Z_4 ));
    LocalMux I__926 (
            .O(N__8511),
            .I(\uu2.r_addrZ0Z_4 ));
    Odrv4 I__925 (
            .O(N__8508),
            .I(\uu2.r_addrZ0Z_4 ));
    InMux I__924 (
            .O(N__8499),
            .I(N__8493));
    InMux I__923 (
            .O(N__8498),
            .I(N__8490));
    InMux I__922 (
            .O(N__8497),
            .I(N__8485));
    InMux I__921 (
            .O(N__8496),
            .I(N__8485));
    LocalMux I__920 (
            .O(N__8493),
            .I(N__8480));
    LocalMux I__919 (
            .O(N__8490),
            .I(N__8480));
    LocalMux I__918 (
            .O(N__8485),
            .I(\uu2.un404_ci ));
    Odrv12 I__917 (
            .O(N__8480),
            .I(\uu2.un404_ci ));
    CascadeMux I__916 (
            .O(N__8475),
            .I(N__8472));
    InMux I__915 (
            .O(N__8472),
            .I(N__8468));
    CascadeMux I__914 (
            .O(N__8471),
            .I(N__8465));
    LocalMux I__913 (
            .O(N__8468),
            .I(N__8461));
    InMux I__912 (
            .O(N__8465),
            .I(N__8455));
    InMux I__911 (
            .O(N__8464),
            .I(N__8455));
    Span4Mux_v I__910 (
            .O(N__8461),
            .I(N__8452));
    InMux I__909 (
            .O(N__8460),
            .I(N__8449));
    LocalMux I__908 (
            .O(N__8455),
            .I(N__8446));
    Odrv4 I__907 (
            .O(N__8452),
            .I(\uu2.r_addrZ0Z_5 ));
    LocalMux I__906 (
            .O(N__8449),
            .I(\uu2.r_addrZ0Z_5 ));
    Odrv12 I__905 (
            .O(N__8446),
            .I(\uu2.r_addrZ0Z_5 ));
    CascadeMux I__904 (
            .O(N__8439),
            .I(\uu2.un404_ci_cascade_ ));
    CascadeMux I__903 (
            .O(N__8436),
            .I(N__8433));
    InMux I__902 (
            .O(N__8433),
            .I(N__8429));
    InMux I__901 (
            .O(N__8432),
            .I(N__8426));
    LocalMux I__900 (
            .O(N__8429),
            .I(\uu2.r_addrZ0Z_8 ));
    LocalMux I__899 (
            .O(N__8426),
            .I(\uu2.r_addrZ0Z_8 ));
    InMux I__898 (
            .O(N__8421),
            .I(N__8418));
    LocalMux I__897 (
            .O(N__8418),
            .I(\uu2.vbuf_raddr.un426_ci_3 ));
    CascadeMux I__896 (
            .O(N__8415),
            .I(\uu2.vbuf_raddr.un426_ci_3_cascade_ ));
    CascadeMux I__895 (
            .O(N__8412),
            .I(N__8409));
    InMux I__894 (
            .O(N__8409),
            .I(N__8404));
    InMux I__893 (
            .O(N__8408),
            .I(N__8401));
    InMux I__892 (
            .O(N__8407),
            .I(N__8398));
    LocalMux I__891 (
            .O(N__8404),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__890 (
            .O(N__8401),
            .I(\uu2.r_addrZ0Z_7 ));
    LocalMux I__889 (
            .O(N__8398),
            .I(\uu2.r_addrZ0Z_7 ));
    InMux I__888 (
            .O(N__8391),
            .I(N__8388));
    LocalMux I__887 (
            .O(N__8388),
            .I(\uu2.vbuf_raddr.un448_ci_0 ));
    CascadeMux I__886 (
            .O(N__8385),
            .I(N__8382));
    InMux I__885 (
            .O(N__8382),
            .I(N__8376));
    InMux I__884 (
            .O(N__8381),
            .I(N__8373));
    InMux I__883 (
            .O(N__8380),
            .I(N__8368));
    InMux I__882 (
            .O(N__8379),
            .I(N__8368));
    LocalMux I__881 (
            .O(N__8376),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__880 (
            .O(N__8373),
            .I(\uu2.r_addrZ0Z_6 ));
    LocalMux I__879 (
            .O(N__8368),
            .I(\uu2.r_addrZ0Z_6 ));
    CascadeMux I__878 (
            .O(N__8361),
            .I(N__8358));
    InMux I__877 (
            .O(N__8358),
            .I(N__8353));
    CascadeMux I__876 (
            .O(N__8357),
            .I(N__8350));
    CascadeMux I__875 (
            .O(N__8356),
            .I(N__8347));
    LocalMux I__874 (
            .O(N__8353),
            .I(N__8344));
    InMux I__873 (
            .O(N__8350),
            .I(N__8339));
    InMux I__872 (
            .O(N__8347),
            .I(N__8339));
    Odrv4 I__871 (
            .O(N__8344),
            .I(\uu2.r_addrZ0Z_3 ));
    LocalMux I__870 (
            .O(N__8339),
            .I(\uu2.r_addrZ0Z_3 ));
    CEMux I__869 (
            .O(N__8334),
            .I(N__8331));
    LocalMux I__868 (
            .O(N__8331),
            .I(\uu2.trig_rd_is_det_0 ));
    CascadeMux I__867 (
            .O(N__8328),
            .I(N__8325));
    InMux I__866 (
            .O(N__8325),
            .I(N__8319));
    CascadeMux I__865 (
            .O(N__8324),
            .I(N__8316));
    InMux I__864 (
            .O(N__8323),
            .I(N__8311));
    InMux I__863 (
            .O(N__8322),
            .I(N__8311));
    LocalMux I__862 (
            .O(N__8319),
            .I(N__8308));
    InMux I__861 (
            .O(N__8316),
            .I(N__8305));
    LocalMux I__860 (
            .O(N__8311),
            .I(N__8302));
    Odrv4 I__859 (
            .O(N__8308),
            .I(\uu2.r_addrZ0Z_2 ));
    LocalMux I__858 (
            .O(N__8305),
            .I(\uu2.r_addrZ0Z_2 ));
    Odrv4 I__857 (
            .O(N__8302),
            .I(\uu2.r_addrZ0Z_2 ));
    InMux I__856 (
            .O(N__8295),
            .I(N__8292));
    LocalMux I__855 (
            .O(N__8292),
            .I(\uu2.mem0.N_31_i ));
    CascadeMux I__854 (
            .O(N__8289),
            .I(\uu2.mem0.N_61_cascade_ ));
    InMux I__853 (
            .O(N__8286),
            .I(N__8283));
    LocalMux I__852 (
            .O(N__8283),
            .I(\uu2.mem0.w_data_1 ));
    InMux I__851 (
            .O(N__8280),
            .I(N__8277));
    LocalMux I__850 (
            .O(N__8277),
            .I(\uu2.mem0.w_data_4 ));
    InMux I__849 (
            .O(N__8274),
            .I(N__8271));
    LocalMux I__848 (
            .O(N__8271),
            .I(\uu2.N_922_tz_tz ));
    InMux I__847 (
            .O(N__8268),
            .I(N__8265));
    LocalMux I__846 (
            .O(N__8265),
            .I(\uu2.bitmap_pmux ));
    CascadeMux I__845 (
            .O(N__8262),
            .I(\uu2.bitmap_pmux_cascade_ ));
    InMux I__844 (
            .O(N__8259),
            .I(N__8256));
    LocalMux I__843 (
            .O(N__8256),
            .I(\uu2.mem0.w_data_3 ));
    InMux I__842 (
            .O(N__8253),
            .I(N__8249));
    CascadeMux I__841 (
            .O(N__8252),
            .I(N__8246));
    LocalMux I__840 (
            .O(N__8249),
            .I(N__8243));
    InMux I__839 (
            .O(N__8246),
            .I(N__8240));
    Odrv4 I__838 (
            .O(N__8243),
            .I(\uu2.N_37 ));
    LocalMux I__837 (
            .O(N__8240),
            .I(\uu2.N_37 ));
    InMux I__836 (
            .O(N__8235),
            .I(N__8232));
    LocalMux I__835 (
            .O(N__8232),
            .I(\uu2.mem0.N_59 ));
    InMux I__834 (
            .O(N__8229),
            .I(N__8226));
    LocalMux I__833 (
            .O(N__8226),
            .I(\uu2.mem0.w_data_0 ));
    CascadeMux I__832 (
            .O(N__8223),
            .I(N__8218));
    InMux I__831 (
            .O(N__8222),
            .I(N__8208));
    InMux I__830 (
            .O(N__8221),
            .I(N__8208));
    InMux I__829 (
            .O(N__8218),
            .I(N__8208));
    InMux I__828 (
            .O(N__8217),
            .I(N__8208));
    LocalMux I__827 (
            .O(N__8208),
            .I(\uu0.un154_ci_9 ));
    InMux I__826 (
            .O(N__8205),
            .I(N__8200));
    InMux I__825 (
            .O(N__8204),
            .I(N__8195));
    InMux I__824 (
            .O(N__8203),
            .I(N__8195));
    LocalMux I__823 (
            .O(N__8200),
            .I(N__8192));
    LocalMux I__822 (
            .O(N__8195),
            .I(\uu0.l_countZ0Z_15 ));
    Odrv4 I__821 (
            .O(N__8192),
            .I(\uu0.l_countZ0Z_15 ));
    CascadeMux I__820 (
            .O(N__8187),
            .I(\uu0.un4_l_count_0_8_cascade_ ));
    CascadeMux I__819 (
            .O(N__8184),
            .I(N__8178));
    InMux I__818 (
            .O(N__8183),
            .I(N__8175));
    InMux I__817 (
            .O(N__8182),
            .I(N__8170));
    InMux I__816 (
            .O(N__8181),
            .I(N__8170));
    InMux I__815 (
            .O(N__8178),
            .I(N__8167));
    LocalMux I__814 (
            .O(N__8175),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__813 (
            .O(N__8170),
            .I(\uu0.l_countZ0Z_14 ));
    LocalMux I__812 (
            .O(N__8167),
            .I(\uu0.l_countZ0Z_14 ));
    InMux I__811 (
            .O(N__8160),
            .I(N__8154));
    InMux I__810 (
            .O(N__8159),
            .I(N__8151));
    InMux I__809 (
            .O(N__8158),
            .I(N__8148));
    InMux I__808 (
            .O(N__8157),
            .I(N__8145));
    LocalMux I__807 (
            .O(N__8154),
            .I(N__8140));
    LocalMux I__806 (
            .O(N__8151),
            .I(N__8140));
    LocalMux I__805 (
            .O(N__8148),
            .I(\uu0.l_countZ0Z_4 ));
    LocalMux I__804 (
            .O(N__8145),
            .I(\uu0.l_countZ0Z_4 ));
    Odrv4 I__803 (
            .O(N__8140),
            .I(\uu0.l_countZ0Z_4 ));
    InMux I__802 (
            .O(N__8133),
            .I(N__8128));
    InMux I__801 (
            .O(N__8132),
            .I(N__8125));
    InMux I__800 (
            .O(N__8131),
            .I(N__8122));
    LocalMux I__799 (
            .O(N__8128),
            .I(N__8119));
    LocalMux I__798 (
            .O(N__8125),
            .I(\uu0.l_countZ0Z_5 ));
    LocalMux I__797 (
            .O(N__8122),
            .I(\uu0.l_countZ0Z_5 ));
    Odrv12 I__796 (
            .O(N__8119),
            .I(\uu0.l_countZ0Z_5 ));
    CascadeMux I__795 (
            .O(N__8112),
            .I(\uu2.N_34_cascade_ ));
    InMux I__794 (
            .O(N__8109),
            .I(N__8106));
    LocalMux I__793 (
            .O(N__8106),
            .I(\uu2.N_114 ));
    InMux I__792 (
            .O(N__8103),
            .I(N__8100));
    LocalMux I__791 (
            .O(N__8100),
            .I(N__8097));
    Odrv4 I__790 (
            .O(N__8097),
            .I(\uu2.mem0.w_data_6 ));
    CascadeMux I__789 (
            .O(N__8094),
            .I(N__8091));
    InMux I__788 (
            .O(N__8091),
            .I(N__8085));
    InMux I__787 (
            .O(N__8090),
            .I(N__8078));
    InMux I__786 (
            .O(N__8089),
            .I(N__8078));
    InMux I__785 (
            .O(N__8088),
            .I(N__8078));
    LocalMux I__784 (
            .O(N__8085),
            .I(\uu0.l_countZ0Z_10 ));
    LocalMux I__783 (
            .O(N__8078),
            .I(\uu0.l_countZ0Z_10 ));
    InMux I__782 (
            .O(N__8073),
            .I(N__8070));
    LocalMux I__781 (
            .O(N__8070),
            .I(N__8067));
    Odrv4 I__780 (
            .O(N__8067),
            .I(\uu0.un143_ci_0 ));
    InMux I__779 (
            .O(N__8064),
            .I(N__8046));
    InMux I__778 (
            .O(N__8063),
            .I(N__8046));
    InMux I__777 (
            .O(N__8062),
            .I(N__8046));
    InMux I__776 (
            .O(N__8061),
            .I(N__8046));
    InMux I__775 (
            .O(N__8060),
            .I(N__8046));
    InMux I__774 (
            .O(N__8059),
            .I(N__8046));
    LocalMux I__773 (
            .O(N__8046),
            .I(\uu0.l_countZ0Z_8 ));
    CascadeMux I__772 (
            .O(N__8043),
            .I(\uu0.un187_ci_1_cascade_ ));
    CascadeMux I__771 (
            .O(N__8040),
            .I(N__8037));
    InMux I__770 (
            .O(N__8037),
            .I(N__8034));
    LocalMux I__769 (
            .O(N__8034),
            .I(\uu0.un165_ci_0 ));
    InMux I__768 (
            .O(N__8031),
            .I(N__8025));
    InMux I__767 (
            .O(N__8030),
            .I(N__8025));
    LocalMux I__766 (
            .O(N__8025),
            .I(\uu0.l_countZ0Z_13 ));
    InMux I__765 (
            .O(N__8022),
            .I(N__8013));
    InMux I__764 (
            .O(N__8021),
            .I(N__8013));
    InMux I__763 (
            .O(N__8020),
            .I(N__8013));
    LocalMux I__762 (
            .O(N__8013),
            .I(\uu0.l_countZ0Z_12 ));
    InMux I__761 (
            .O(N__8010),
            .I(N__8005));
    InMux I__760 (
            .O(N__8009),
            .I(N__8000));
    InMux I__759 (
            .O(N__8008),
            .I(N__8000));
    LocalMux I__758 (
            .O(N__8005),
            .I(\uu0.un4_l_count_0_8 ));
    LocalMux I__757 (
            .O(N__8000),
            .I(\uu0.un4_l_count_0_8 ));
    CascadeMux I__756 (
            .O(N__7995),
            .I(\uu0.un55_ci_cascade_ ));
    CascadeMux I__755 (
            .O(N__7992),
            .I(N__7985));
    InMux I__754 (
            .O(N__7991),
            .I(N__7971));
    InMux I__753 (
            .O(N__7990),
            .I(N__7971));
    InMux I__752 (
            .O(N__7989),
            .I(N__7971));
    InMux I__751 (
            .O(N__7988),
            .I(N__7971));
    InMux I__750 (
            .O(N__7985),
            .I(N__7971));
    InMux I__749 (
            .O(N__7984),
            .I(N__7971));
    LocalMux I__748 (
            .O(N__7971),
            .I(\uu0.l_countZ0Z_0 ));
    InMux I__747 (
            .O(N__7968),
            .I(N__7955));
    InMux I__746 (
            .O(N__7967),
            .I(N__7955));
    InMux I__745 (
            .O(N__7966),
            .I(N__7955));
    InMux I__744 (
            .O(N__7965),
            .I(N__7955));
    InMux I__743 (
            .O(N__7964),
            .I(N__7952));
    LocalMux I__742 (
            .O(N__7955),
            .I(\uu0.l_countZ0Z_1 ));
    LocalMux I__741 (
            .O(N__7952),
            .I(\uu0.l_countZ0Z_1 ));
    CascadeMux I__740 (
            .O(N__7947),
            .I(N__7943));
    CascadeMux I__739 (
            .O(N__7946),
            .I(N__7940));
    InMux I__738 (
            .O(N__7943),
            .I(N__7931));
    InMux I__737 (
            .O(N__7940),
            .I(N__7931));
    InMux I__736 (
            .O(N__7939),
            .I(N__7931));
    InMux I__735 (
            .O(N__7938),
            .I(N__7928));
    LocalMux I__734 (
            .O(N__7931),
            .I(\uu0.l_countZ0Z_2 ));
    LocalMux I__733 (
            .O(N__7928),
            .I(\uu0.l_countZ0Z_2 ));
    CascadeMux I__732 (
            .O(N__7923),
            .I(N__7918));
    CascadeMux I__731 (
            .O(N__7922),
            .I(N__7912));
    InMux I__730 (
            .O(N__7921),
            .I(N__7909));
    InMux I__729 (
            .O(N__7918),
            .I(N__7906));
    InMux I__728 (
            .O(N__7917),
            .I(N__7897));
    InMux I__727 (
            .O(N__7916),
            .I(N__7897));
    InMux I__726 (
            .O(N__7915),
            .I(N__7897));
    InMux I__725 (
            .O(N__7912),
            .I(N__7897));
    LocalMux I__724 (
            .O(N__7909),
            .I(N__7894));
    LocalMux I__723 (
            .O(N__7906),
            .I(\uu0.l_precountZ0Z_0 ));
    LocalMux I__722 (
            .O(N__7897),
            .I(\uu0.l_precountZ0Z_0 ));
    Odrv4 I__721 (
            .O(N__7894),
            .I(\uu0.l_precountZ0Z_0 ));
    CascadeMux I__720 (
            .O(N__7887),
            .I(\uu0.un4_l_count_14_cascade_ ));
    InMux I__719 (
            .O(N__7884),
            .I(N__7881));
    LocalMux I__718 (
            .O(N__7881),
            .I(N__7878));
    Odrv4 I__717 (
            .O(N__7878),
            .I(\uu0.un4_l_count_18 ));
    InMux I__716 (
            .O(N__7875),
            .I(N__7870));
    InMux I__715 (
            .O(N__7874),
            .I(N__7865));
    InMux I__714 (
            .O(N__7873),
            .I(N__7865));
    LocalMux I__713 (
            .O(N__7870),
            .I(\uu0.l_countZ0Z_11 ));
    LocalMux I__712 (
            .O(N__7865),
            .I(\uu0.l_countZ0Z_11 ));
    CascadeMux I__711 (
            .O(N__7860),
            .I(\uu0.un154_ci_9_cascade_ ));
    InMux I__710 (
            .O(N__7857),
            .I(N__7846));
    InMux I__709 (
            .O(N__7856),
            .I(N__7846));
    InMux I__708 (
            .O(N__7855),
            .I(N__7846));
    InMux I__707 (
            .O(N__7854),
            .I(N__7841));
    InMux I__706 (
            .O(N__7853),
            .I(N__7841));
    LocalMux I__705 (
            .O(N__7846),
            .I(\uu0.l_precountZ0Z_1 ));
    LocalMux I__704 (
            .O(N__7841),
            .I(\uu0.l_precountZ0Z_1 ));
    CascadeMux I__703 (
            .O(N__7836),
            .I(N__7831));
    InMux I__702 (
            .O(N__7835),
            .I(N__7828));
    InMux I__701 (
            .O(N__7834),
            .I(N__7823));
    InMux I__700 (
            .O(N__7831),
            .I(N__7823));
    LocalMux I__699 (
            .O(N__7828),
            .I(\uu0.l_precountZ0Z_3 ));
    LocalMux I__698 (
            .O(N__7823),
            .I(\uu0.l_precountZ0Z_3 ));
    CascadeMux I__697 (
            .O(N__7818),
            .I(\uu0.un4_l_count_11_cascade_ ));
    CascadeMux I__696 (
            .O(N__7815),
            .I(\uu0.un4_l_count_16_cascade_ ));
    InMux I__695 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__694 (
            .O(N__7809),
            .I(\uu0.delay_lineZ0Z_1 ));
    CascadeMux I__693 (
            .O(N__7806),
            .I(\uu0.un4_l_count_0_cascade_ ));
    InMux I__692 (
            .O(N__7803),
            .I(N__7799));
    InMux I__691 (
            .O(N__7802),
            .I(N__7796));
    LocalMux I__690 (
            .O(N__7799),
            .I(\uu0.delay_lineZ0Z_0 ));
    LocalMux I__689 (
            .O(N__7796),
            .I(\uu0.delay_lineZ0Z_0 ));
    IoInMux I__688 (
            .O(N__7791),
            .I(N__7788));
    LocalMux I__687 (
            .O(N__7788),
            .I(\uu0.un11_l_count_i ));
    CascadeMux I__686 (
            .O(N__7785),
            .I(N__7782));
    InMux I__685 (
            .O(N__7782),
            .I(N__7776));
    InMux I__684 (
            .O(N__7781),
            .I(N__7773));
    InMux I__683 (
            .O(N__7780),
            .I(N__7768));
    InMux I__682 (
            .O(N__7779),
            .I(N__7768));
    LocalMux I__681 (
            .O(N__7776),
            .I(N__7765));
    LocalMux I__680 (
            .O(N__7773),
            .I(\uu0.l_precountZ0Z_2 ));
    LocalMux I__679 (
            .O(N__7768),
            .I(\uu0.l_precountZ0Z_2 ));
    Odrv4 I__678 (
            .O(N__7765),
            .I(\uu0.l_precountZ0Z_2 ));
    InMux I__677 (
            .O(N__7758),
            .I(N__7755));
    LocalMux I__676 (
            .O(N__7755),
            .I(\uu0.un4_l_count_13 ));
    CascadeMux I__675 (
            .O(N__7752),
            .I(N__7749));
    InMux I__674 (
            .O(N__7749),
            .I(N__7746));
    LocalMux I__673 (
            .O(N__7746),
            .I(N__7743));
    Span4Mux_s2_v I__672 (
            .O(N__7743),
            .I(N__7740));
    Odrv4 I__671 (
            .O(N__7740),
            .I(\uu2.mem0.N_139 ));
    InMux I__670 (
            .O(N__7737),
            .I(N__7734));
    LocalMux I__669 (
            .O(N__7734),
            .I(N__7731));
    IoSpan4Mux I__668 (
            .O(N__7731),
            .I(N__7728));
    Odrv4 I__667 (
            .O(N__7728),
            .I(uart_RXD));
    CascadeMux I__666 (
            .O(N__7725),
            .I(N__7722));
    InMux I__665 (
            .O(N__7722),
            .I(N__7719));
    LocalMux I__664 (
            .O(N__7719),
            .I(N__7716));
    Odrv4 I__663 (
            .O(N__7716),
            .I(\uu2.mem0.N_137 ));
    CascadeMux I__662 (
            .O(N__7713),
            .I(N__7710));
    InMux I__661 (
            .O(N__7710),
            .I(N__7707));
    LocalMux I__660 (
            .O(N__7707),
            .I(N__7704));
    Odrv4 I__659 (
            .O(N__7704),
            .I(\uu2.mem0.N_141 ));
    CascadeMux I__658 (
            .O(N__7701),
            .I(\uu2.bitmap_pmux_u_0_a2_0_cascade_ ));
    CascadeMux I__657 (
            .O(N__7698),
            .I(N__7695));
    InMux I__656 (
            .O(N__7695),
            .I(N__7692));
    LocalMux I__655 (
            .O(N__7692),
            .I(N__7689));
    Odrv4 I__654 (
            .O(N__7689),
            .I(\uu2.mem0.N_140 ));
    IoInMux I__653 (
            .O(N__7686),
            .I(N__7683));
    LocalMux I__652 (
            .O(N__7683),
            .I(N__7680));
    IoSpan4Mux I__651 (
            .O(N__7680),
            .I(N__7677));
    Odrv4 I__650 (
            .O(N__7677),
            .I(clk_in_c));
    INV \INVuu2.w_addr_user_7C  (
            .O(\INVuu2.w_addr_user_7C_net ),
            .I(N__21656));
    INV \INVuu2.w_addr_user_nesr_5C  (
            .O(\INVuu2.w_addr_user_nesr_5C_net ),
            .I(N__21622));
    INV \INVuu2.bitmap_308C  (
            .O(\INVuu2.bitmap_308C_net ),
            .I(N__21645));
    INV \INVuu2.bitmap_296C  (
            .O(\INVuu2.bitmap_296C_net ),
            .I(N__21653));
    INV \INVuu2.bitmap_168C  (
            .O(\INVuu2.bitmap_168C_net ),
            .I(N__21659));
    INV \INVuu2.bitmap_314C  (
            .O(\INVuu2.bitmap_314C_net ),
            .I(N__21649));
    INV \INVuu2.w_addr_displaying_3_rep1C  (
            .O(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .I(N__21662));
    INV \INVuu2.bitmap_194C  (
            .O(\INVuu2.bitmap_194C_net ),
            .I(N__21669));
    INV \INVuu2.r_data_reg_0C  (
            .O(\INVuu2.r_data_reg_0C_net ),
            .I(N__21625));
    INV \INVuu2.w_addr_user_nesr_8C  (
            .O(\INVuu2.w_addr_user_nesr_8C_net ),
            .I(N__21648));
    INV \INVuu2.w_addr_displaying_nesr_7C  (
            .O(\INVuu2.w_addr_displaying_nesr_7C_net ),
            .I(N__21655));
    INV \INVuu2.bitmap_186C  (
            .O(\INVuu2.bitmap_186C_net ),
            .I(N__21661));
    INV \INVuu2.w_addr_displaying_fast_2C  (
            .O(\INVuu2.w_addr_displaying_fast_2C_net ),
            .I(N__21668));
    INV \INVuu2.w_addr_displaying_nesr_4C  (
            .O(\INVuu2.w_addr_displaying_nesr_4C_net ),
            .I(N__21672));
    INV \INVuu2.w_addr_user_4C  (
            .O(\INVuu2.w_addr_user_4C_net ),
            .I(N__21654));
    INV \INVuu2.w_addr_user_1C  (
            .O(\INVuu2.w_addr_user_1C_net ),
            .I(N__21660));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    ICE_GB \latticehx1k_pll_inst.latticehx1k_pll_inst_RNIQV8B  (
            .USERSIGNALTOGLOBALBUFFER(N__9759),
            .GLOBALBUFFEROUTPUT(clk_g));
    ICE_GB bu_rx_data_rdy_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__19437),
            .GLOBALBUFFEROUTPUT(bu_rx_data_rdy_0_g));
    ICE_GB \buart.Z_rx.bitcount_es_RNIV4M42_0_0  (
            .USERSIGNALTOGLOBALBUFFER(N__11844),
            .GLOBALBUFFEROUTPUT(\buart.Z_rx.sample_g ));
    ICE_GB \uu0.delay_line_RNILLLG7_0_1  (
            .USERSIGNALTOGLOBALBUFFER(N__7791),
            .GLOBALBUFFEROUTPUT(\uu0.un11_l_count_i_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB \resetGen.rst_RNI4PQ1  (
            .USERSIGNALTOGLOBALBUFFER(N__15585),
            .GLOBALBUFFEROUTPUT(rst_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_1_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_3_LC_1_3_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_3_LC_1_3_0  (
            .in0(N__10329),
            .in1(N__11257),
            .in2(N__12927),
            .in3(N__9399),
            .lcout(\uu2.mem0.N_137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_1_3_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_LC_1_3_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_LC_1_3_2  (
            .in0(N__10330),
            .in1(N__12381),
            .in2(N__9585),
            .in3(N__11259),
            .lcout(\uu2.mem0.N_141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIFPHP1_3_LC_1_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIFPHP1_3_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIFPHP1_3_LC_1_3_3 .LUT_INIT=16'b0100000000001000;
    LogicCell40 \uu2.w_addr_displaying_RNIFPHP1_3_LC_1_3_3  (
            .in0(N__10706),
            .in1(N__9411),
            .in2(N__10604),
            .in3(N__10402),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_u_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIUI3J3_3_LC_1_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIUI3J3_3_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIUI3J3_3_LC_1_3_4 .LUT_INIT=16'b1111011011110000;
    LogicCell40 \uu2.w_addr_displaying_RNIUI3J3_3_LC_1_3_4  (
            .in0(N__10403),
            .in1(N__10600),
            .in2(N__7701),
            .in3(N__8109),
            .lcout(\uu2.N_922_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_1_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_0_LC_1_3_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_0_LC_1_3_6  (
            .in0(N__10404),
            .in1(N__10331),
            .in2(N__9637),
            .in3(N__11258),
            .lcout(\uu2.mem0.N_140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_1_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_1_LC_1_3_7 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_1_LC_1_3_7  (
            .in0(N__11256),
            .in1(N__9858),
            .in2(N__10710),
            .in3(N__10328),
            .lcout(\uu2.mem0.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_1_LC_1_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_1_LC_1_6_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_1_LC_1_6_3 .LUT_INIT=16'b0001001011110000;
    LogicCell40 \uu2.w_addr_user_1_LC_1_6_3  (
            .in0(N__9584),
            .in1(N__14084),
            .in2(N__9631),
            .in3(N__13997),
            .lcout(\uu2.w_addr_userZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_1C_net ),
            .ce(),
            .sr(N__19166));
    defparam \uu0.l_count_6_LC_1_8_3 .C_ON=1'b0;
    defparam \uu0.l_count_6_LC_1_8_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_6_LC_1_8_3 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_6_LC_1_8_3  (
            .in0(N__8951),
            .in1(N__8809),
            .in2(N__9123),
            .in3(N__9084),
            .lcout(\uu0.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21646),
            .ce(N__8725),
            .sr(N__19216));
    defparam \buart.Z_rx.hh_1_LC_1_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_1_LC_1_9_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_1_LC_1_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_1_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11558),
            .lcout(\buart.Z_rx.hhZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \buart.Z_rx.hh_0_LC_1_9_1 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_0_LC_1_9_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.hh_0_LC_1_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.hh_0_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7737),
            .lcout(\buart.Z_rx.hhZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.l_precount_0_LC_1_9_2 .C_ON=1'b0;
    defparam \uu0.l_precount_0_LC_1_9_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_0_LC_1_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uu0.l_precount_0_LC_1_9_2  (
            .in0(N__7915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu0.l_precountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.delay_line_1_LC_1_9_3 .C_ON=1'b0;
    defparam \uu0.delay_line_1_LC_1_9_3 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_1_LC_1_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu0.delay_line_1_LC_1_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7803),
            .lcout(\uu0.delay_lineZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.delay_line_0_LC_1_9_4 .C_ON=1'b0;
    defparam \uu0.delay_line_0_LC_1_9_4 .SEQ_MODE=4'b1010;
    defparam \uu0.delay_line_0_LC_1_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.delay_line_0_LC_1_9_4  (
            .in0(N__7779),
            .in1(N__7835),
            .in2(N__7922),
            .in3(N__7855),
            .lcout(\uu0.delay_lineZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.l_precount_2_LC_1_9_5 .C_ON=1'b0;
    defparam \uu0.l_precount_2_LC_1_9_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_2_LC_1_9_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_precount_2_LC_1_9_5  (
            .in0(N__7857),
            .in1(N__7917),
            .in2(_gnd_net_),
            .in3(N__7780),
            .lcout(\uu0.l_precountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.l_precount_1_LC_1_9_7 .C_ON=1'b0;
    defparam \uu0.l_precount_1_LC_1_9_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_1_LC_1_9_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_precount_1_LC_1_9_7  (
            .in0(N__7856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7916),
            .lcout(\uu0.l_precountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21641),
            .ce(),
            .sr(N__19217));
    defparam \uu0.l_precount_3_LC_1_10_1 .C_ON=1'b0;
    defparam \uu0.l_precount_3_LC_1_10_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_precount_3_LC_1_10_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu0.l_precount_3_LC_1_10_1  (
            .in0(N__7781),
            .in1(N__7834),
            .in2(N__7923),
            .in3(N__7854),
            .lcout(\uu0.l_precountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21632),
            .ce(),
            .sr(N__19218));
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_4 .C_ON=1'b0;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \uu0.l_precount_RNI85Q91_3_LC_1_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_precount_RNI85Q91_3_LC_1_10_4  (
            .in0(N__7853),
            .in1(N__8133),
            .in2(N__7836),
            .in3(N__7964),
            .lcout(),
            .ltout(\uu0.un4_l_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI96A32_18_LC_1_10_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNI96A32_18_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI96A32_18_LC_1_10_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI96A32_18_LC_1_10_5  (
            .in0(N__8205),
            .in1(N__8741),
            .in2(N__7818),
            .in3(N__9085),
            .lcout(),
            .ltout(\uu0.un4_l_count_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_10_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI8ORT6_11_LC_1_10_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.l_count_RNI8ORT6_11_LC_1_10_6  (
            .in0(N__7758),
            .in1(N__8625),
            .in2(N__7815),
            .in3(N__7884),
            .lcout(\uu0.un4_l_count_0 ),
            .ltout(\uu0.un4_l_count_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_7 .C_ON=1'b0;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \uu0.delay_line_RNILLLG7_1_LC_1_10_7 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \uu0.delay_line_RNILLLG7_1_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__7812),
            .in2(N__7806),
            .in3(N__7802),
            .lcout(\uu0.un11_l_count_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2CNU_11_LC_1_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2CNU_11_LC_1_11_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uu0.l_count_RNI2CNU_11_LC_1_11_0  (
            .in0(N__8832),
            .in1(N__7873),
            .in2(N__7785),
            .in3(N__7984),
            .lcout(\uu0.un4_l_count_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_6_LC_1_11_1  (
            .in0(N__8639),
            .in1(N__7939),
            .in2(N__7992),
            .in3(N__7965),
            .lcout(\uu0.un66_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_2_LC_1_11_2 .C_ON=1'b0;
    defparam \uu0.l_count_2_LC_1_11_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_2_LC_1_11_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uu0.l_count_2_LC_1_11_2  (
            .in0(N__7968),
            .in1(_gnd_net_),
            .in2(N__7947),
            .in3(N__7991),
            .lcout(\uu0.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__8726),
            .sr(N__19220));
    defparam \uu0.l_count_0_LC_1_11_3 .C_ON=1'b0;
    defparam \uu0.l_count_0_LC_1_11_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_0_LC_1_11_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uu0.l_count_0_LC_1_11_3  (
            .in0(N__7989),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8803),
            .lcout(\uu0.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__8726),
            .sr(N__19220));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_3__un55_ci_LC_1_11_4  (
            .in0(N__7966),
            .in1(_gnd_net_),
            .in2(N__7946),
            .in3(N__7988),
            .lcout(),
            .ltout(\uu0.un55_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_3_LC_1_11_5 .C_ON=1'b0;
    defparam \uu0.l_count_3_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_3_LC_1_11_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \uu0.l_count_3_LC_1_11_5  (
            .in0(N__8640),
            .in1(_gnd_net_),
            .in2(N__7995),
            .in3(N__8805),
            .lcout(\uu0.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__8726),
            .sr(N__19220));
    defparam \uu0.l_count_1_LC_1_11_6 .C_ON=1'b0;
    defparam \uu0.l_count_1_LC_1_11_6 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_1_LC_1_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_1_LC_1_11_6  (
            .in0(N__7967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7990),
            .lcout(\uu0.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__8726),
            .sr(N__19220));
    defparam \uu0.l_count_11_LC_1_11_7 .C_ON=1'b0;
    defparam \uu0.l_count_11_LC_1_11_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_11_LC_1_11_7 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \uu0.l_count_11_LC_1_11_7  (
            .in0(N__7874),
            .in1(N__8073),
            .in2(N__8899),
            .in3(N__8804),
            .lcout(\uu0.l_countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21623),
            .ce(N__8726),
            .sr(N__19220));
    defparam \uu0.l_count_RNI04591_10_LC_1_12_0 .C_ON=1'b0;
    defparam \uu0.l_count_RNI04591_10_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI04591_10_LC_1_12_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu0.l_count_RNI04591_10_LC_1_12_0  (
            .in0(N__8088),
            .in1(N__8059),
            .in2(N__8184),
            .in3(N__7938),
            .lcout(),
            .ltout(\uu0.un4_l_count_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNI2GS72_4_LC_1_12_1 .C_ON=1'b0;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNI2GS72_4_LC_1_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu0.l_count_RNI2GS72_4_LC_1_12_1  (
            .in0(N__7921),
            .in1(N__8159),
            .in2(N__7887),
            .in3(N__8008),
            .lcout(\uu0.un4_l_count_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_12_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_12__un154_ci_9_LC_1_12_2  (
            .in0(N__8089),
            .in1(N__7875),
            .in2(N__8702),
            .in3(N__8060),
            .lcout(\uu0.un154_ci_9 ),
            .ltout(\uu0.un154_ci_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_14_LC_1_12_3 .C_ON=1'b0;
    defparam \uu0.l_count_14_LC_1_12_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_14_LC_1_12_3 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uu0.l_count_14_LC_1_12_3  (
            .in0(N__8183),
            .in1(N__8883),
            .in2(N__7860),
            .in3(N__8009),
            .lcout(\uu0.l_countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(N__8727),
            .sr(N__19222));
    defparam \uu0.l_count_8_LC_1_12_4 .C_ON=1'b0;
    defparam \uu0.l_count_8_LC_1_12_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_8_LC_1_12_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu0.l_count_8_LC_1_12_4  (
            .in0(N__8882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8063),
            .lcout(\uu0.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(N__8727),
            .sr(N__19222));
    defparam \uu0.l_count_10_LC_1_12_5 .C_ON=1'b0;
    defparam \uu0.l_count_10_LC_1_12_5 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_10_LC_1_12_5 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu0.l_count_10_LC_1_12_5  (
            .in0(N__8062),
            .in1(N__8700),
            .in2(N__8094),
            .in3(N__8885),
            .lcout(\uu0.l_countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(N__8727),
            .sr(N__19222));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_11__un143_ci_0_LC_1_12_6  (
            .in0(N__8090),
            .in1(_gnd_net_),
            .in2(N__8703),
            .in3(N__8061),
            .lcout(\uu0.un143_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_9_LC_1_12_7 .C_ON=1'b0;
    defparam \uu0.l_count_9_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_9_LC_1_12_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_9_LC_1_12_7  (
            .in0(N__8064),
            .in1(N__8884),
            .in2(_gnd_net_),
            .in3(N__8701),
            .lcout(\uu0.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21616),
            .ce(N__8727),
            .sr(N__19222));
    defparam \uu0.l_count_13_LC_1_13_0 .C_ON=1'b0;
    defparam \uu0.l_count_13_LC_1_13_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_13_LC_1_13_0 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \uu0.l_count_13_LC_1_13_0  (
            .in0(N__8031),
            .in1(N__8813),
            .in2(N__8040),
            .in3(N__8909),
            .lcout(\uu0.l_countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21611),
            .ce(N__8729),
            .sr(N__19226));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_13_1 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_15__un187_ci_1_LC_1_13_1  (
            .in0(N__8182),
            .in1(N__8221),
            .in2(_gnd_net_),
            .in3(N__8010),
            .lcout(),
            .ltout(\uu0.un187_ci_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_15_LC_1_13_2 .C_ON=1'b0;
    defparam \uu0.l_count_15_LC_1_13_2 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_15_LC_1_13_2 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_15_LC_1_13_2  (
            .in0(N__8910),
            .in1(N__8814),
            .in2(N__8043),
            .in3(N__8204),
            .lcout(\uu0.l_countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21611),
            .ce(N__8729),
            .sr(N__19226));
    defparam \uu0.l_count_12_LC_1_13_3 .C_ON=1'b0;
    defparam \uu0.l_count_12_LC_1_13_3 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_12_LC_1_13_3 .LUT_INIT=16'b0000011000001100;
    LogicCell40 \uu0.l_count_12_LC_1_13_3  (
            .in0(N__8908),
            .in1(N__8022),
            .in2(N__8817),
            .in3(N__8222),
            .lcout(\uu0.l_countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21611),
            .ce(N__8729),
            .sr(N__19226));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_13_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_13_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_13__un165_ci_0_LC_1_13_4  (
            .in0(N__8021),
            .in1(_gnd_net_),
            .in2(N__8223),
            .in3(_gnd_net_),
            .lcout(\uu0.un165_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_13_5 .C_ON=1'b0;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIFAQ9_13_LC_1_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.l_count_RNIFAQ9_13_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__8030),
            .in2(_gnd_net_),
            .in3(N__8020),
            .lcout(\uu0.un4_l_count_0_8 ),
            .ltout(\uu0.un4_l_count_0_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_13_6 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_16__un198_ci_2_LC_1_13_6  (
            .in0(N__8217),
            .in1(N__8203),
            .in2(N__8187),
            .in3(N__8181),
            .lcout(\uu0.un198_ci_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_4_LC_1_13_7 .C_ON=1'b0;
    defparam \uu0.l_count_4_LC_1_13_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_4_LC_1_13_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \uu0.l_count_4_LC_1_13_7  (
            .in0(N__8949),
            .in1(N__8815),
            .in2(_gnd_net_),
            .in3(N__8157),
            .lcout(\uu0.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21611),
            .ce(N__8729),
            .sr(N__19226));
    defparam \uu0.l_count_5_LC_1_14_0 .C_ON=1'b0;
    defparam \uu0.l_count_5_LC_1_14_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_5_LC_1_14_0 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu0.l_count_5_LC_1_14_0  (
            .in0(N__8950),
            .in1(N__8158),
            .in2(_gnd_net_),
            .in3(N__8132),
            .lcout(\uu0.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21604),
            .ce(N__8730),
            .sr(N__19229));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_15_4 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_15_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_3_LC_1_15_4  (
            .in0(_gnd_net_),
            .in1(N__8160),
            .in2(_gnd_net_),
            .in3(N__8131),
            .lcout(\uu0.un88_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_2_1_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_2_1_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_2_1_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_2_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_2_LC_2_2_0 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_2_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_2_LC_2_2_0 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_2_LC_2_2_0  (
            .in0(N__12377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10400),
            .lcout(\uu2.N_34 ),
            .ltout(\uu2.N_34_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_5_LC_2_2_1 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_5_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_5_LC_2_2_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_5_LC_2_2_1  (
            .in0(N__10700),
            .in1(N__10595),
            .in2(N__8112),
            .in3(N__9398),
            .lcout(\uu2.N_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIDKOL_0_LC_2_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIDKOL_0_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIDKOL_0_LC_2_2_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uu2.w_addr_displaying_RNIDKOL_0_LC_2_2_2  (
            .in0(N__12376),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10399),
            .lcout(\uu2.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_RNIV1P31_4_LC_2_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNIV1P31_4_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNIV1P31_4_LC_2_2_3 .LUT_INIT=16'b1000100000010001;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNIV1P31_4_LC_2_2_3  (
            .in0(N__10699),
            .in1(N__12375),
            .in2(_gnd_net_),
            .in3(N__9397),
            .lcout(\uu2.N_114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_2_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_14_LC_2_2_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_14_LC_2_2_7  (
            .in0(N__10401),
            .in1(N__9042),
            .in2(N__12735),
            .in3(N__9716),
            .lcout(\uu2.mem0.w_data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_2_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_13_LC_2_3_0 .LUT_INIT=16'b0111010011111100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_13_LC_2_3_0  (
            .in0(N__9040),
            .in1(N__9709),
            .in2(N__11166),
            .in3(N__8253),
            .lcout(\uu2.mem0.N_31_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_3_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_15_LC_2_3_1 .LUT_INIT=16'b0000000010001100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_15_LC_2_3_1  (
            .in0(N__11255),
            .in1(N__9038),
            .in2(N__10335),
            .in3(N__10435),
            .lcout(),
            .ltout(\uu2.mem0.N_61_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_2_3_2 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_9_LC_2_3_2 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_9_LC_2_3_2  (
            .in0(N__9714),
            .in1(N__13266),
            .in2(N__8289),
            .in3(N__8268),
            .lcout(\uu2.mem0.w_data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_2_3_3 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_12_LC_2_3_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_12_LC_2_3_3  (
            .in0(N__9710),
            .in1(N__9039),
            .in2(N__11331),
            .in3(N__10436),
            .lcout(\uu2.mem0.w_data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIPAN5U_3_LC_2_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIPAN5U_3_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIPAN5U_3_LC_2_3_4 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \uu2.w_addr_displaying_RNIPAN5U_3_LC_2_3_4  (
            .in0(N__8274),
            .in1(N__10857),
            .in2(N__9423),
            .in3(N__10719),
            .lcout(\uu2.bitmap_pmux ),
            .ltout(\uu2.bitmap_pmux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_2_3_5 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_11_LC_2_3_5 .LUT_INIT=16'b1111101011101110;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_11_LC_2_3_5  (
            .in0(N__8235),
            .in1(N__12783),
            .in2(N__8262),
            .in3(N__9715),
            .lcout(\uu2.mem0.w_data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_2_3_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_16_LC_2_3_6 .LUT_INIT=16'b1010000000100000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_16_LC_2_3_6  (
            .in0(N__9037),
            .in1(N__10324),
            .in2(N__8252),
            .in3(N__11254),
            .lcout(\uu2.mem0.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_2_3_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_8_LC_2_3_7 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_8_LC_2_3_7  (
            .in0(N__11283),
            .in1(N__10437),
            .in2(N__9717),
            .in3(N__9041),
            .lcout(\uu2.mem0.w_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_4_0 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_4_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_4__un404_ci_LC_2_4_0  (
            .in0(N__8569),
            .in1(N__8322),
            .in2(N__8356),
            .in3(N__8611),
            .lcout(\uu2.un404_ci ),
            .ltout(\uu2.un404_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_8_LC_2_4_1 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_8_LC_2_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_8_LC_2_4_1 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_8_LC_2_4_1  (
            .in0(N__8421),
            .in1(N__8432),
            .in2(N__8439),
            .in3(N__8391),
            .lcout(\uu2.r_addrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21665),
            .ce(N__8334),
            .sr(N__19202));
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_4_2 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_4_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_6__un426_ci_3_LC_2_4_2  (
            .in0(_gnd_net_),
            .in1(N__8464),
            .in2(_gnd_net_),
            .in3(N__8532),
            .lcout(\uu2.vbuf_raddr.un426_ci_3 ),
            .ltout(\uu2.vbuf_raddr.un426_ci_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_7_LC_2_4_3 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_7_LC_2_4_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_7_LC_2_4_3 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_7_LC_2_4_3  (
            .in0(N__8380),
            .in1(N__8408),
            .in2(N__8415),
            .in3(N__8497),
            .lcout(\uu2.r_addrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21665),
            .ce(N__8334),
            .sr(N__19202));
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_4_4 .C_ON=1'b0;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu2.vbuf_raddr.counter_gen_label_8__un448_ci_0_LC_2_4_4  (
            .in0(_gnd_net_),
            .in1(N__8407),
            .in2(_gnd_net_),
            .in3(N__8379),
            .lcout(\uu2.vbuf_raddr.un448_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_addr_esr_6_LC_2_4_5 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_6_LC_2_4_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_6_LC_2_4_5 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.r_addr_esr_6_LC_2_4_5  (
            .in0(N__8533),
            .in1(N__8381),
            .in2(N__8471),
            .in3(N__8496),
            .lcout(\uu2.r_addrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21665),
            .ce(N__8334),
            .sr(N__19202));
    defparam \uu2.r_addr_esr_3_LC_2_4_6 .C_ON=1'b0;
    defparam \uu2.r_addr_esr_3_LC_2_4_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_esr_3_LC_2_4_6 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_esr_3_LC_2_4_6  (
            .in0(N__8570),
            .in1(N__8323),
            .in2(N__8357),
            .in3(N__8612),
            .lcout(\uu2.r_addrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21665),
            .ce(N__8334),
            .sr(N__19202));
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_5_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNINBDQ_1_LC_2_5_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.trig_rd_det_RNINBDQ_1_LC_2_5_2  (
            .in0(_gnd_net_),
            .in1(N__10121),
            .in2(_gnd_net_),
            .in3(N__19284),
            .lcout(\uu2.trig_rd_is_det_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_4_LC_2_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_4_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_4_LC_2_6_1 .LUT_INIT=16'b0010000110101010;
    LogicCell40 \uu2.w_addr_user_4_LC_2_6_1  (
            .in0(N__12921),
            .in1(N__14076),
            .in2(N__12885),
            .in3(N__13990),
            .lcout(\uu2.w_addr_userZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_4C_net ),
            .ce(),
            .sr(N__19167));
    defparam \uu2.r_addr_2_LC_2_7_0 .C_ON=1'b0;
    defparam \uu2.r_addr_2_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_2_LC_2_7_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu2.r_addr_2_LC_2_7_0  (
            .in0(N__10114),
            .in1(N__8607),
            .in2(N__8324),
            .in3(N__8565),
            .lcout(\uu2.r_addrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21647),
            .ce(),
            .sr(N__19200));
    defparam \uu2.r_addr_4_LC_2_7_5 .C_ON=1'b0;
    defparam \uu2.r_addr_4_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_4_LC_2_7_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_4_LC_2_7_5  (
            .in0(N__8525),
            .in1(N__8498),
            .in2(_gnd_net_),
            .in3(N__10115),
            .lcout(\uu2.r_addrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21647),
            .ce(),
            .sr(N__19200));
    defparam \uu0.sec_clk_LC_2_7_6 .C_ON=1'b0;
    defparam \uu0.sec_clk_LC_2_7_6 .SEQ_MODE=4'b1010;
    defparam \uu0.sec_clk_LC_2_7_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu0.sec_clk_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__13915),
            .in2(_gnd_net_),
            .in3(N__8816),
            .lcout(o_One_Sec_Pulse),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21647),
            .ce(),
            .sr(N__19200));
    defparam \uu2.r_addr_0_LC_2_8_1 .C_ON=1'b0;
    defparam \uu2.r_addr_0_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_0_LC_2_8_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.r_addr_0_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__8605),
            .in2(_gnd_net_),
            .in3(N__10116),
            .lcout(\uu2.r_addrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21642),
            .ce(),
            .sr(N__19199));
    defparam \uu2.r_addr_1_LC_2_8_5 .C_ON=1'b0;
    defparam \uu2.r_addr_1_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_1_LC_2_8_5 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.r_addr_1_LC_2_8_5  (
            .in0(N__8564),
            .in1(N__8606),
            .in2(_gnd_net_),
            .in3(N__10117),
            .lcout(\uu2.r_addrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21642),
            .ce(),
            .sr(N__19199));
    defparam \uu0.l_count_7_LC_2_9_7 .C_ON=1'b0;
    defparam \uu0.l_count_7_LC_2_9_7 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_7_LC_2_9_7 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_7_LC_2_9_7  (
            .in0(N__8952),
            .in1(N__8802),
            .in2(N__9057),
            .in3(N__8674),
            .lcout(\uu0.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21633),
            .ce(N__8724),
            .sr(N__19219));
    defparam \uu2.r_addr_5_LC_2_10_0 .C_ON=1'b0;
    defparam \uu2.r_addr_5_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_addr_5_LC_2_10_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \uu2.r_addr_5_LC_2_10_0  (
            .in0(N__8534),
            .in1(N__8499),
            .in2(N__10122),
            .in3(N__8460),
            .lcout(\uu2.r_addrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu2.trig_rd_det_0_LC_2_10_1 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_0_LC_2_10_1 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_0_LC_2_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_0_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__13860),
            .in2(_gnd_net_),
            .in3(N__10898),
            .lcout(\uu2.trig_rd_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu2.trig_rd_det_1_LC_2_10_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_1_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \uu2.trig_rd_det_1_LC_2_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.trig_rd_det_1_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10136),
            .lcout(\uu2.trig_rd_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu2.vram_rd_clk_LC_2_10_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_LC_2_10_3 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_LC_2_10_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.vram_rd_clk_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__13861),
            .in2(_gnd_net_),
            .in3(N__8997),
            .lcout(\uu2.vram_rd_clkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu2.l_count_5_LC_2_10_4 .C_ON=1'b0;
    defparam \uu2.l_count_5_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_5_LC_2_10_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \uu2.l_count_5_LC_2_10_4  (
            .in0(N__10027),
            .in1(N__10061),
            .in2(_gnd_net_),
            .in3(N__9269),
            .lcout(\uu2.l_countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu2.l_count_6_LC_2_10_5 .C_ON=1'b0;
    defparam \uu2.l_count_6_LC_2_10_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_6_LC_2_10_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \uu2.l_count_6_LC_2_10_5  (
            .in0(N__9268),
            .in1(N__10003),
            .in2(_gnd_net_),
            .in3(N__9221),
            .lcout(\uu2.l_countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21624),
            .ce(),
            .sr(N__19201));
    defparam \uu0.l_count_17_LC_2_11_0 .C_ON=1'b0;
    defparam \uu0.l_count_17_LC_2_11_0 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_17_LC_2_11_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \uu0.l_count_17_LC_2_11_0  (
            .in0(N__8835),
            .in1(N__8889),
            .in2(N__8658),
            .in3(N__8853),
            .lcout(\uu0.l_countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21617),
            .ce(N__8728),
            .sr(N__19223));
    defparam \uu0.l_count_16_LC_2_11_1 .C_ON=1'b0;
    defparam \uu0.l_count_16_LC_2_11_1 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_16_LC_2_11_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \uu0.l_count_16_LC_2_11_1  (
            .in0(N__8852),
            .in1(N__8801),
            .in2(N__8898),
            .in3(N__8834),
            .lcout(\uu0.l_countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21617),
            .ce(N__8728),
            .sr(N__19223));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_10__un132_ci_8_LC_2_11_2  (
            .in0(N__8936),
            .in1(N__9086),
            .in2(N__9122),
            .in3(N__8676),
            .lcout(\uu0.un110_ci ),
            .ltout(\uu0.un110_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_18__un220_ci_LC_2_11_3  (
            .in0(N__8851),
            .in1(N__8653),
            .in2(N__8838),
            .in3(N__8833),
            .lcout(),
            .ltout(\uu0.un220_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.l_count_18_LC_2_11_4 .C_ON=1'b0;
    defparam \uu0.l_count_18_LC_2_11_4 .SEQ_MODE=4'b1010;
    defparam \uu0.l_count_18_LC_2_11_4 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uu0.l_count_18_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__8800),
            .in2(N__8745),
            .in3(N__8742),
            .lcout(\uu0.l_countZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21617),
            .ce(N__8728),
            .sr(N__19223));
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_6 .C_ON=1'b0;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \uu0.l_count_RNIRLTJ1_17_LC_2_11_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uu0.l_count_RNIRLTJ1_17_LC_2_11_6  (
            .in0(N__8693),
            .in1(N__8675),
            .in2(N__8657),
            .in3(N__8638),
            .lcout(\uu0.un4_l_count_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_12_0 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_0_1_LC_2_12_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_0_1_LC_2_12_0  (
            .in0(N__9338),
            .in1(N__9006),
            .in2(N__9186),
            .in3(N__8958),
            .lcout(\uu2.un1_l_count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_12_1 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_9_LC_2_12_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_9_LC_2_12_1  (
            .in0(N__9223),
            .in1(N__10050),
            .in2(N__8978),
            .in3(N__9314),
            .lcout(),
            .ltout(\uu2.un1_l_count_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_RNI9S834_1_LC_2_12_2 .C_ON=1'b0;
    defparam \uu2.l_count_RNI9S834_1_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNI9S834_1_LC_2_12_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.l_count_RNI9S834_1_LC_2_12_2  (
            .in0(N__9184),
            .in1(N__9342),
            .in2(N__9012),
            .in3(N__9005),
            .lcout(\uu2.un1_l_count_2_0 ),
            .ltout(\uu2.un1_l_count_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_4_LC_2_12_3 .C_ON=1'b0;
    defparam \uu2.l_count_4_LC_2_12_3 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_4_LC_2_12_3 .LUT_INIT=16'b0000001100001100;
    LogicCell40 \uu2.l_count_4_LC_2_12_3  (
            .in0(_gnd_net_),
            .in1(N__9267),
            .in2(N__9009),
            .in3(N__10051),
            .lcout(\uu2.l_countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21612),
            .ce(),
            .sr(N__19227));
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_12_4 .C_ON=1'b0;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIFGGK1_3_LC_2_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.l_count_RNIFGGK1_3_LC_2_12_4  (
            .in0(N__9241),
            .in1(N__10028),
            .in2(N__9144),
            .in3(N__9286),
            .lcout(\uu2.un1_l_count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_9_LC_2_12_5 .C_ON=1'b0;
    defparam \uu2.l_count_9_LC_2_12_5 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_9_LC_2_12_5 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uu2.l_count_9_LC_2_12_5  (
            .in0(N__8996),
            .in1(N__9143),
            .in2(N__8979),
            .in3(N__9156),
            .lcout(\uu2.l_countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21612),
            .ce(),
            .sr(N__19227));
    defparam \uu2.l_count_3_LC_2_12_6 .C_ON=1'b0;
    defparam \uu2.l_count_3_LC_2_12_6 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_3_LC_2_12_6 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \uu2.l_count_3_LC_2_12_6  (
            .in0(N__9185),
            .in1(N__8995),
            .in2(N__9294),
            .in3(N__9198),
            .lcout(\uu2.l_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21612),
            .ce(),
            .sr(N__19227));
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_12_7 .C_ON=1'b0;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \uu2.l_count_RNIBCGK1_0_9_LC_2_12_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uu2.l_count_RNIBCGK1_0_9_LC_2_12_7  (
            .in0(N__9222),
            .in1(N__10049),
            .in2(N__8977),
            .in3(N__9313),
            .lcout(\uu2.un1_l_count_1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_7_LC_2_13_0 .C_ON=1'b0;
    defparam \uu2.l_count_7_LC_2_13_0 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_7_LC_2_13_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \uu2.l_count_7_LC_2_13_0  (
            .in0(N__10005),
            .in1(N__9243),
            .in2(N__9270),
            .in3(N__9225),
            .lcout(\uu2.l_countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21605),
            .ce(),
            .sr(N__19230));
    defparam \uu2.l_count_1_LC_2_13_1 .C_ON=1'b0;
    defparam \uu2.l_count_1_LC_2_13_1 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_1_LC_2_13_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \uu2.l_count_1_LC_2_13_1  (
            .in0(N__9341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9318),
            .lcout(\uu2.l_countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21605),
            .ce(),
            .sr(N__19230));
    defparam \uu2.l_count_0_LC_2_13_2 .C_ON=1'b0;
    defparam \uu2.l_count_0_LC_2_13_2 .SEQ_MODE=4'b1010;
    defparam \uu2.l_count_0_LC_2_13_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uu2.l_count_0_LC_2_13_2  (
            .in0(N__9317),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.l_countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21605),
            .ce(),
            .sr(N__19230));
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_13_3 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_13_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_2__un284_ci_LC_2_13_3  (
            .in0(N__9340),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9316),
            .lcout(\uu2.un284_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_13_5 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_4__un306_ci_LC_2_13_5  (
            .in0(N__9339),
            .in1(N__9315),
            .in2(N__9293),
            .in3(N__9179),
            .lcout(\uu2.un306_ci ),
            .ltout(\uu2.un306_ci_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_13_6 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_8__un350_ci_LC_2_13_6  (
            .in0(N__10004),
            .in1(N__9242),
            .in2(N__9228),
            .in3(N__9224),
            .lcout(\uu2.un350_ci ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.l_count_2_LC_2_14_1 .C_ON=1'b0;
    defparam \uu2.l_count_2_LC_2_14_1 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_2_LC_2_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_2_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__9197),
            .in2(_gnd_net_),
            .in3(N__9180),
            .lcout(\uu2.l_countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21599),
            .ce(),
            .sr(N__19232));
    defparam \uu2.l_count_8_LC_2_14_2 .C_ON=1'b0;
    defparam \uu2.l_count_8_LC_2_14_2 .SEQ_MODE=4'b1011;
    defparam \uu2.l_count_8_LC_2_14_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.l_count_8_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(N__9139),
            .in2(_gnd_net_),
            .in3(N__9155),
            .lcout(\uu2.l_countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21599),
            .ce(),
            .sr(N__19232));
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_15_3 .C_ON=1'b0;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uu0.vbuf_count_cntrl1.counter_gen_label_7__un99_ci_0_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__9109),
            .in2(_gnd_net_),
            .in3(N__9090),
            .lcout(\uu0.un99_ci_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIJQOL_2_LC_4_1_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIJQOL_2_LC_4_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIJQOL_2_LC_4_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.w_addr_displaying_RNIJQOL_2_LC_4_1_1  (
            .in0(N__10685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10831),
            .lcout(),
            .ltout(\uu2.w_data_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI37MM2_3_LC_4_1_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI37MM2_3_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI37MM2_3_LC_4_1_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.w_addr_displaying_RNI37MM2_3_LC_4_1_2  (
            .in0(N__9380),
            .in1(N__10573),
            .in2(N__9045),
            .in3(N__10876),
            .lcout(\uu2.w_data_0_a2_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_4_LC_4_1_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_4_LC_4_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_4_LC_4_1_3 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_nesr_4_LC_4_1_3  (
            .in0(N__10686),
            .in1(N__10586),
            .in2(N__10653),
            .in3(N__9381),
            .lcout(\uu2.w_addr_displayingZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_4C_net ),
            .ce(N__9515),
            .sr(N__19174));
    defparam \uu2.w_addr_displaying_nesr_RNI7MSO_4_LC_4_1_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_RNI7MSO_4_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_nesr_RNI7MSO_4_LC_4_1_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_nesr_RNI7MSO_4_LC_4_1_5  (
            .in0(_gnd_net_),
            .in1(N__12358),
            .in2(_gnd_net_),
            .in3(N__9376),
            .lcout(\uu2.bitmap_pmux_u_0_a2_0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIPFLE1_3_LC_4_1_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIPFLE1_3_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIPFLE1_3_LC_4_1_6 .LUT_INIT=16'b0111001010000000;
    LogicCell40 \uu2.w_addr_displaying_RNIPFLE1_3_LC_4_1_6  (
            .in0(N__10379),
            .in1(N__10572),
            .in2(N__9388),
            .in3(N__10684),
            .lcout(\uu2.bitmap_pmux_sn_N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIDKOL_0_0_LC_4_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIDKOL_0_0_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIDKOL_0_0_LC_4_1_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uu2.w_addr_displaying_RNIDKOL_0_0_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(N__12359),
            .in2(_gnd_net_),
            .in3(N__10378),
            .lcout(\uu2.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_RNIC9NT_LC_4_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_RNIC9NT_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_RNIC9NT_LC_4_2_1 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_RNIC9NT_LC_4_2_1  (
            .in0(N__10374),
            .in1(N__12252),
            .in2(_gnd_net_),
            .in3(N__12183),
            .lcout(\uu2.bitmap_pmux_sn_N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI4GV31_2_LC_4_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI4GV31_2_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI4GV31_2_LC_4_2_2 .LUT_INIT=16'b0101100110011010;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI4GV31_2_LC_4_2_2  (
            .in0(N__9474),
            .in1(N__9375),
            .in2(N__12263),
            .in3(N__10377),
            .lcout(\uu2.N_112_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI7JV31_2_LC_4_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI7JV31_2_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI7JV31_2_LC_4_2_3 .LUT_INIT=16'b0000010100001110;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI7JV31_2_LC_4_2_3  (
            .in0(N__10376),
            .in1(N__12253),
            .in2(N__12579),
            .in3(N__9475),
            .lcout(\uu2.bitmap_pmux_sn_N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIGD5V_2_LC_4_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIGD5V_2_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIGD5V_2_LC_4_2_4 .LUT_INIT=16'b1111111001111111;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIGD5V_2_LC_4_2_4  (
            .in0(N__10380),
            .in1(N__12486),
            .in2(N__9477),
            .in3(N__9374),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_u_0_82_tz_tz_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_RNIT30I1_LC_4_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_RNIT30I1_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_RNIT30I1_LC_4_2_5 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_RNIT30I1_LC_4_2_5  (
            .in0(_gnd_net_),
            .in1(N__12257),
            .in2(N__9345),
            .in3(N__12360),
            .lcout(\uu2.N_921_tz_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_2_LC_4_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_2_LC_4_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_2_LC_4_2_6 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uu2.w_addr_displaying_fast_2_LC_4_2_6  (
            .in0(N__9476),
            .in1(N__10636),
            .in2(_gnd_net_),
            .in3(N__10476),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_fast_2C_net ),
            .ce(),
            .sr(N__19173));
    defparam \uu2.w_addr_displaying_fast_RNI245H_2_LC_4_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI245H_2_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI245H_2_LC_4_2_7 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI245H_2_LC_4_2_7  (
            .in0(N__10375),
            .in1(N__12091),
            .in2(_gnd_net_),
            .in3(N__9470),
            .lcout(\uu2.bitmap_pmux_sn_N_54_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_186_LC_4_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_186_LC_4_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_186_LC_4_3_0 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_186_LC_4_3_0  (
            .in0(N__11100),
            .in1(N__11130),
            .in2(N__11062),
            .in3(N__12666),
            .lcout(\uu2.bitmapZ0Z_186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__19171));
    defparam \uu2.bitmap_RNIBG4K_58_LC_4_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIBG4K_58_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIBG4K_58_LC_4_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uu2.bitmap_RNIBG4K_58_LC_4_3_1  (
            .in0(N__9456),
            .in1(N__9450),
            .in2(_gnd_net_),
            .in3(N__10970),
            .lcout(\uu2.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_58_LC_4_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_58_LC_4_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_58_LC_4_3_2 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_58_LC_4_3_2  (
            .in0(N__11102),
            .in1(N__11132),
            .in2(N__11064),
            .in3(N__12668),
            .lcout(\uu2.bitmapZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__19171));
    defparam \uu2.bitmap_93_LC_4_3_3 .C_ON=1'b0;
    defparam \uu2.bitmap_93_LC_4_3_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_93_LC_4_3_3 .LUT_INIT=16'b0010100101111111;
    LogicCell40 \uu2.bitmap_93_LC_4_3_3  (
            .in0(N__12669),
            .in1(N__11060),
            .in2(N__11136),
            .in3(N__11103),
            .lcout(\uu2.bitmapZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__19171));
    defparam \uu2.bitmap_221_LC_4_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_221_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_221_LC_4_3_4 .LUT_INIT=16'b0111111101011011;
    LogicCell40 \uu2.bitmap_221_LC_4_3_4  (
            .in0(N__11101),
            .in1(N__11131),
            .in2(N__11063),
            .in3(N__12667),
            .lcout(\uu2.bitmapZ0Z_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_186C_net ),
            .ce(),
            .sr(N__19171));
    defparam \uu2.bitmap_RNIRETJ1_93_LC_4_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIRETJ1_93_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIRETJ1_93_LC_4_3_5 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \uu2.bitmap_RNIRETJ1_93_LC_4_3_5  (
            .in0(N__12362),
            .in1(N__9444),
            .in2(N__9438),
            .in3(N__10986),
            .lcout(),
            .ltout(\uu2.bitmap_RNIRETJ1Z0Z_93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNIHPJ64_3_LC_4_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNIHPJ64_3_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNIHPJ64_3_LC_4_3_6 .LUT_INIT=16'b0011001100011101;
    LogicCell40 \uu2.w_addr_displaying_RNIHPJ64_3_LC_4_3_6  (
            .in0(N__10212),
            .in1(N__10579),
            .in2(N__9429),
            .in3(N__10426),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_27_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIIU8Q8_72_LC_4_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIIU8Q8_72_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIIU8Q8_72_LC_4_3_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uu2.bitmap_RNIIU8Q8_72_LC_4_3_7  (
            .in0(N__10427),
            .in1(N__12318),
            .in2(N__9426),
            .in3(N__10884),
            .lcout(\uu2.N_404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_4_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_5_LC_4_4_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_5_LC_4_4_0  (
            .in0(N__10316),
            .in1(N__10789),
            .in2(N__12966),
            .in3(N__11250),
            .lcout(\uu2.mem0.N_135 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_4_1 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_6_LC_4_4_1 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_6_LC_4_4_1  (
            .in0(N__11251),
            .in1(N__10317),
            .in2(N__13962),
            .in3(N__12558),
            .lcout(\uu2.mem0.N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_nesr_7_LC_4_4_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_nesr_7_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_nesr_7_LC_4_4_2 .LUT_INIT=16'b1010011010101010;
    LogicCell40 \uu2.w_addr_displaying_nesr_7_LC_4_4_2  (
            .in0(N__12560),
            .in1(N__10793),
            .in2(N__10527),
            .in3(N__10847),
            .lcout(\uu2.w_addr_displayingZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_7C_net ),
            .ce(N__9516),
            .sr(N__19169));
    defparam \uu2.w_addr_displaying_ness_6_LC_4_4_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_6_LC_4_4_3 .SEQ_MODE=4'b1001;
    defparam \uu2.w_addr_displaying_ness_6_LC_4_4_3 .LUT_INIT=16'b1111110011011110;
    LogicCell40 \uu2.w_addr_displaying_ness_6_LC_4_4_3  (
            .in0(N__10848),
            .in1(N__10878),
            .in2(N__10800),
            .in3(N__10524),
            .lcout(\uu2.w_addr_displayingZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_7C_net ),
            .ce(N__9516),
            .sr(N__19169));
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_4_4_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_nesr_7_LC_4_4_4 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_fast_nesr_7_LC_4_4_4  (
            .in0(N__10797),
            .in1(N__10846),
            .in2(N__10526),
            .in3(N__10980),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_nesr_7C_net ),
            .ce(N__9516),
            .sr(N__19169));
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_8_LC_4_4_5 .C_ON=1'b0;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_8_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_w_addr_displaying.result_1_0_o2_8_LC_4_4_5 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \uu2.vbuf_w_addr_displaying.result_1_0_o2_8_LC_4_4_5  (
            .in0(N__10845),
            .in1(N__10517),
            .in2(N__10799),
            .in3(N__12559),
            .lcout(\uu2.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI0ES07_5_LC_4_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI0ES07_5_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI0ES07_5_LC_4_4_6 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \uu2.w_addr_displaying_RNI0ES07_5_LC_4_4_6  (
            .in0(N__10877),
            .in1(N__10844),
            .in2(N__10525),
            .in3(N__9685),
            .lcout(\uu2.w_addr_displaying_RNI0ES07Z0Z_5 ),
            .ltout(\uu2.w_addr_displaying_RNI0ES07Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI47N27_5_LC_4_4_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI47N27_5_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI47N27_5_LC_4_4_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uu2.w_addr_displaying_RNI47N27_5_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9519),
            .in3(N__15584),
            .lcout(\uu2.N_32_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_0 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_7_LC_4_5_0  (
            .in0(N__12200),
            .in1(N__9661),
            .in2(N__10333),
            .in3(N__11252),
            .lcout(\uu2.mem0.N_133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNI20V6_8_LC_4_5_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNI20V6_8_LC_4_5_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNI20V6_8_LC_4_5_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNI20V6_8_LC_4_5_1  (
            .in0(N__13954),
            .in1(N__9632),
            .in2(N__9663),
            .in3(N__9564),
            .lcout(\uu2.w_addr_user_3_i_a2_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_8_LC_4_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_8_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_8_LC_4_5_2 .LUT_INIT=16'b0000000010100110;
    LogicCell40 \uu2.w_addr_user_nesr_8_LC_4_5_2  (
            .in0(N__9662),
            .in1(N__13955),
            .in2(N__14030),
            .in3(N__14063),
            .lcout(\uu2.w_addr_userZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12815),
            .sr(N__19168));
    defparam \uu2.w_addr_user_nesr_2_LC_4_5_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_2_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_2_LC_4_5_3 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \uu2.w_addr_user_nesr_2_LC_4_5_3  (
            .in0(N__14060),
            .in1(N__9636),
            .in2(N__9857),
            .in3(N__9566),
            .lcout(\uu2.w_addr_userZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12815),
            .sr(N__19168));
    defparam \uu2.w_addr_user_nesr_0_LC_4_5_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_0_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_0_LC_4_5_4 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \uu2.w_addr_user_nesr_0_LC_4_5_4  (
            .in0(N__9567),
            .in1(N__9815),
            .in2(N__12971),
            .in3(N__14059),
            .lcout(\uu2.w_addr_userZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12815),
            .sr(N__19168));
    defparam \uu2.w_addr_user_nesr_6_LC_4_5_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_6_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_6_LC_4_5_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \uu2.w_addr_user_nesr_6_LC_4_5_5  (
            .in0(N__14062),
            .in1(N__14023),
            .in2(N__9870),
            .in3(N__9816),
            .lcout(\uu2.w_addr_userZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12815),
            .sr(N__19168));
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_4_5_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_4_5_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_3_LC_4_5_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_3_LC_4_5_6  (
            .in0(N__9565),
            .in1(N__9798),
            .in2(N__9639),
            .in3(N__9850),
            .lcout(),
            .ltout(\uu2.N_161_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_3_LC_4_5_7 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_3_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_3_LC_4_5_7 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \uu2.w_addr_user_nesr_3_LC_4_5_7  (
            .in0(N__14061),
            .in1(_gnd_net_),
            .in2(N__9645),
            .in3(N__12873),
            .lcout(\uu2.w_addr_userZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_8C_net ),
            .ce(N__12815),
            .sr(N__19168));
    defparam \uu2.un28_w_addr_user_i_0_o2_LC_4_6_0 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_o2_LC_4_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_o2_LC_4_6_0 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \uu2.un28_w_addr_user_i_0_o2_LC_4_6_0  (
            .in0(N__11276),
            .in1(N__11007),
            .in2(N__11019),
            .in3(N__11206),
            .lcout(\uu2.N_101 ),
            .ltout(\uu2.N_101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIE43C7_6_LC_4_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIE43C7_6_LC_4_6_1 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIE43C7_6_LC_4_6_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \uu2.w_addr_user_nesr_RNIE43C7_6_LC_4_6_1  (
            .in0(N__12967),
            .in1(N__9814),
            .in2(N__9642),
            .in3(N__10275),
            .lcout(\uu2.un28_w_addr_user_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_4_6_3 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIFBD5_3_LC_4_6_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIFBD5_3_LC_4_6_3  (
            .in0(N__9797),
            .in1(N__9846),
            .in2(N__9638),
            .in3(N__9574),
            .lcout(\uu2.N_106 ),
            .ltout(\uu2.N_106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_4_6_4 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNO_0_6_LC_4_6_4 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \uu2.w_addr_user_nesr_RNO_0_6_LC_4_6_4  (
            .in0(N__12962),
            .in1(N__12849),
            .in2(N__9873),
            .in3(N__12912),
            .lcout(\uu2.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_4_6_5 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNINJD5_3_LC_4_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.w_addr_user_nesr_RNINJD5_3_LC_4_6_5  (
            .in0(N__12911),
            .in1(N__9795),
            .in2(N__12852),
            .in3(N__9845),
            .lcout(),
            .ltout(\uu2.w_addr_user_3_i_a2_2_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIPJCC_3_LC_4_6_6 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIPJCC_3_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIPJCC_3_LC_4_6_6 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \uu2.w_addr_user_nesr_RNIPJCC_3_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__9825),
            .in2(N__9819),
            .in3(_gnd_net_),
            .lcout(\uu2.N_230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_6_7 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_2_LC_4_6_7 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_2_LC_4_6_7  (
            .in0(N__11207),
            .in1(N__9796),
            .in2(N__10334),
            .in3(N__10605),
            .lcout(\uu2.mem0.N_138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_RNISDHD_LC_4_7_0 .C_ON=1'b0;
    defparam \uu0.sec_clkD_RNISDHD_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \uu0.sec_clkD_RNISDHD_LC_4_7_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu0.sec_clkD_RNISDHD_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__12691),
            .in2(_gnd_net_),
            .in3(N__13916),
            .lcout(oneSecStrb),
            .ltout(oneSecStrb_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.rdy_LC_4_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.rdy_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.rdy_LC_4_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dispString.rdy_LC_4_7_1  (
            .in0(N__13090),
            .in1(N__14362),
            .in2(N__9762),
            .in3(N__14480),
            .lcout(L3_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21634),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_wr_en_0_i_LC_4_7_2 .C_ON=1'b0;
    defparam \uu2.vram_wr_en_0_i_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_wr_en_0_i_LC_4_7_2 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \uu2.vram_wr_en_0_i_LC_4_7_2  (
            .in0(N__9758),
            .in1(N__10274),
            .in2(_gnd_net_),
            .in3(N__11204),
            .lcout(\uu2.vram_wr_en_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu0.sec_clkD_LC_4_7_3 .C_ON=1'b0;
    defparam \uu0.sec_clkD_LC_4_7_3 .SEQ_MODE=4'b1000;
    defparam \uu0.sec_clkD_LC_4_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu0.sec_clkD_LC_4_7_3  (
            .in0(N__13917),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(uu0_sec_clkD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21634),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un4_w_user_data_rdy_i_o2_0_LC_4_7_4 .C_ON=1'b0;
    defparam \uu2.un4_w_user_data_rdy_i_o2_0_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \uu2.un4_w_user_data_rdy_i_o2_0_LC_4_7_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \uu2.un4_w_user_data_rdy_i_o2_0_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__10273),
            .in2(_gnd_net_),
            .in3(N__11203),
            .lcout(\uu2.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_7_6 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_10_LC_4_7_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_10_LC_4_7_6  (
            .in0(N__10297),
            .in1(N__11304),
            .in2(_gnd_net_),
            .in3(N__11205),
            .lcout(\uu2.mem0.N_54_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_0_LC_4_8_0 .C_ON=1'b0;
    defparam \uu2.r_data_reg_0_LC_4_8_0 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_0_LC_4_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_0_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9969),
            .lcout(vbuf_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_1_LC_4_8_1 .C_ON=1'b0;
    defparam \uu2.r_data_reg_1_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_1_LC_4_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_1_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9957),
            .lcout(vbuf_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_2_LC_4_8_2 .C_ON=1'b0;
    defparam \uu2.r_data_reg_2_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_2_LC_4_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_2_LC_4_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9945),
            .lcout(vbuf_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_3_LC_4_8_3 .C_ON=1'b0;
    defparam \uu2.r_data_reg_3_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_3_LC_4_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_3_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9933),
            .lcout(vbuf_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_4_LC_4_8_4 .C_ON=1'b0;
    defparam \uu2.r_data_reg_4_LC_4_8_4 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_4_LC_4_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_4_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9921),
            .lcout(vbuf_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_5_LC_4_8_5 .C_ON=1'b0;
    defparam \uu2.r_data_reg_5_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_5_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_5_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9909),
            .lcout(vbuf_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_6_LC_4_8_6 .C_ON=1'b0;
    defparam \uu2.r_data_reg_6_LC_4_8_6 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_6_LC_4_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_6_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9897),
            .lcout(vbuf_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \uu2.r_data_reg_7_LC_4_8_7 .C_ON=1'b0;
    defparam \uu2.r_data_reg_7_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_reg_7_LC_4_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.r_data_reg_7_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9885),
            .lcout(vbuf_tx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.r_data_reg_0C_net ),
            .ce(N__11343),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_1_LC_4_9_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_1_LC_4_9_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_1_LC_4_9_0 .LUT_INIT=16'b1111110111001110;
    LogicCell40 \buart.Z_tx.bitcount_1_LC_4_9_0  (
            .in0(N__11543),
            .in1(N__13217),
            .in2(N__11523),
            .in3(N__11480),
            .lcout(\buart.Z_tx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(N__19224));
    defparam \buart.Z_tx.bitcount_0_LC_4_9_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_0_LC_4_9_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_0_LC_4_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.bitcount_0_LC_4_9_1  (
            .in0(N__13216),
            .in1(N__11519),
            .in2(_gnd_net_),
            .in3(N__11542),
            .lcout(\buart.Z_tx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(N__19224));
    defparam \buart.Z_tx.bitcount_3_LC_4_9_2 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_3_LC_4_9_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_3_LC_4_9_2 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \buart.Z_tx.bitcount_3_LC_4_9_2  (
            .in0(N__11544),
            .in1(N__11580),
            .in2(N__13218),
            .in3(N__11457),
            .lcout(\buart.Z_tx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(N__19224));
    defparam \buart.Z_tx.bitcount_2_LC_4_9_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_2_LC_4_9_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.bitcount_2_LC_4_9_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \buart.Z_tx.bitcount_2_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__13212),
            .in2(_gnd_net_),
            .in3(N__11586),
            .lcout(\buart.Z_tx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21618),
            .ce(),
            .sr(N__19224));
    defparam \buart.Z_rx.bitcount_es_1_LC_4_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_1_LC_4_10_0 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_1_LC_4_10_0 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_es_1_LC_4_10_0  (
            .in0(N__10182),
            .in1(N__12053),
            .in2(N__11685),
            .in3(N__11820),
            .lcout(\buart.Z_rx.bitcountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21613),
            .ce(N__12025),
            .sr(N__19228));
    defparam \buart.Z_rx.bitcount_es_2_LC_4_10_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_2_LC_4_10_1 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_2_LC_4_10_1 .LUT_INIT=16'b0101001101011100;
    LogicCell40 \buart.Z_rx.bitcount_es_2_LC_4_10_1  (
            .in0(N__11819),
            .in1(N__10173),
            .in2(N__12060),
            .in3(N__11628),
            .lcout(\buart.Z_rx.bitcountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21613),
            .ce(N__12025),
            .sr(N__19228));
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_10_2 .C_ON=1'b0;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \uu2.trig_rd_det_RNIJIIO_1_LC_4_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.trig_rd_det_RNIJIIO_1_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__10146),
            .in2(_gnd_net_),
            .in3(N__10137),
            .lcout(\uu2.trig_rd_is_det ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_10_4 .C_ON=1'b0;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_10_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uu2.vbuf_count.counter_gen_label_6__un328_ci_3_LC_4_10_4  (
            .in0(N__10062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10029),
            .lcout(\uu2.vbuf_count.un328_ci_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_11_0 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_c_0_LC_4_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_c_0_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__11867),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\buart.Z_rx.bitcount_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_11_1 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_0_THRU_LUT4_0_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__11681),
            .in2(_gnd_net_),
            .in3(N__10176),
            .lcout(\buart.Z_rx.bitcount_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_0 ),
            .carryout(\buart.Z_rx.bitcount_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_11_2 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_1_THRU_LUT4_0_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__11627),
            .in2(_gnd_net_),
            .in3(N__10167),
            .lcout(\buart.Z_rx.bitcount_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_1 ),
            .carryout(\buart.Z_rx.bitcount_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_11_3 .C_ON=1'b1;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.bitcount_cry_2_THRU_LUT4_0_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__11711),
            .in2(_gnd_net_),
            .in3(N__10164),
            .lcout(\buart.Z_rx.bitcount_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.bitcount_cry_2 ),
            .carryout(\buart.Z_rx.bitcount_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_4_LC_4_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_4_LC_4_11_4 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_4_LC_4_11_4 .LUT_INIT=16'b0010011101110010;
    LogicCell40 \buart.Z_rx.bitcount_es_4_LC_4_11_4  (
            .in0(N__12057),
            .in1(N__11827),
            .in2(N__11655),
            .in3(N__10161),
            .lcout(\buart.Z_rx.bitcountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21606),
            .ce(N__12030),
            .sr(N__19231));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_12_0 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_c_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__11940),
            .in2(N__11772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_12_1 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_LUT4_0_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__11921),
            .in2(_gnd_net_),
            .in3(N__10158),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_1 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_12_2 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_12_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_3_LC_4_12_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_3_LC_4_12_2  (
            .in0(N__11821),
            .in1(N__11970),
            .in2(_gnd_net_),
            .in3(N__10155),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_2 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .clk(N__21600),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_12_3 .C_ON=1'b1;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_LUT4_0_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__11987),
            .in2(_gnd_net_),
            .in3(N__10152),
            .lcout(\buart.Z_rx.Z_baudgen.un5_counter_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\buart.Z_rx.Z_baudgen.un5_counter_cry_3 ),
            .carryout(\buart.Z_rx.Z_baudgen.un5_counter_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_12_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_5_LC_4_12_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_5_LC_4_12_4  (
            .in0(N__11823),
            .in1(N__11898),
            .in2(N__11958),
            .in3(N__10149),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21600),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_12_6 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_2_LC_4_12_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_2_LC_4_12_6  (
            .in0(N__11822),
            .in1(N__10227),
            .in2(N__11925),
            .in3(N__11899),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21600),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_194_LC_5_1_0 .C_ON=1'b0;
    defparam \uu2.bitmap_194_LC_5_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_194_LC_5_1_0 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \uu2.bitmap_194_LC_5_1_0  (
            .in0(N__12437),
            .in1(N__13670),
            .in2(N__13420),
            .in3(N__13634),
            .lcout(\uu2.bitmapZ0Z_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.bitmap_RNII0BN_69_LC_5_1_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNII0BN_69_LC_5_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNII0BN_69_LC_5_1_1 .LUT_INIT=16'b0001100100111011;
    LogicCell40 \uu2.bitmap_RNII0BN_69_LC_5_1_1  (
            .in0(N__12479),
            .in1(N__10979),
            .in2(N__10203),
            .in3(N__10188),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_25_i_m2_am_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIG91I1_66_LC_5_1_2 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIG91I1_66_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIG91I1_66_LC_5_1_2 .LUT_INIT=16'b0000111110101100;
    LogicCell40 \uu2.bitmap_RNIG91I1_66_LC_5_1_2  (
            .in0(N__10221),
            .in1(N__10194),
            .in2(N__10215),
            .in3(N__12361),
            .lcout(\uu2.bitmap_RNIG91I1Z0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_34_LC_5_1_3 .C_ON=1'b0;
    defparam \uu2.bitmap_34_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_34_LC_5_1_3 .LUT_INIT=16'b1111011101101101;
    LogicCell40 \uu2.bitmap_34_LC_5_1_3  (
            .in0(N__13636),
            .in1(N__13414),
            .in2(N__13679),
            .in3(N__12439),
            .lcout(\uu2.bitmapZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.bitmap_69_LC_5_1_4 .C_ON=1'b0;
    defparam \uu2.bitmap_69_LC_5_1_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_69_LC_5_1_4 .LUT_INIT=16'b0101101100110111;
    LogicCell40 \uu2.bitmap_69_LC_5_1_4  (
            .in0(N__12441),
            .in1(N__13678),
            .in2(N__13422),
            .in3(N__13638),
            .lcout(\uu2.bitmapZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.bitmap_66_LC_5_1_5 .C_ON=1'b0;
    defparam \uu2.bitmap_66_LC_5_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_66_LC_5_1_5 .LUT_INIT=16'b0001000000111101;
    LogicCell40 \uu2.bitmap_66_LC_5_1_5  (
            .in0(N__13637),
            .in1(N__13415),
            .in2(N__13680),
            .in3(N__12440),
            .lcout(\uu2.bitmapZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.bitmap_197_LC_5_1_6 .C_ON=1'b0;
    defparam \uu2.bitmap_197_LC_5_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_197_LC_5_1_6 .LUT_INIT=16'b0111111100111101;
    LogicCell40 \uu2.bitmap_197_LC_5_1_6  (
            .in0(N__12438),
            .in1(N__13671),
            .in2(N__13421),
            .in3(N__13635),
            .lcout(\uu2.bitmapZ0Z_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.w_addr_displaying_fast_0_LC_5_1_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_0_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_0_LC_5_1_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \uu2.w_addr_displaying_fast_0_LC_5_1_7  (
            .in0(N__10485),
            .in1(_gnd_net_),
            .in2(N__12488),
            .in3(_gnd_net_),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_194C_net ),
            .ce(),
            .sr(N__19177));
    defparam \uu2.w_addr_displaying_3_rep1_LC_5_2_0 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_LC_5_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_rep1_LC_5_2_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_LC_5_2_0  (
            .in0(N__10695),
            .in1(N__10483),
            .in2(N__10648),
            .in3(N__12262),
            .lcout(\uu2.w_addr_displaying_3_repZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_2_LC_5_2_1 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_2_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_2_LC_5_2_1 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uu2.w_addr_displaying_2_LC_5_2_1  (
            .in0(N__10479),
            .in1(N__10637),
            .in2(_gnd_net_),
            .in3(N__10697),
            .lcout(\uu2.w_addr_displayingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_fast_3_LC_5_2_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_3_LC_5_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_fast_3_LC_5_2_2 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \uu2.w_addr_displaying_fast_3_LC_5_2_2  (
            .in0(N__10696),
            .in1(N__10484),
            .in2(N__10649),
            .in3(N__12095),
            .lcout(\uu2.w_addr_displaying_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_3_LC_5_2_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_LC_5_2_3 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_3_LC_5_2_3 .LUT_INIT=16'b1111000001111000;
    LogicCell40 \uu2.w_addr_displaying_3_LC_5_2_3  (
            .in0(N__10482),
            .in1(N__10698),
            .in2(N__10596),
            .in3(N__10638),
            .lcout(\uu2.w_addr_displayingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_0_LC_5_2_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_0_LC_5_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_0_LC_5_2_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uu2.w_addr_displaying_0_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__10477),
            .in2(_gnd_net_),
            .in3(N__12374),
            .lcout(\uu2.w_addr_displayingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_8_LC_5_2_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_8_LC_5_2_5 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_8_LC_5_2_5 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uu2.w_addr_displaying_8_LC_5_2_5  (
            .in0(N__10481),
            .in1(N__10539),
            .in2(_gnd_net_),
            .in3(N__12195),
            .lcout(\uu2.w_addr_displayingZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_5_LC_5_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_5_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_5_LC_5_2_6 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \uu2.w_addr_displaying_5_LC_5_2_6  (
            .in0(N__10513),
            .in1(N__10480),
            .in2(_gnd_net_),
            .in3(N__10843),
            .lcout(\uu2.w_addr_displayingZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.w_addr_displaying_1_LC_5_2_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_1_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_displaying_1_LC_5_2_7 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \uu2.w_addr_displaying_1_LC_5_2_7  (
            .in0(N__10478),
            .in1(N__10425),
            .in2(_gnd_net_),
            .in3(N__10391),
            .lcout(\uu2.w_addr_displayingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_displaying_3_rep1C_net ),
            .ce(),
            .sr(N__19175));
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_0 .C_ON=1'b0;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_0 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \uu2.mem0.ram512X8_inst_RNO_4_LC_5_3_0  (
            .in0(N__10332),
            .in1(N__10830),
            .in2(N__11253),
            .in3(N__12850),
            .lcout(\uu2.mem0.N_136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIFJI02_212_LC_5_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIFJI02_212_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIFJI02_212_LC_5_3_1 .LUT_INIT=16'b0010001011111100;
    LogicCell40 \uu2.bitmap_RNIFJI02_212_LC_5_3_1  (
            .in0(N__13689),
            .in1(N__12547),
            .in2(N__13791),
            .in3(N__12447),
            .lcout(\uu2.bitmap_RNIFJI02Z0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNI6J081_6_LC_5_3_2 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI6J081_6_LC_5_3_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI6J081_6_LC_5_3_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI6J081_6_LC_5_3_2  (
            .in0(N__12191),
            .in1(_gnd_net_),
            .in2(N__12567),
            .in3(N__10783),
            .lcout(\uu2.N_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_0_6_LC_5_3_3 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_0_6_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_0_6_LC_5_3_3 .LUT_INIT=16'b0000011101110000;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI12TI1_0_6_LC_5_3_3  (
            .in0(N__10829),
            .in1(N__10788),
            .in2(N__12581),
            .in3(N__12194),
            .lcout(\uu2.bitmap_pmux_u_0_83_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_1_6_LC_5_3_4 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_1_6_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_1_6_LC_5_3_4 .LUT_INIT=16'b0000011001000010;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI12TI1_1_6_LC_5_3_4  (
            .in0(N__12192),
            .in1(N__12571),
            .in2(N__10798),
            .in3(N__10828),
            .lcout(\uu2.bitmap_pmux_sn_N_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_6_LC_5_3_5 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_6_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_ness_RNI12TI1_6_LC_5_3_5 .LUT_INIT=16'b1111011101110111;
    LogicCell40 \uu2.w_addr_displaying_ness_RNI12TI1_6_LC_5_3_5  (
            .in0(N__10827),
            .in1(N__10787),
            .in2(N__12582),
            .in3(N__12193),
            .lcout(),
            .ltout(\uu2.N_100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNI3OPR5_2_LC_5_3_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNI3OPR5_2_LC_5_3_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNI3OPR5_2_LC_5_3_6 .LUT_INIT=16'b1010111000001100;
    LogicCell40 \uu2.w_addr_displaying_fast_RNI3OPR5_2_LC_5_3_6  (
            .in0(N__10752),
            .in1(N__10746),
            .in2(N__10740),
            .in3(N__10737),
            .lcout(),
            .ltout(\uu2.N_923_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_RNI8ND5G_3_LC_5_3_7 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_RNI8ND5G_3_LC_5_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_RNI8ND5G_3_LC_5_3_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \uu2.w_addr_displaying_RNI8ND5G_3_LC_5_3_7  (
            .in0(N__10731),
            .in1(N__10932),
            .in2(N__10722),
            .in3(N__12279),
            .lcout(\uu2.w_addr_displaying_RNI8ND5GZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_314_LC_5_4_0 .C_ON=1'b0;
    defparam \uu2.bitmap_314_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_314_LC_5_4_0 .LUT_INIT=16'b0001001000100111;
    LogicCell40 \uu2.bitmap_314_LC_5_4_0  (
            .in0(N__11119),
            .in1(N__11049),
            .in2(N__11089),
            .in3(N__12652),
            .lcout(\uu2.bitmapZ0Z_314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__19172));
    defparam \uu2.bitmap_218_LC_5_4_1 .C_ON=1'b0;
    defparam \uu2.bitmap_218_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_218_LC_5_4_1 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \uu2.bitmap_218_LC_5_4_1  (
            .in0(N__12651),
            .in1(N__11079),
            .in2(N__11061),
            .in3(N__11118),
            .lcout(\uu2.bitmapZ0Z_218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__19172));
    defparam \uu2.bitmap_90_LC_5_4_2 .C_ON=1'b0;
    defparam \uu2.bitmap_90_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_90_LC_5_4_2 .LUT_INIT=16'b0001010000110101;
    LogicCell40 \uu2.bitmap_90_LC_5_4_2  (
            .in0(N__11120),
            .in1(N__11050),
            .in2(N__11090),
            .in3(N__12653),
            .lcout(\uu2.bitmapZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_314C_net ),
            .ce(),
            .sr(N__19172));
    defparam \uu2.bitmap_RNI6H8O_90_LC_5_4_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI6H8O_90_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI6H8O_90_LC_5_4_3 .LUT_INIT=16'b0100010101100111;
    LogicCell40 \uu2.bitmap_RNI6H8O_90_LC_5_4_3  (
            .in0(N__10978),
            .in1(N__12489),
            .in2(N__11001),
            .in3(N__10992),
            .lcout(\uu2.bitmap_pmux_25_i_m2_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIU0UJ_314_LC_5_4_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIU0UJ_314_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIU0UJ_314_LC_5_4_4 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \uu2.bitmap_RNIU0UJ_314_LC_5_4_4  (
            .in0(N__12096),
            .in1(N__10977),
            .in2(_gnd_net_),
            .in3(N__10925),
            .lcout(),
            .ltout(\uu2.bitmap_pmux_21_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIBNS22_180_LC_5_4_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIBNS22_180_LC_5_4_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIBNS22_180_LC_5_4_5 .LUT_INIT=16'b0011111000001110;
    LogicCell40 \uu2.bitmap_RNIBNS22_180_LC_5_4_5  (
            .in0(N__13806),
            .in1(N__12264),
            .in2(N__10950),
            .in3(N__12135),
            .lcout(),
            .ltout(\uu2.N_393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_3_rep1_RNIN52C4_LC_5_4_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_3_rep1_RNIN52C4_LC_5_4_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_3_rep1_RNIN52C4_LC_5_4_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_3_rep1_RNIN52C4_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__10947),
            .in2(N__10935),
            .in3(N__10911),
            .lcout(\uu2.N_397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNI05EB1_314_LC_5_4_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI05EB1_314_LC_5_4_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI05EB1_314_LC_5_4_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uu2.bitmap_RNI05EB1_314_LC_5_4_7  (
            .in0(N__10926),
            .in1(N__12199),
            .in2(_gnd_net_),
            .in3(N__10917),
            .lcout(\uu2.N_131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.r_data_rdy_LC_5_5_1 .C_ON=1'b0;
    defparam \uu2.r_data_rdy_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \uu2.r_data_rdy_LC_5_5_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \uu2.r_data_rdy_LC_5_5_1  (
            .in0(N__13875),
            .in1(N__10905),
            .in2(N__13199),
            .in3(N__19287),
            .lcout(vbuf_tx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21643),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_RNIITTD7_6_LC_5_5_2 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIITTD7_6_LC_5_5_2 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIITTD7_6_LC_5_5_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \uu2.w_addr_user_nesr_RNIITTD7_6_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__15574),
            .in2(_gnd_net_),
            .in3(N__13980),
            .lcout(\uu2.un28_w_addr_user_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_5_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_0_LC_5_5_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_0_LC_5_5_3  (
            .in0(N__18006),
            .in1(N__18046),
            .in2(_gnd_net_),
            .in3(N__19949),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_0_LC_5_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_0_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_0_LC_5_5_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce1.q_0_LC_5_5_4  (
            .in0(N__18047),
            .in1(N__15810),
            .in2(N__11139),
            .in3(N__15843),
            .lcout(\Lab_UT.didp.di_Sones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21643),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIFKHR3_1_LC_5_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIFKHR3_1_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIFKHR3_1_LC_5_5_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIFKHR3_1_LC_5_5_5  (
            .in0(N__17964),
            .in1(N__14571),
            .in2(_gnd_net_),
            .in3(N__17319),
            .lcout(\Lab_UT.sec2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIHMHR3_2_LC_5_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIHMHR3_2_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIHMHR3_2_LC_5_5_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIHMHR3_2_LC_5_5_6  (
            .in0(N__14570),
            .in1(N__16044),
            .in2(_gnd_net_),
            .in3(N__17295),
            .lcout(\Lab_UT.sec2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJOHR3_3_LC_5_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJOHR3_3_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIJOHR3_3_LC_5_5_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIJOHR3_3_LC_5_5_7  (
            .in0(N__15999),
            .in1(N__14572),
            .in2(_gnd_net_),
            .in3(N__17265),
            .lcout(\Lab_UT.sec2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_a2_0_4_LC_5_6_0 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_4_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_4_LC_5_6_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a2_0_4_LC_5_6_0  (
            .in0(N__11303),
            .in1(N__11156),
            .in2(N__12779),
            .in3(N__11321),
            .lcout(\uu2.un28_w_addr_user_i_0_a2_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_6_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \Lab_UT.dispString.cnt_RNIOG7L_2_LC_5_6_1  (
            .in0(N__13079),
            .in1(N__14356),
            .in2(_gnd_net_),
            .in3(N__14483),
            .lcout(\Lab_UT.dispString.un42_dOutP ),
            .ltout(\Lab_UT.dispString.un42_dOutP_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_2_LC_5_6_2 .LUT_INIT=16'b1000100000001000;
    LogicCell40 \Lab_UT.dispString.dOut_2_LC_5_6_2  (
            .in0(N__11355),
            .in1(N__11349),
            .in2(N__11010),
            .in3(N__12636),
            .lcout(L3_tx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21635),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un28_w_addr_user_i_0_a2_0_0_LC_5_6_3 .C_ON=1'b0;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_0_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \uu2.un28_w_addr_user_i_0_a2_0_0_LC_5_6_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uu2.un28_w_addr_user_i_0_a2_0_0_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__12721),
            .in2(_gnd_net_),
            .in3(N__13256),
            .lcout(\uu2.un28_w_addr_user_i_0_a2_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_4 .LUT_INIT=16'b1101111111010101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_2_LC_5_6_4  (
            .in0(N__14481),
            .in1(N__17577),
            .in2(N__14366),
            .in3(N__17436),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_5 .LUT_INIT=16'b1101100010111010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_2_LC_5_6_5  (
            .in0(N__13080),
            .in1(N__14357),
            .in2(N__11358),
            .in3(N__14482),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_0_LC_5_6_6 .LUT_INIT=16'b0010001011101110;
    LogicCell40 \Lab_UT.dispString.dOut_0_LC_5_6_6  (
            .in0(N__12612),
            .in1(N__13084),
            .in2(_gnd_net_),
            .in3(N__12621),
            .lcout(L3_tx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21635),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_6_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_2_LC_5_6_7 .LUT_INIT=16'b1111101100111011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_2_LC_5_6_7  (
            .in0(N__12411),
            .in1(N__11600),
            .in2(N__13091),
            .in3(N__17294),
            .lcout(\Lab_UT.dispString.dOutP_0_iv_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_4_LC_5_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_4_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_4_LC_5_7_0 .LUT_INIT=16'b0101101011001111;
    LogicCell40 \Lab_UT.dispString.dOut_4_LC_5_7_0  (
            .in0(N__14476),
            .in1(N__11601),
            .in2(N__13092),
            .in3(N__13239),
            .lcout(L3_tx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21626),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_7_1 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \uu2.vram_rd_clk_det_RNI95711_1_LC_5_7_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uu2.vram_rd_clk_det_RNI95711_1_LC_5_7_1  (
            .in0(N__13839),
            .in1(N__13821),
            .in2(_gnd_net_),
            .in3(N__19278),
            .lcout(\uu2.vram_rd_clk_det_RNI95711Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_3_LC_5_7_2 .LUT_INIT=16'b0101110101010101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_3_LC_5_7_2  (
            .in0(N__14253),
            .in1(N__14965),
            .in2(N__14488),
            .in3(N__16638),
            .lcout(\Lab_UT.dispString.N_219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_0_a3_4_LC_5_7_5 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_0_a3_4_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_0_a3_4_LC_5_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uu2.un1_w_user_cr_0_a3_4_LC_5_7_5  (
            .in0(N__11155),
            .in1(N__11320),
            .in2(N__12725),
            .in3(N__13255),
            .lcout(),
            .ltout(\uu2.un1_w_user_cr_0_a3Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.un1_w_user_cr_0_a3_LC_5_7_6 .C_ON=1'b0;
    defparam \uu2.un1_w_user_cr_0_a3_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \uu2.un1_w_user_cr_0_a3_LC_5_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uu2.un1_w_user_cr_0_a3_LC_5_7_6  (
            .in0(N__12766),
            .in1(N__11302),
            .in2(N__11286),
            .in3(N__11275),
            .lcout(\uu2.un1_w_user_cr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_5_LC_5_7_7 .LUT_INIT=16'b0111011101111110;
    LogicCell40 \Lab_UT.dispString.dOut_5_LC_5_7_7  (
            .in0(N__14365),
            .in1(N__13089),
            .in2(N__14489),
            .in3(N__12675),
            .lcout(L3_tx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21626),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_1_LC_5_8_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_1_LC_5_8_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_1_LC_5_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_1_LC_5_8_0  (
            .in0(N__13183),
            .in1(N__11412),
            .in2(_gnd_net_),
            .in3(N__11451),
            .lcout(\buart.Z_tx.shifterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_0_LC_5_8_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_0_LC_5_8_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_0_LC_5_8_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \buart.Z_tx.shifter_0_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__11445),
            .in2(_gnd_net_),
            .in3(N__13181),
            .lcout(\buart.Z_tx.shifterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.uart_tx_LC_5_8_2 .C_ON=1'b0;
    defparam \buart.Z_tx.uart_tx_LC_5_8_2 .SEQ_MODE=4'b1011;
    defparam \buart.Z_tx.uart_tx_LC_5_8_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \buart.Z_tx.uart_tx_LC_5_8_2  (
            .in0(N__13182),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11439),
            .lcout(o_serial_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_2_LC_5_8_3 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_2_LC_5_8_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_2_LC_5_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_2_LC_5_8_3  (
            .in0(N__11400),
            .in1(N__13184),
            .in2(_gnd_net_),
            .in3(N__11418),
            .lcout(\buart.Z_tx.shifterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_3_LC_5_8_4 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_3_LC_5_8_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_3_LC_5_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_3_LC_5_8_4  (
            .in0(N__13185),
            .in1(N__11388),
            .in2(_gnd_net_),
            .in3(N__11406),
            .lcout(\buart.Z_tx.shifterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_4_LC_5_8_5 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_4_LC_5_8_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_4_LC_5_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_4_LC_5_8_5  (
            .in0(N__11376),
            .in1(N__13186),
            .in2(_gnd_net_),
            .in3(N__11394),
            .lcout(\buart.Z_tx.shifterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_5_LC_5_8_6 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_5_LC_5_8_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_5_LC_5_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_5_LC_5_8_6  (
            .in0(N__13187),
            .in1(N__11364),
            .in2(_gnd_net_),
            .in3(N__11382),
            .lcout(\buart.Z_tx.shifterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.shifter_6_LC_5_8_7 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_6_LC_5_8_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_6_LC_5_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \buart.Z_tx.shifter_6_LC_5_8_7  (
            .in0(N__13224),
            .in1(N__13188),
            .in2(_gnd_net_),
            .in3(N__11370),
            .lcout(\buart.Z_tx.shifterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21619),
            .ce(N__13115),
            .sr(N__19221));
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_9_0 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_9_0 .LUT_INIT=16'b1111101100000000;
    LogicCell40 \buart.Z_tx.bitcount_RNIVE1P1_2_LC_5_9_0  (
            .in0(N__11475),
            .in1(N__11568),
            .in2(N__11498),
            .in3(N__13338),
            .lcout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2 ),
            .ltout(\buart.Z_tx.bitcount_RNIVE1P1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_5_9_1 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNI22V22_2_LC_5_9_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \buart.Z_tx.bitcount_RNI22V22_2_LC_5_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11604),
            .in3(N__13180),
            .lcout(\buart.Z_tx.un1_uart_wr_i_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_5_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.cnt_RNIFV4E_1_LC_5_9_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dispString.cnt_RNIFV4E_1_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(N__14297),
            .in2(_gnd_net_),
            .in3(N__14407),
            .lcout(\Lab_UT.dispString.N_191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_9_3 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_2_LC_5_9_3 .LUT_INIT=16'b1100100111001100;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_2_LC_5_9_3  (
            .in0(N__11517),
            .in1(N__11494),
            .in2(N__11481),
            .in3(N__11540),
            .lcout(\buart.Z_tx.bitcount_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_9_4 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_9_4 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \buart.Z_tx.bitcount_RNIDCDL_3_LC_5_9_4  (
            .in0(N__11579),
            .in1(N__11516),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\buart.Z_tx.uart_busy_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_9_5 .C_ON=1'b0;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.hh_RNIJ3K62_0_LC_5_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \buart.Z_rx.hh_RNIJ3K62_0_LC_5_9_5  (
            .in0(N__14653),
            .in1(N__11562),
            .in2(_gnd_net_),
            .in3(N__11745),
            .lcout(\buart.Z_rx.startbit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_9_6 .C_ON=1'b0;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.bitcount_RNO_0_3_LC_5_9_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \buart.Z_tx.bitcount_RNO_0_3_LC_5_9_6  (
            .in0(N__11541),
            .in1(N__11518),
            .in2(N__11499),
            .in3(N__11479),
            .lcout(\buart.Z_tx.un1_bitcount_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_10_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_sbtinv_4_LC_5_10_0 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \buart.Z_rx.bitcount_sbtinv_4_LC_5_10_0  (
            .in0(N__18987),
            .in1(N__11796),
            .in2(N__11904),
            .in3(N__11744),
            .lcout(\buart.Z_rx.bitcounte_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_10_1 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_1_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_1_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__13009),
            .in2(_gnd_net_),
            .in3(N__12986),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21607),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_10_2 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNI5M6E_1_LC_5_10_2  (
            .in0(N__12985),
            .in1(N__13364),
            .in2(N__13011),
            .in3(N__13272),
            .lcout(\buart.Z_tx.ser_clk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_5_10_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_5_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIOP0V3_0_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__11743),
            .in2(_gnd_net_),
            .in3(N__18986),
            .lcout(\buart.Z_rx.N_27_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.rst_LC_5_10_4 .C_ON=1'b0;
    defparam \resetGen.rst_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \resetGen.rst_LC_5_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \resetGen.rst_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21399),
            .lcout(rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21607),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_10_7 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_0_LC_5_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_0_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13008),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21607),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_5_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_5_11_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIIVPI1_4_LC_5_11_0  (
            .in0(N__11626),
            .in1(N__11651),
            .in2(N__11712),
            .in3(N__11679),
            .lcout(\buart.Z_rx.un1_sample_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIQ0DP_4_LC_5_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIQ0DP_4_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIQ0DP_4_LC_5_11_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIQ0DP_4_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(N__11650),
            .in2(_gnd_net_),
            .in3(N__11624),
            .lcout(),
            .ltout(\buart.Z_rx.idle_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_11_2 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_11_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_0_LC_5_11_2  (
            .in0(N__11680),
            .in1(N__11706),
            .in2(N__11748),
            .in3(N__11865),
            .lcout(\buart.Z_rx.idle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_3_LC_5_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_3_LC_5_11_3 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_3_LC_5_11_3 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_es_3_LC_5_11_3  (
            .in0(N__11707),
            .in1(N__12059),
            .in2(N__11724),
            .in3(N__11829),
            .lcout(\buart.Z_rx.bitcountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21601),
            .ce(N__12026),
            .sr(N__19233));
    defparam \buart.Z_rx.bitcount_es_RNINTCP_0_LC_5_11_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNINTCP_0_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNINTCP_0_LC_5_11_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.bitcount_es_RNINTCP_0_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(N__11705),
            .in2(_gnd_net_),
            .in3(N__11864),
            .lcout(),
            .ltout(\buart.Z_rx.valid_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_11_5 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_11_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNISCGV1_4_LC_5_11_5  (
            .in0(N__11678),
            .in1(N__11649),
            .in2(N__11631),
            .in3(N__11625),
            .lcout(bu_rx_data_rdy),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_0_LC_5_11_7 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_0_LC_5_11_7 .SEQ_MODE=4'b1011;
    defparam \buart.Z_rx.bitcount_es_0_LC_5_11_7 .LUT_INIT=16'b0001001011011110;
    LogicCell40 \buart.Z_rx.bitcount_es_0_LC_5_11_7  (
            .in0(N__11866),
            .in1(N__12058),
            .in2(N__15759),
            .in3(N__11828),
            .lcout(\buart.Z_rx.bitcountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21601),
            .ce(N__12026),
            .sr(N__19233));
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_1_LC_5_12_0 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_1_LC_5_12_0  (
            .in0(N__11824),
            .in1(_gnd_net_),
            .in2(N__11771),
            .in3(N__11939),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21595),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_4_LC_5_12_1 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_4_LC_5_12_1  (
            .in0(N__11900),
            .in1(N__11825),
            .in2(N__11991),
            .in3(N__11997),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21595),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_12_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI5JE3_5_LC_5_12_2  (
            .in0(N__11986),
            .in1(N__11969),
            .in2(N__11957),
            .in3(N__11938),
            .lcout(),
            .ltout(\buart.Z_rx.Z_baudgen.ser_clk_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_12_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_RNI3O55_2_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__11920),
            .in2(N__11907),
            .in3(N__11763),
            .lcout(\buart.Z_rx.ser_clk ),
            .ltout(\buart.Z_rx.ser_clk_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_12_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \buart.Z_rx.bitcount_es_RNIV4M42_0_LC_5_12_4  (
            .in0(N__11877),
            .in1(_gnd_net_),
            .in2(N__11871),
            .in3(N__11868),
            .lcout(\buart.Z_rx.sample ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \buart.Z_rx.Z_baudgen.counter_0_LC_5_12_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \buart.Z_rx.Z_baudgen.counter_0_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__11764),
            .in2(_gnd_net_),
            .in3(N__11826),
            .lcout(\buart.Z_rx.Z_baudgen.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21595),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g1_5_LC_5_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_5_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_5_LC_5_13_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.g1_5_LC_5_13_4  (
            .in0(N__18875),
            .in1(N__20161),
            .in2(N__21355),
            .in3(N__19933),
            .lcout(\Lab_UT.dictrl.g1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJAJ21_LC_5_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJAJ21_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIJAJ21_LC_5_13_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIJAJ21_LC_5_13_5  (
            .in0(N__18494),
            .in1(N__21348),
            .in2(N__20937),
            .in3(N__18876),
            .lcout(\Lab_UT.dictrl.g0_17_a6_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_168_LC_6_1_0 .C_ON=1'b0;
    defparam \uu2.bitmap_168_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_168_LC_6_1_0 .LUT_INIT=16'b0001011001010110;
    LogicCell40 \uu2.bitmap_168_LC_6_1_0  (
            .in0(N__13437),
            .in1(N__13603),
            .in2(N__13547),
            .in3(N__13576),
            .lcout(\uu2.bitmapZ0Z_168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__19180));
    defparam \uu2.bitmap_RNISSSN_162_LC_6_1_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNISSSN_162_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNISSSN_162_LC_6_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNISSSN_162_LC_6_1_1  (
            .in0(N__12108),
            .in1(N__12090),
            .in2(_gnd_net_),
            .in3(N__12129),
            .lcout(\uu2.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_75_LC_6_1_2 .C_ON=1'b0;
    defparam \uu2.bitmap_75_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_75_LC_6_1_2 .LUT_INIT=16'b0110011100011111;
    LogicCell40 \uu2.bitmap_75_LC_6_1_2  (
            .in0(N__13439),
            .in1(N__13607),
            .in2(N__13548),
            .in3(N__13578),
            .lcout(\uu2.bitmapZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__19180));
    defparam \uu2.bitmap_203_LC_6_1_3 .C_ON=1'b0;
    defparam \uu2.bitmap_203_LC_6_1_3 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_203_LC_6_1_3 .LUT_INIT=16'b0011101111101111;
    LogicCell40 \uu2.bitmap_203_LC_6_1_3  (
            .in0(N__13577),
            .in1(N__13530),
            .in2(N__13608),
            .in3(N__13438),
            .lcout(\uu2.bitmapZ0Z_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__19180));
    defparam \uu2.bitmap_RNIM9P11_75_LC_6_1_4 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIM9P11_75_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIM9P11_75_LC_6_1_4 .LUT_INIT=16'b0010011101010101;
    LogicCell40 \uu2.bitmap_RNIM9P11_75_LC_6_1_4  (
            .in0(N__12578),
            .in1(N__12123),
            .in2(N__12117),
            .in3(N__12475),
            .lcout(\uu2.bitmap_pmux_24_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_162_LC_6_1_5 .C_ON=1'b0;
    defparam \uu2.bitmap_162_LC_6_1_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_162_LC_6_1_5 .LUT_INIT=16'b0001011000110110;
    LogicCell40 \uu2.bitmap_162_LC_6_1_5  (
            .in0(N__12435),
            .in1(N__13404),
            .in2(N__13658),
            .in3(N__13621),
            .lcout(\uu2.bitmapZ0Z_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__19180));
    defparam \uu2.bitmap_290_LC_6_1_6 .C_ON=1'b0;
    defparam \uu2.bitmap_290_LC_6_1_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_290_LC_6_1_6 .LUT_INIT=16'b0000011100011001;
    LogicCell40 \uu2.bitmap_290_LC_6_1_6  (
            .in0(N__13622),
            .in1(N__13654),
            .in2(N__13419),
            .in3(N__12436),
            .lcout(\uu2.bitmapZ0Z_290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_168C_net ),
            .ce(),
            .sr(N__19180));
    defparam \uu2.bitmap_RNI4LQU_34_LC_6_1_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI4LQU_34_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI4LQU_34_LC_6_1_7 .LUT_INIT=16'b0000110100111101;
    LogicCell40 \uu2.bitmap_RNI4LQU_34_LC_6_1_7  (
            .in0(N__12102),
            .in1(N__12089),
            .in2(N__12201),
            .in3(N__12066),
            .lcout(\uu2.bitmap_pmux_15_i_m2_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_296_LC_6_2_0 .C_ON=1'b0;
    defparam \uu2.bitmap_296_LC_6_2_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_296_LC_6_2_0 .LUT_INIT=16'b0001001000100111;
    LogicCell40 \uu2.bitmap_296_LC_6_2_0  (
            .in0(N__13600),
            .in1(N__13452),
            .in2(N__13549),
            .in3(N__13573),
            .lcout(\uu2.bitmapZ0Z_296 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__19178));
    defparam \uu2.bitmap_200_LC_6_2_1 .C_ON=1'b0;
    defparam \uu2.bitmap_200_LC_6_2_1 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_200_LC_6_2_1 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \uu2.bitmap_200_LC_6_2_1  (
            .in0(N__13572),
            .in1(N__13537),
            .in2(N__13455),
            .in3(N__13599),
            .lcout(\uu2.bitmapZ0Z_200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__19178));
    defparam \uu2.bitmap_72_LC_6_2_2 .C_ON=1'b0;
    defparam \uu2.bitmap_72_LC_6_2_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_72_LC_6_2_2 .LUT_INIT=16'b0001010000110101;
    LogicCell40 \uu2.bitmap_72_LC_6_2_2  (
            .in0(N__13602),
            .in1(N__13454),
            .in2(N__13551),
            .in3(N__13575),
            .lcout(\uu2.bitmapZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__19178));
    defparam \uu2.bitmap_RNI5T9T1_72_LC_6_2_3 .C_ON=1'b0;
    defparam \uu2.bitmap_RNI5T9T1_72_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNI5T9T1_72_LC_6_2_3 .LUT_INIT=16'b0101010111100100;
    LogicCell40 \uu2.bitmap_RNI5T9T1_72_LC_6_2_3  (
            .in0(N__12402),
            .in1(N__12396),
            .in2(N__12390),
            .in3(N__12373),
            .lcout(\uu2.bitmap_RNI5T9T1Z0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_40_LC_6_2_4 .C_ON=1'b0;
    defparam \uu2.bitmap_40_LC_6_2_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_40_LC_6_2_4 .LUT_INIT=16'b1011011011101111;
    LogicCell40 \uu2.bitmap_40_LC_6_2_4  (
            .in0(N__13601),
            .in1(N__13453),
            .in2(N__13550),
            .in3(N__13574),
            .lcout(\uu2.bitmapZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_296C_net ),
            .ce(),
            .sr(N__19178));
    defparam \uu2.bitmap_RNIGQ8J1_111_LC_6_2_5 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIGQ8J1_111_LC_6_2_5 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIGQ8J1_111_LC_6_2_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uu2.bitmap_RNIGQ8J1_111_LC_6_2_5  (
            .in0(N__12306),
            .in1(N__13881),
            .in2(_gnd_net_),
            .in3(N__12297),
            .lcout(),
            .ltout(\uu2.N_395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_displaying_fast_RNIL9SE4_2_LC_6_2_6 .C_ON=1'b0;
    defparam \uu2.w_addr_displaying_fast_RNIL9SE4_2_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_displaying_fast_RNIL9SE4_2_LC_6_2_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uu2.w_addr_displaying_fast_RNIL9SE4_2_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__12291),
            .in2(N__12282),
            .in3(N__12207),
            .lcout(\uu2.N_401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_RNIURJN1_40_LC_6_2_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIURJN1_40_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIURJN1_40_LC_6_2_7 .LUT_INIT=16'b1100000010111011;
    LogicCell40 \uu2.bitmap_RNIURJN1_40_LC_6_2_7  (
            .in0(N__12270),
            .in1(N__12258),
            .in2(N__12225),
            .in3(N__12213),
            .lcout(\uu2.N_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_308_LC_6_3_0 .C_ON=1'b0;
    defparam \uu2.bitmap_308_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_308_LC_6_3_0 .LUT_INIT=16'b0000011000011101;
    LogicCell40 \uu2.bitmap_308_LC_6_3_0  (
            .in0(N__13773),
            .in1(N__13746),
            .in2(N__14232),
            .in3(N__13716),
            .lcout(\uu2.bitmapZ0Z_308 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__19176));
    defparam \uu2.bitmap_RNIU2IS_52_LC_6_3_1 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIU2IS_52_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIU2IS_52_LC_6_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uu2.bitmap_RNIU2IS_52_LC_6_3_1  (
            .in0(N__12588),
            .in1(N__12190),
            .in2(_gnd_net_),
            .in3(N__12141),
            .lcout(\uu2.bitmap_RNIU2ISZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.bitmap_52_LC_6_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_52_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_52_LC_6_3_2 .LUT_INIT=16'b1001111011111101;
    LogicCell40 \uu2.bitmap_52_LC_6_3_2  (
            .in0(N__13774),
            .in1(N__13747),
            .in2(N__14233),
            .in3(N__13717),
            .lcout(\uu2.bitmapZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__19176));
    defparam \uu2.bitmap_84_LC_6_3_4 .C_ON=1'b0;
    defparam \uu2.bitmap_84_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_84_LC_6_3_4 .LUT_INIT=16'b0001001000011011;
    LogicCell40 \uu2.bitmap_84_LC_6_3_4  (
            .in0(N__13775),
            .in1(N__13748),
            .in2(N__14234),
            .in3(N__13718),
            .lcout(\uu2.bitmapZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__19176));
    defparam \uu2.bitmap_87_LC_6_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_87_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_87_LC_6_3_6 .LUT_INIT=16'b0011110101010111;
    LogicCell40 \uu2.bitmap_87_LC_6_3_6  (
            .in0(N__13776),
            .in1(N__13749),
            .in2(N__14235),
            .in3(N__13719),
            .lcout(\uu2.bitmapZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.bitmap_308C_net ),
            .ce(),
            .sr(N__19176));
    defparam \uu2.bitmap_RNIG5UR_84_LC_6_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_RNIG5UR_84_LC_6_3_7 .SEQ_MODE=4'b0000;
    defparam \uu2.bitmap_RNIG5UR_84_LC_6_3_7 .LUT_INIT=16'b0000101001110111;
    LogicCell40 \uu2.bitmap_RNIG5UR_84_LC_6_3_7  (
            .in0(N__12580),
            .in1(N__12504),
            .in2(N__12498),
            .in3(N__12487),
            .lcout(\uu2.bitmap_pmux_24_am_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI8CKM3_1_LC_6_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI8CKM3_1_LC_6_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI8CKM3_1_LC_6_4_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI8CKM3_1_LC_6_4_0  (
            .in0(N__16823),
            .in1(N__14564),
            .in2(_gnd_net_),
            .in3(N__15386),
            .lcout(\Lab_UT.sec1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNIAEKM3_2_LC_6_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNIAEKM3_2_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNIAEKM3_2_LC_6_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNIAEKM3_2_LC_6_4_1  (
            .in0(N__14563),
            .in1(N__15633),
            .in2(_gnd_net_),
            .in3(N__17573),
            .lcout(\Lab_UT.sec1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNILUSP3_1_LC_6_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNILUSP3_1_LC_6_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNILUSP3_1_LC_6_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNILUSP3_1_LC_6_4_4  (
            .in0(N__14580),
            .in1(N__14125),
            .in2(_gnd_net_),
            .in3(N__14180),
            .lcout(\Lab_UT.min1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_6_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_1_LC_6_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_1_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20303),
            .lcout(\Lab_UT.di_AMtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21638),
            .ce(N__16604),
            .sr(N__19209));
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_6_4_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_6_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_3_2_LC_6_4_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_3_2_LC_6_4_6  (
            .in0(N__12702),
            .in1(N__13928),
            .in2(_gnd_net_),
            .in3(N__14159),
            .lcout(\Lab_UT.dispString.un46_dOutP_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_6_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_2_LC_6_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_2_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20766),
            .lcout(\Lab_UT.di_AMtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21638),
            .ce(N__16604),
            .sr(N__19209));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH9JB1_0_LC_6_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH9JB1_0_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIH9JB1_0_LC_6_5_0 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIH9JB1_0_LC_6_5_0  (
            .in0(N__15426),
            .in1(N__16843),
            .in2(N__12606),
            .in3(N__18034),
            .lcout(\Lab_UT.didp.did_alarmMatch_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIDIHR3_0_LC_6_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIDIHR3_0_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIDIHR3_0_LC_6_5_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIDIHR3_0_LC_6_5_1  (
            .in0(N__12604),
            .in1(N__14561),
            .in2(_gnd_net_),
            .in3(N__18035),
            .lcout(\Lab_UT.sec2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNI6AKM3_0_LC_6_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNI6AKM3_0_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNI6AKM3_0_LC_6_5_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNI6AKM3_0_LC_6_5_2  (
            .in0(N__14562),
            .in1(_gnd_net_),
            .in2(N__15435),
            .in3(N__16844),
            .lcout(\Lab_UT.sec1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_0_LC_6_5_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_0_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_0_LC_6_5_3 .LUT_INIT=16'b1100100011111111;
    LogicCell40 \Lab_UT.alarmchar_latch_0_LC_6_5_3  (
            .in0(N__12635),
            .in1(N__17768),
            .in2(N__19290),
            .in3(N__17834),
            .lcout(G_190),
            .ltout(G_190_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_0_LC_6_5_4 .LUT_INIT=16'b0110010001110101;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_0_LC_6_5_4  (
            .in0(N__14335),
            .in1(N__14456),
            .in2(N__12624),
            .in3(N__12605),
            .lcout(\Lab_UT.dispString.i21_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_0_LC_6_5_5 .LUT_INIT=16'b0001110100110011;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_0_LC_6_5_5  (
            .in0(N__17505),
            .in1(N__14334),
            .in2(N__16848),
            .in3(N__14471),
            .lcout(),
            .ltout(\Lab_UT.dispString.m28_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_0_LC_6_5_6 .LUT_INIT=16'b0100101000001010;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_0_LC_6_5_6  (
            .in0(N__14472),
            .in1(N__15011),
            .in2(N__12615),
            .in3(N__17172),
            .lcout(\Lab_UT.dispString.N_204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_0_LC_6_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_0_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19955),
            .lcout(\Lab_UT.di_ASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21629),
            .ce(N__18663),
            .sr(N__19206));
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_6_0 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_6_0 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \uu2.w_addr_user_nesr_RNIF1S9_5_LC_6_6_0  (
            .in0(N__12972),
            .in1(N__12842),
            .in2(N__12881),
            .in3(N__12925),
            .lcout(\uu2.N_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_nesr_5_LC_6_6_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_nesr_5_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_nesr_5_LC_6_6_1 .LUT_INIT=16'b0000000011010010;
    LogicCell40 \uu2.w_addr_user_nesr_5_LC_6_6_1  (
            .in0(N__12926),
            .in1(N__12877),
            .in2(N__12851),
            .in3(N__14077),
            .lcout(\uu2.w_addr_userZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_nesr_5C_net ),
            .ce(N__12816),
            .sr(N__19170));
    defparam \Lab_UT.dictrl.m59_ns_1_ns_LC_6_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m59_ns_1_ns_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m59_ns_1_ns_LC_6_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.dictrl.m59_ns_1_ns_LC_6_6_5  (
            .in0(N__16223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16203),
            .lcout(\Lab_UT.dictrl.m59_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_3_LC_6_7_0 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_3_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_3_LC_6_7_0 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.alarmchar_latch_3_LC_6_7_0  (
            .in0(N__15752),
            .in1(N__15774),
            .in2(N__12804),
            .in3(N__14625),
            .lcout(G_193),
            .ltout(G_193_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_3_LC_6_7_1 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_3_LC_6_7_1  (
            .in0(N__14340),
            .in1(N__14441),
            .in2(N__12795),
            .in3(N__17264),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_3_LC_6_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_3_LC_6_7_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_3_LC_6_7_2 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \Lab_UT.dispString.dOut_3_LC_6_7_2  (
            .in0(N__12792),
            .in1(_gnd_net_),
            .in2(N__12786),
            .in3(N__13069),
            .lcout(L3_tx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21615),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_6_LC_6_7_3 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_6_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_6_LC_6_7_3 .LUT_INIT=16'b0011000100100010;
    LogicCell40 \Lab_UT.alarmchar_latch_6_LC_6_7_3  (
            .in0(N__17769),
            .in1(N__15500),
            .in2(N__12753),
            .in3(N__17835),
            .lcout(G_189),
            .ltout(G_189_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_6_LC_6_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_6_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_6_LC_6_7_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \Lab_UT.dispString.dOut_6_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12744),
            .in3(N__12741),
            .lcout(L3_tx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21615),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_6_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_5_LC_6_7_5 .LUT_INIT=16'b0000010011110100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_5_LC_6_7_5  (
            .in0(N__12701),
            .in1(N__13918),
            .in2(N__14361),
            .in3(N__14615),
            .lcout(\Lab_UT.dispString.m44_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_1_LC_6_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_1_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.dOut_1_LC_6_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.dispString.dOut_1_LC_6_7_6  (
            .in0(N__13506),
            .in1(N__13068),
            .in2(_gnd_net_),
            .in3(N__14496),
            .lcout(L3_tx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21615),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_6_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_4_LC_6_7_7 .LUT_INIT=16'b0000000111110001;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_4_LC_6_7_7  (
            .in0(N__14336),
            .in1(N__15005),
            .in2(N__13085),
            .in3(N__14614),
            .lcout(\Lab_UT.dispString.m42_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.shifter_7_LC_6_8_0 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_7_LC_6_8_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_7_LC_6_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \buart.Z_tx.shifter_7_LC_6_8_0  (
            .in0(N__13201),
            .in1(N__13125),
            .in2(_gnd_net_),
            .in3(N__13233),
            .lcout(\buart.Z_tx.shifterZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21610),
            .ce(N__13119),
            .sr(N__19225));
    defparam \buart.Z_tx.shifter_8_LC_6_8_1 .C_ON=1'b0;
    defparam \buart.Z_tx.shifter_8_LC_6_8_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_tx.shifter_8_LC_6_8_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \buart.Z_tx.shifter_8_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__13200),
            .in2(_gnd_net_),
            .in3(N__13134),
            .lcout(\buart.Z_tx.shifterZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21610),
            .ce(N__13119),
            .sr(N__19225));
    defparam \Lab_UT.dispString.cnt_1_LC_6_9_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_1_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_1_LC_6_9_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.dispString.cnt_1_LC_6_9_0  (
            .in0(N__14311),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14455),
            .lcout(\Lab_UT.dispString.cntZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21603),
            .ce(),
            .sr(N__19204));
    defparam \Lab_UT.dispString.cnt_0_LC_6_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_0_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_0_LC_6_9_2 .LUT_INIT=16'b0011001100110010;
    LogicCell40 \Lab_UT.dispString.cnt_0_LC_6_9_2  (
            .in0(N__14310),
            .in1(N__14454),
            .in2(N__13078),
            .in3(N__15012),
            .lcout(\Lab_UT.dispString.cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21603),
            .ce(),
            .sr(N__19204));
    defparam \Lab_UT.dispString.cnt_2_LC_6_9_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.cnt_2_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dispString.cnt_2_LC_6_9_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \Lab_UT.dispString.cnt_2_LC_6_9_7  (
            .in0(N__14453),
            .in1(N__14312),
            .in2(_gnd_net_),
            .in3(N__13055),
            .lcout(\Lab_UT.dispString.cntZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21603),
            .ce(),
            .sr(N__19204));
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_10_0 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \buart.Z_tx.Z_baudgen.un2_counter_cry_1_c_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(N__13010),
            .in2(N__12990),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_10_1 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_2_LC_6_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_2_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(N__13365),
            .in2(_gnd_net_),
            .in3(N__13353),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_2 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_1 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .clk(N__21598),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_10_2 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_3_LC_6_10_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_3_LC_6_10_2  (
            .in0(N__13340),
            .in1(N__13281),
            .in2(_gnd_net_),
            .in3(N__13350),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_3 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_2 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .clk(N__21598),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_10_3 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_4_LC_6_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_4_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13308),
            .in3(N__13347),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_4 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_3 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .clk(N__21598),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_10_4 .C_ON=1'b1;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_5_LC_6_10_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_5_LC_6_10_4  (
            .in0(N__13341),
            .in1(_gnd_net_),
            .in2(N__13320),
            .in3(N__13344),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_5 ),
            .ltout(),
            .carryin(\buart.Z_tx.Z_baudgen.un2_counter_cry_4 ),
            .carryout(\buart.Z_tx.Z_baudgen.un2_counter_cry_5 ),
            .clk(N__21598),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_10_5 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \buart.Z_tx.Z_baudgen.counter_6_LC_6_10_5 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_6_LC_6_10_5  (
            .in0(N__13295),
            .in1(N__13339),
            .in2(_gnd_net_),
            .in3(N__13323),
            .lcout(\buart.Z_tx.Z_baudgen.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21598),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_6_10_6 .C_ON=1'b0;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_6_10_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \buart.Z_tx.Z_baudgen.counter_RNII048_6_LC_6_10_6  (
            .in0(N__13316),
            .in1(N__13304),
            .in2(N__13296),
            .in3(N__13280),
            .lcout(\buart.Z_tx.Z_baudgen.ser_clk_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUJLP6_1_LC_6_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUJLP6_1_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUJLP6_1_LC_6_10_7 .LUT_INIT=16'b0000010011001000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUJLP6_1_LC_6_10_7  (
            .in0(N__16290),
            .in1(N__14844),
            .in2(N__21261),
            .in3(N__19641),
            .lcout(\Lab_UT.dictrl.N_95_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_LC_6_11_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_LC_6_11_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_LC_6_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14660),
            .lcout(bu_rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21594),
            .ce(N__19316),
            .sr(N__19235));
    defparam \buart.Z_rx.shifter_fast_7_LC_6_11_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_7_LC_6_11_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_7_LC_6_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_7_LC_6_11_1  (
            .in0(N__14661),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21594),
            .ce(N__19316),
            .sr(N__19235));
    defparam \buart.Z_rx.shifter_fast_6_LC_6_11_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_6_LC_6_11_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_6_LC_6_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_6_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20362),
            .lcout(buart__rx_shifter_fast_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21594),
            .ce(N__19316),
            .sr(N__19235));
    defparam \buart.Z_rx.shifter_6_LC_6_11_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_6_LC_6_11_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_6_LC_6_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_6_LC_6_11_6  (
            .in0(N__20363),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21594),
            .ce(N__19316),
            .sr(N__19235));
    defparam \Lab_UT.dictrl.state_0_esr_RNIU7683_2_LC_6_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIU7683_2_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIU7683_2_LC_6_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIU7683_2_LC_6_12_0  (
            .in0(N__16449),
            .in1(N__20029),
            .in2(N__19810),
            .in3(N__13377),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI88DT7_1_LC_6_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI88DT7_1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI88DT7_1_LC_6_12_1 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI88DT7_1_LC_6_12_1  (
            .in0(N__19665),
            .in1(N__21250),
            .in2(N__13371),
            .in3(N__14877),
            .lcout(\Lab_UT.dictrl.N_90_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m30_0_0_LC_6_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m30_0_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m30_0_0_LC_6_12_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \Lab_UT.dictrl.m30_0_0_LC_6_12_2  (
            .in0(N__14896),
            .in1(_gnd_net_),
            .in2(N__18429),
            .in3(N__18941),
            .lcout(\Lab_UT.dictrl.m30_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_17_LC_6_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_17_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_17_LC_6_12_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_17_LC_6_12_4  (
            .in0(N__18424),
            .in1(N__16131),
            .in2(N__16519),
            .in3(N__18942),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_14_LC_6_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_14_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_14_LC_6_12_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_14_LC_6_12_5  (
            .in0(N__16732),
            .in1(N__16448),
            .in2(N__13368),
            .in3(N__19497),
            .lcout(\Lab_UT.dictrl.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIHC6L_1_LC_6_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIHC6L_1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIHC6L_1_LC_6_12_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIHC6L_1_LC_6_12_7  (
            .in0(N__14734),
            .in1(N__16367),
            .in2(N__21044),
            .in3(N__20929),
            .lcout(\Lab_UT.dictrl.g0_17_a6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNINEHL_LC_6_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNINEHL_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNINEHL_LC_6_13_0 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNINEHL_LC_6_13_0  (
            .in0(N__18868),
            .in1(N__16259),
            .in2(N__21104),
            .in3(N__18381),
            .lcout(\Lab_UT.dictrl.g0_17_a6_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_17_a6_1_6_LC_6_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_a6_1_6_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_a6_1_6_LC_6_13_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.g0_17_a6_1_6_LC_6_13_1  (
            .in0(N__19496),
            .in1(N__20374),
            .in2(N__21356),
            .in3(N__20595),
            .lcout(\Lab_UT.dictrl.g0_17_a6_1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI7FC61_LC_6_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI7FC61_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI7FC61_LC_6_13_2 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNI7FC61_LC_6_13_2  (
            .in0(N__16380),
            .in1(N__18753),
            .in2(N__20163),
            .in3(N__20934),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_17_a6_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIU4P66_LC_6_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIU4P66_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIU4P66_LC_6_13_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIU4P66_LC_6_13_3  (
            .in0(N__13491),
            .in1(N__13485),
            .in2(N__13479),
            .in3(N__13467),
            .lcout(\Lab_UT.dictrl.g0_17_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_17_o6_1_4_LC_6_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_o6_1_4_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_o6_1_4_LC_6_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \Lab_UT.dictrl.g0_17_o6_1_4_LC_6_13_4  (
            .in0(N__19495),
            .in1(N__20142),
            .in2(N__18633),
            .in3(N__18380),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_17_o6_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIG3243_1_LC_6_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIG3243_1_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIG3243_1_LC_6_13_5 .LUT_INIT=16'b1111110000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIG3243_1_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__13461),
            .in2(N__13476),
            .in3(N__13473),
            .lcout(\Lab_UT.dictrl.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIO3GC_LC_6_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIO3GC_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNIO3GC_LC_6_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNIO3GC_LC_6_13_6  (
            .in0(_gnd_net_),
            .in1(N__16710),
            .in2(_gnd_net_),
            .in3(N__16258),
            .lcout(\Lab_UT.dictrl.g0_17_a6_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_17_o6_1_5_LC_6_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_o6_1_5_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_o6_1_5_LC_6_13_7 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \Lab_UT.dictrl.g0_17_o6_1_5_LC_6_13_7  (
            .in0(N__18428),
            .in1(N__18867),
            .in2(N__16731),
            .in3(N__20594),
            .lcout(\Lab_UT.dictrl.g0_17_o6_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_1_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_1_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_3_LC_7_1_3  (
            .in0(N__15062),
            .in1(N__17208),
            .in2(_gnd_net_),
            .in3(N__14135),
            .lcout(\Lab_UT.didp.countrce4.un20_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNIEQ8R3_3_LC_7_1_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNIEQ8R3_3_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNIEQ8R3_3_LC_7_1_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNIEQ8R3_3_LC_7_1_4  (
            .in0(N__14568),
            .in1(N__17088),
            .in2(_gnd_net_),
            .in3(N__17358),
            .lcout(\Lab_UT.min2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIP2TP3_3_LC_7_1_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIP2TP3_3_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIP2TP3_3_LC_7_1_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIP2TP3_3_LC_7_1_5  (
            .in0(N__15476),
            .in1(N__14569),
            .in2(_gnd_net_),
            .in3(N__16634),
            .lcout(\Lab_UT.min1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIN0TP3_2_LC_7_1_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIN0TP3_2_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIN0TP3_2_LC_7_1_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIN0TP3_2_LC_7_1_6  (
            .in0(N__14566),
            .in1(N__15061),
            .in2(_gnd_net_),
            .in3(N__14163),
            .lcout(\Lab_UT.min1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIJSSP3_0_LC_7_1_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIJSSP3_0_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIJSSP3_0_LC_7_1_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIJSSP3_0_LC_7_1_7  (
            .in0(N__17171),
            .in1(N__17207),
            .in2(_gnd_net_),
            .in3(N__14567),
            .lcout(\Lab_UT.min1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_2_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_2_0 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_0_LC_7_2_0  (
            .in0(N__17203),
            .in1(N__15184),
            .in2(_gnd_net_),
            .in3(N__19948),
            .lcout(\Lab_UT.didp.countrce4.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_7_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_1_LC_7_2_1 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_1_LC_7_2_1  (
            .in0(N__17051),
            .in1(N__20304),
            .in2(N__16953),
            .in3(N__17004),
            .lcout(\Lab_UT.didp.countrce3.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.reset_RNO_0_3_LC_7_2_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \Lab_UT.didp.reset_RNO_0_3_LC_7_2_2  (
            .in0(N__17204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14136),
            .lcout(\Lab_UT.didp.reset_12_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNIAM8R3_1_LC_7_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNIAM8R3_1_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNIAM8R3_1_LC_7_2_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNIAM8R3_1_LC_7_2_3  (
            .in0(N__14583),
            .in1(N__17003),
            .in2(_gnd_net_),
            .in3(N__17465),
            .lcout(\Lab_UT.min2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNI8K8R3_0_LC_7_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNI8K8R3_0_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNI8K8R3_0_LC_7_2_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNI8K8R3_0_LC_7_2_4  (
            .in0(N__17050),
            .in1(N__14582),
            .in2(_gnd_net_),
            .in3(N__17504),
            .lcout(\Lab_UT.min2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNICO8R3_2_LC_7_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNICO8R3_2_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNICO8R3_2_LC_7_2_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNICO8R3_2_LC_7_2_5  (
            .in0(N__14581),
            .in1(N__16904),
            .in2(_gnd_net_),
            .in3(N__17435),
            .lcout(\Lab_UT.min2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_2_6 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_1_LC_7_2_6 .LUT_INIT=16'b0101001101011111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_1_LC_7_2_6  (
            .in0(N__17466),
            .in1(N__15013),
            .in2(N__14490),
            .in3(N__14184),
            .lcout(),
            .ltout(\Lab_UT.dispString.N_18_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_7_2_7 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_0_1_LC_7_2_7 .LUT_INIT=16'b1010111100100111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_0_1_LC_7_2_7  (
            .in0(N__14367),
            .in1(N__14487),
            .in2(N__13509),
            .in3(N__16824),
            .lcout(\Lab_UT.dispString.dOut_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uu2.w_addr_user_7_LC_7_3_1 .C_ON=1'b0;
    defparam \uu2.w_addr_user_7_LC_7_3_1 .SEQ_MODE=4'b1000;
    defparam \uu2.w_addr_user_7_LC_7_3_1 .LUT_INIT=16'b0010000110101010;
    LogicCell40 \uu2.w_addr_user_7_LC_7_3_1  (
            .in0(N__13953),
            .in1(N__14085),
            .in2(N__14031),
            .in3(N__13998),
            .lcout(\uu2.w_addr_userZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.bitmap_111_LC_7_3_2 .C_ON=1'b0;
    defparam \uu2.bitmap_111_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_111_LC_7_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.bitmap_111_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13929),
            .lcout(\uu2.bitmapZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.vram_rd_clk_det_0_LC_7_3_3 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_0_LC_7_3_3 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_0_LC_7_3_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uu2.vram_rd_clk_det_0_LC_7_3_3  (
            .in0(N__13871),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uu2.vram_rd_clk_detZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.vram_rd_clk_det_1_LC_7_3_4 .C_ON=1'b0;
    defparam \uu2.vram_rd_clk_det_1_LC_7_3_4 .SEQ_MODE=4'b1011;
    defparam \uu2.vram_rd_clk_det_1_LC_7_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uu2.vram_rd_clk_det_1_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13835),
            .lcout(\uu2.vram_rd_clk_detZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.bitmap_180_LC_7_3_5 .C_ON=1'b0;
    defparam \uu2.bitmap_180_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_180_LC_7_3_5 .LUT_INIT=16'b0001011000011110;
    LogicCell40 \uu2.bitmap_180_LC_7_3_5  (
            .in0(N__13777),
            .in1(N__13750),
            .in2(N__14229),
            .in3(N__13720),
            .lcout(\uu2.bitmapZ0Z_180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.bitmap_215_LC_7_3_6 .C_ON=1'b0;
    defparam \uu2.bitmap_215_LC_7_3_6 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_215_LC_7_3_6 .LUT_INIT=16'b0011111010111111;
    LogicCell40 \uu2.bitmap_215_LC_7_3_6  (
            .in0(N__13722),
            .in1(N__13779),
            .in2(N__14231),
            .in3(N__13752),
            .lcout(\uu2.bitmapZ0Z_215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \uu2.bitmap_212_LC_7_3_7 .C_ON=1'b0;
    defparam \uu2.bitmap_212_LC_7_3_7 .SEQ_MODE=4'b1000;
    defparam \uu2.bitmap_212_LC_7_3_7 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \uu2.bitmap_212_LC_7_3_7  (
            .in0(N__13778),
            .in1(N__13751),
            .in2(N__14230),
            .in3(N__13721),
            .lcout(\uu2.bitmapZ0Z_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuu2.w_addr_user_7C_net ),
            .ce(),
            .sr(N__19179));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_7_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_7_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_0_LC_7_4_0 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_0_LC_7_4_0  (
            .in0(N__16941),
            .in1(N__17052),
            .in2(_gnd_net_),
            .in3(N__19929),
            .lcout(\Lab_UT.didp.countrce3.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNICGKM3_3_LC_7_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNICGKM3_3_LC_7_4_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNICGKM3_3_LC_7_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNICGKM3_3_LC_7_4_1  (
            .in0(N__14565),
            .in1(N__15339),
            .in2(_gnd_net_),
            .in3(N__17543),
            .lcout(\Lab_UT.sec1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIAC7D1_1_LC_7_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIAC7D1_1_LC_7_4_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIAC7D1_1_LC_7_4_2 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIAC7D1_1_LC_7_4_2  (
            .in0(N__14179),
            .in1(N__15050),
            .in2(N__14134),
            .in3(N__14155),
            .lcout(\Lab_UT.didp.did_alarmMatch_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_4_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_4_3 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_1_LC_7_4_3  (
            .in0(N__14132),
            .in1(N__20302),
            .in2(N__15196),
            .in3(N__17206),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_1_LC_7_4_4 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \Lab_UT.didp.countrce4.q_1_LC_7_4_4  (
            .in0(N__15097),
            .in1(N__15138),
            .in2(N__14139),
            .in3(N__14133),
            .lcout(\Lab_UT.didp.di_Mtens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21650),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_1_2_LC_7_4_5  (
            .in0(_gnd_net_),
            .in1(N__14124),
            .in2(_gnd_net_),
            .in3(N__17205),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_4_6 .LUT_INIT=16'b1100110001011010;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_2_LC_7_4_6  (
            .in0(N__15060),
            .in1(N__20765),
            .in2(N__14094),
            .in3(N__15188),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_2_LC_7_4_7 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_2_LC_7_4_7  (
            .in0(N__15051),
            .in1(N__15137),
            .in2(N__14091),
            .in3(N__15098),
            .lcout(\Lab_UT.didp.di_Mtens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21650),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_1_LC_7_5_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_1_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_1_LC_7_5_3 .LUT_INIT=16'b0001010100001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_1_LC_7_5_3  (
            .in0(N__21260),
            .in1(N__14598),
            .in2(N__17853),
            .in3(N__19647),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_5_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_5_4 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_2_ess_LC_7_5_4 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_LC_7_5_4  (
            .in0(N__19332),
            .in1(N__21100),
            .in2(N__14088),
            .in3(N__20924),
            .lcout(\Lab_UT.dictrl.state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21644),
            .ce(N__15872),
            .sr(N__19210));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI036C1_LC_7_5_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI036C1_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNI036C1_LC_7_5_5 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNI036C1_LC_7_5_5  (
            .in0(N__19418),
            .in1(N__18738),
            .in2(N__18477),
            .in3(N__19757),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_21_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIH9933_0_LC_7_5_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH9933_0_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIH9933_0_LC_7_5_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIH9933_0_LC_7_5_6  (
            .in0(_gnd_net_),
            .in1(N__20923),
            .in2(N__14586),
            .in3(N__14502),
            .lcout(\Lab_UT.i16_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIRKP91_LC_7_5_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIRKP91_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIRKP91_LC_7_5_7 .LUT_INIT=16'b0101010101000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNIRKP91_LC_7_5_7  (
            .in0(N__19417),
            .in1(N__19646),
            .in2(N__18258),
            .in3(N__14694),
            .lcout(\Lab_UT.dictrl.i18_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_7_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_1_1_LC_7_6_0 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_1_1_LC_7_6_0  (
            .in0(N__14458),
            .in1(N__17318),
            .in2(N__14364),
            .in3(N__15704),
            .lcout(\Lab_UT.dispString.dOut_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_7_6_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_7_6_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUC6L1_1_LC_7_6_1  (
            .in0(N__20930),
            .in1(N__19649),
            .in2(N__21259),
            .in3(N__19774),
            .lcout(\Lab_UT.LdMones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_7_6_2 .C_ON=1'b0;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dispString.dOut_RNO_2_3_LC_7_6_2 .LUT_INIT=16'b0010010100101111;
    LogicCell40 \Lab_UT.dispString.dOut_RNO_2_3_LC_7_6_2  (
            .in0(N__14457),
            .in1(N__17544),
            .in2(N__14363),
            .in3(N__17357),
            .lcout(\Lab_UT.dispString.m49_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_7_6_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_2_LC_7_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_2_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__18060),
            .in2(_gnd_net_),
            .in3(N__17950),
            .lcout(\Lab_UT.didp.countrce1.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_6_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_6_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_1_3_LC_7_6_5  (
            .in0(N__18061),
            .in1(N__16035),
            .in2(_gnd_net_),
            .in3(N__17951),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_6_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_6_6 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_3_LC_7_6_6  (
            .in0(N__17998),
            .in1(N__20491),
            .in2(N__14241),
            .in3(N__15993),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_6_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_3_LC_7_6_7 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_3_LC_7_6_7  (
            .in0(N__15806),
            .in1(N__15994),
            .in2(N__14238),
            .in3(N__15842),
            .lcout(\Lab_UT.didp.di_Sones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21636),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_7_7_0 .C_ON=1'b0;
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_idle_1_0_iclk_LC_7_7_0 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \Lab_UT.un1_idle_1_0_iclk_LC_7_7_0  (
            .in0(N__15582),
            .in1(N__17761),
            .in2(_gnd_net_),
            .in3(N__17819),
            .lcout(\Lab_UT.un1_idle_1_0_iclkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_7_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_7_7_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNI6H8A1_LC_7_7_2  (
            .in0(N__21217),
            .in1(N__19648),
            .in2(N__17628),
            .in3(N__19743),
            .lcout(\Lab_UT.LdMtens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.dicAlarmTrig_LC_7_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.dicAlarmTrig_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.dicAlarmTrig_LC_7_7_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.dicAlarmTrig_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__17762),
            .in2(_gnd_net_),
            .in3(N__17820),
            .lcout(G_186),
            .ltout(G_186_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_4_LC_7_7_5 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_4_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_4_LC_7_7_5 .LUT_INIT=16'b0000111100001101;
    LogicCell40 \Lab_UT.alarmchar_latch_4_LC_7_7_5  (
            .in0(N__17763),
            .in1(N__19282),
            .in2(N__14619),
            .in3(N__14616),
            .lcout(G_191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_10_LC_7_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_10_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_10_LC_7_7_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_10_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__20167),
            .in2(_gnd_net_),
            .in3(N__20608),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_2_ess_RNOZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_4_LC_7_7_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_4_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_4_LC_7_7_7 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_4_LC_7_7_7  (
            .in0(N__19744),
            .in1(N__19650),
            .in2(N__14601),
            .in3(N__20386),
            .lcout(\Lab_UT.dictrl.G_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNIRFD0E_LC_7_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNIRFD0E_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNIRFD0E_LC_7_8_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNIRFD0E_LC_7_8_0  (
            .in0(N__17901),
            .in1(N__16106),
            .in2(N__18175),
            .in3(N__16073),
            .lcout(),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_8_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_3_LC_7_8_1 .LUT_INIT=16'b0011011100000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_3_LC_7_8_1  (
            .in0(N__15918),
            .in1(N__19009),
            .in2(N__14589),
            .in3(N__14693),
            .lcout(\Lab_UT.dicRun_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21620),
            .ce(),
            .sr(N__19203));
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_3 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_ctle_3_LC_7_8_3  (
            .in0(N__19286),
            .in1(N__20886),
            .in2(N__21237),
            .in3(N__14691),
            .lcout(\Lab_UT.didp.regrce4.LdAMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_0_LC_7_8_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_0_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_0_LC_7_8_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.ce_0_LC_7_8_4  (
            .in0(N__14692),
            .in1(N__17634),
            .in2(N__15024),
            .in3(N__21204),
            .lcout(\Lab_UT.didp.ceZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21620),
            .ce(),
            .sr(N__19203));
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_7_8_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI51AM_0_LC_7_8_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI51AM_0_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(N__14673),
            .in2(_gnd_net_),
            .in3(N__15927),
            .lcout(\Lab_UT.didp.un1_dicLdSones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_1_LC_7_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_1_LC_7_8_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_1_LC_7_8_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.ce_1_LC_7_8_6  (
            .in0(N__15020),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15941),
            .lcout(\Lab_UT.didp.ceZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21620),
            .ce(),
            .sr(N__19203));
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_7_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI5U3I_1_LC_7_8_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.didp.ce_RNI5U3I_1_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__14667),
            .in2(_gnd_net_),
            .in3(N__14748),
            .lcout(\Lab_UT.didp.un1_dicLdStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_9_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_7_rep1_LC_7_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_LC_7_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14654),
            .lcout(bu_rx_data_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21614),
            .ce(N__19318),
            .sr(N__19234));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_LC_7_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_LC_7_10_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_LC_7_10_1  (
            .in0(N__18720),
            .in1(_gnd_net_),
            .in2(N__16376),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.dictrl.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_0_LC_7_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_0_LC_7_10_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIBOOF_0_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__16359),
            .in2(_gnd_net_),
            .in3(N__18719),
            .lcout(\Lab_UT.dictrl.N_189 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_10_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_LC_7_10_3  (
            .in0(N__20883),
            .in1(N__14800),
            .in2(N__14783),
            .in3(N__21098),
            .lcout(\Lab_UT.dictrl.state_1_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(N__15871),
            .sr(N__19207));
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_10_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_10_4 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_1_LC_7_10_4  (
            .in0(N__14802),
            .in1(N__21021),
            .in2(N__14782),
            .in3(N__20885),
            .lcout(\Lab_UT.dictrl.state_fast_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(N__15871),
            .sr(N__19207));
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_1_LC_7_10_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_1_LC_7_10_5  (
            .in0(N__20884),
            .in1(N__14801),
            .in2(N__14784),
            .in3(N__21099),
            .lcout(\Lab_UT.dictrl.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(N__15871),
            .sr(N__19207));
    defparam \Lab_UT.dictrl.state_ret_11_RNITTE7F_LC_7_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNITTE7F_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNITTE7F_LC_7_10_6 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNITTE7F_LC_7_10_6  (
            .in0(N__14799),
            .in1(N__21020),
            .in2(N__14781),
            .in3(N__20882),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_1 ),
            .ltout(\Lab_UT.dictrl.next_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_7_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_7_10_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_7_ess_LC_7_10_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \Lab_UT.dictrl.state_ret_7_ess_LC_7_10_7  (
            .in0(N__18302),
            .in1(N__21097),
            .in2(N__14751),
            .in3(N__16179),
            .lcout(\Lab_UT.LdStens_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21608),
            .ce(N__15871),
            .sr(N__19207));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_12_LC_7_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_12_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_12_LC_7_11_0 .LUT_INIT=16'b0100000001001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_12_LC_7_11_0  (
            .in0(N__16271),
            .in1(N__14853),
            .in2(N__14738),
            .in3(N__16159),
            .lcout(\Lab_UT.dictrl.N_81_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_10_LC_7_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_10_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_10_LC_7_11_3 .LUT_INIT=16'b0001111000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_10_LC_7_11_3  (
            .in0(N__16272),
            .in1(N__16283),
            .in2(N__14739),
            .in3(N__14837),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_95_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_6_LC_7_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_6_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_6_LC_7_11_4 .LUT_INIT=16'b1010111010111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_6_LC_7_11_4  (
            .in0(N__21048),
            .in1(N__20906),
            .in2(N__14712),
            .in3(N__14859),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_3_LC_7_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_3_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_3_LC_7_11_5 .LUT_INIT=16'b1111000111111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_3_LC_7_11_5  (
            .in0(N__20907),
            .in1(N__16301),
            .in2(N__14709),
            .in3(N__16386),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_0_LC_7_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_0_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_0_LC_7_11_6 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_0_LC_7_11_6  (
            .in0(N__14700),
            .in1(N__18198),
            .in2(N__14706),
            .in3(N__14910),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_ret_11and_0_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_LC_7_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_LC_7_11_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_11_LC_7_11_7 .LUT_INIT=16'b0000000001000110;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_LC_7_11_7  (
            .in0(N__18999),
            .in1(N__21049),
            .in2(N__14703),
            .in3(N__15583),
            .lcout(\Lab_UT.dictrl.un1_next_state66_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21602),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_2_LC_7_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_2_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_2_LC_7_12_0 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_2_LC_7_12_0  (
            .in0(N__18684),
            .in1(N__21022),
            .in2(N__21255),
            .in3(N__19802),
            .lcout(\Lab_UT.dictrl.g2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_2_5_LC_7_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_2_5_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_2_5_LC_7_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.g0_2_5_LC_7_12_1  (
            .in0(N__16469),
            .in1(N__16434),
            .in2(N__14901),
            .in3(N__16781),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_2Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIQOJQ3_LC_7_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIQOJQ3_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIQOJQ3_LC_7_12_2 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIQOJQ3_LC_7_12_2  (
            .in0(N__16378),
            .in1(N__16560),
            .in2(N__14880),
            .in3(N__18944),
            .lcout(\Lab_UT.dictrl.g2_0 ),
            .ltout(\Lab_UT.dictrl.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_9_LC_7_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_9_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_9_LC_7_12_3 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_9_LC_7_12_3  (
            .in0(N__19395),
            .in1(N__14868),
            .in2(N__14862),
            .in3(N__18747),
            .lcout(\Lab_UT.dictrl.N_90_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_15_LC_7_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_15_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_15_LC_7_12_4 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_15_LC_7_12_4  (
            .in0(N__18945),
            .in1(N__18786),
            .in2(N__16746),
            .in3(N__18375),
            .lcout(\Lab_UT.dictrl.m40_N_5_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g2_1_LC_7_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g2_1_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g2_1_LC_7_12_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \Lab_UT.dictrl.g2_1_LC_7_12_6  (
            .in0(N__16780),
            .in1(N__14900),
            .in2(_gnd_net_),
            .in3(N__18943),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI416J3_LC_7_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI416J3_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_RNI416J3_LC_7_12_7 .LUT_INIT=16'b0011000100111011;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_RNI416J3_LC_7_12_7  (
            .in0(N__18787),
            .in1(N__16270),
            .in2(N__14847),
            .in3(N__16379),
            .lcout(\Lab_UT.dictrl.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIVJEO_LC_7_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIVJEO_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNIVJEO_LC_7_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNIVJEO_LC_7_13_0  (
            .in0(N__19376),
            .in1(N__20375),
            .in2(N__21091),
            .in3(N__18382),
            .lcout(\Lab_UT.dictrl.g0_17_a6_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIE4AI_LC_7_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIE4AI_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIE4AI_LC_7_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIE4AI_LC_7_13_2  (
            .in0(N__14826),
            .in1(N__16377),
            .in2(N__21092),
            .in3(N__18383),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFEKI3_LC_7_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFEKI3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFEKI3_LC_7_13_3 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNIFEKI3_LC_7_13_3  (
            .in0(N__14820),
            .in1(N__14811),
            .in2(N__14805),
            .in3(N__18441),
            .lcout(\Lab_UT.dictrl.g0_17_0 ),
            .ltout(\Lab_UT.dictrl.g0_17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_1_LC_7_13_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_1_LC_7_13_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_1_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14913),
            .in3(N__16060),
            .lcout(\Lab_UT.dictrl.g2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_13_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep1_esr_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__18310),
            .in2(_gnd_net_),
            .in3(N__21057),
            .lcout(\Lab_UT.dictrl.state_3_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21593),
            .ce(N__15873),
            .sr(N__19212));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_13_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_13_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_LC_7_13_6  (
            .in0(N__21056),
            .in1(_gnd_net_),
            .in2(N__18315),
            .in3(_gnd_net_),
            .lcout(Lab_UT_dictrl_state_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21593),
            .ce(N__15873),
            .sr(N__19212));
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_13_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_13_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_3_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__18314),
            .in2(_gnd_net_),
            .in3(N__21058),
            .lcout(\Lab_UT.dictrl.state_fast_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21593),
            .ce(N__15873),
            .sr(N__19212));
    defparam \buart.Z_rx.shifter_4_LC_7_14_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_LC_7_14_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_LC_7_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20577),
            .lcout(bu_rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21592),
            .ce(N__19313),
            .sr(N__19238));
    defparam \buart.Z_rx.shifter_3_rep1_LC_7_14_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep1_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep1_LC_7_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep1_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20012),
            .lcout(bu_rx_data_3_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21592),
            .ce(N__19313),
            .sr(N__19238));
    defparam \buart.Z_rx.shifter_fast_4_LC_7_14_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_4_LC_7_14_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_4_LC_7_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_4_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20578),
            .lcout(bu_rx_data_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21592),
            .ce(N__19313),
            .sr(N__19238));
    defparam \buart.Z_rx.shifter_fast_3_LC_7_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_3_LC_7_14_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_3_LC_7_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_3_LC_7_14_6  (
            .in0(N__20013),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21592),
            .ce(N__19313),
            .sr(N__19238));
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_8_1_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNIDJKH1_3_LC_8_1_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNIDJKH1_3_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__14924),
            .in2(_gnd_net_),
            .in3(N__15197),
            .lcout(\Lab_UT.didp.un1_dicLdMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.ce_3_LC_8_2_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_3_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_3_LC_8_2_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.ce_3_LC_8_2_1  (
            .in0(N__15018),
            .in1(N__15959),
            .in2(N__15227),
            .in3(N__16652),
            .lcout(\Lab_UT.didp.ceZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_2_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_2_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIE21V3_3_LC_8_2_2  (
            .in0(N__15955),
            .in1(N__16651),
            .in2(N__15226),
            .in3(N__15014),
            .lcout(),
            .ltout(\Lab_UT.didp.ce_12_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.reset_3_LC_8_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_3_LC_8_2_3 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_3_LC_8_2_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.didp.reset_3_LC_8_2_3  (
            .in0(N__15069),
            .in1(N__15063),
            .in2(N__15027),
            .in3(N__15477),
            .lcout(\Lab_UT.didp.resetZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.ce_2_LC_8_2_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_2_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.ce_2_LC_8_2_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.ce_2_LC_8_2_4  (
            .in0(N__15956),
            .in1(N__15219),
            .in2(_gnd_net_),
            .in3(N__15016),
            .lcout(\Lab_UT.didp.ceZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.reset_1_LC_8_2_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_1_LC_8_2_5 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_1_LC_8_2_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.reset_1_LC_8_2_5  (
            .in0(N__15017),
            .in1(N__15218),
            .in2(_gnd_net_),
            .in3(N__15958),
            .lcout(\Lab_UT.didp.resetZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.reset_0_LC_8_2_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_0_LC_8_2_6 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_0_LC_8_2_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.reset_0_LC_8_2_6  (
            .in0(N__15957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15015),
            .lcout(\Lab_UT.didp.resetZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.reset_2_LC_8_2_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.reset_2_LC_8_2_7 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.didp.reset_2_LC_8_2_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.reset_2_LC_8_2_7  (
            .in0(N__15019),
            .in1(N__15960),
            .in2(N__15228),
            .in3(N__16653),
            .lcout(\Lab_UT.didp.resetZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21670),
            .ce(),
            .sr(N__19214));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_8_3_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_3_LC_8_3_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_3_LC_8_3_0  (
            .in0(N__15430),
            .in1(N__15631),
            .in2(_gnd_net_),
            .in3(N__15380),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce2.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_8_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_3_LC_8_3_1 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_3_LC_8_3_1  (
            .in0(N__15901),
            .in1(N__15341),
            .in2(N__14937),
            .in3(N__20507),
            .lcout(\Lab_UT.didp.countrce2.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_0_LC_8_3_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_0_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_0_LC_8_3_3 .LUT_INIT=16'b0010001000100001;
    LogicCell40 \Lab_UT.didp.countrce4.q_0_LC_8_3_3  (
            .in0(N__14934),
            .in1(N__15118),
            .in2(N__14928),
            .in3(N__15198),
            .lcout(\Lab_UT.didp.di_Mtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21663),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_3_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_3_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNI6SFG_3_LC_8_3_4  (
            .in0(N__15432),
            .in1(N__15340),
            .in2(N__15387),
            .in3(N__15632),
            .lcout(\Lab_UT.didp.un24_ce_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_8_3_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_1_LC_8_3_5 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_1_LC_8_3_5  (
            .in0(N__15381),
            .in1(N__20298),
            .in2(N__15903),
            .in3(N__15433),
            .lcout(\Lab_UT.didp.countrce2.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_3_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_3_7 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_0_LC_8_3_7  (
            .in0(N__15897),
            .in1(N__15431),
            .in2(_gnd_net_),
            .in3(N__19928),
            .lcout(\Lab_UT.didp.countrce2.q_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_8_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce4.q_RNO_0_3_LC_8_4_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Lab_UT.didp.countrce4.q_RNO_0_3_LC_8_4_0  (
            .in0(N__20499),
            .in1(N__15189),
            .in2(N__15153),
            .in3(N__15468),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce4.q_5_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce4.q_3_LC_8_4_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce4.q_3_LC_8_4_1  (
            .in0(N__15469),
            .in1(N__15136),
            .in2(N__15105),
            .in3(N__15102),
            .lcout(\Lab_UT.didp.di_Mtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21657),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_1_LC_8_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_1_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_1_LC_8_4_2 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \Lab_UT.didp.countrce2.q_1_LC_8_4_2  (
            .in0(N__15379),
            .in1(N__15282),
            .in2(N__15260),
            .in3(N__15078),
            .lcout(\Lab_UT.didp.di_Stens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21657),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_4_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_4_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_3_LC_8_4_3  (
            .in0(N__16898),
            .in1(N__17039),
            .in2(_gnd_net_),
            .in3(N__16992),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un20_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_4_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_3_LC_8_4_4  (
            .in0(N__20498),
            .in1(N__16942),
            .in2(N__15072),
            .in3(N__17076),
            .lcout(\Lab_UT.didp.countrce3.q_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_1_2_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__15413),
            .in2(_gnd_net_),
            .in3(N__15378),
            .lcout(\Lab_UT.didp.countrce2.un13_qPone ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5AJE1_3_LC_8_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5AJE1_3_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNI5AJE1_3_LC_8_4_6 .LUT_INIT=16'b1001000000001001;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNI5AJE1_3_LC_8_4_6  (
            .in0(N__17337),
            .in1(N__17075),
            .in2(N__16627),
            .in3(N__15467),
            .lcout(\Lab_UT.didp.did_alarmMatch_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_4_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_3_LC_8_4_7 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \Lab_UT.didp.countrce2.q_3_LC_8_4_7  (
            .in0(N__15450),
            .in1(N__15252),
            .in2(N__15288),
            .in3(N__15342),
            .lcout(\Lab_UT.didp.di_Stens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21657),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_0_LC_8_5_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.didp.countrce2.q_0_LC_8_5_0  (
            .in0(N__15286),
            .in1(N__15444),
            .in2(N__15434),
            .in3(N__15259),
            .lcout(\Lab_UT.didp.di_Stens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21651),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_8_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_8_5_2 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNIKRUF1_1_LC_8_5_2  (
            .in0(N__16879),
            .in1(N__17452),
            .in2(N__16996),
            .in3(N__17421),
            .lcout(\Lab_UT.didp.regrce3.did_alarmMatch_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_5_3 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.didp.regrce2.q_RNIG7M61_1_LC_8_5_3  (
            .in0(N__15385),
            .in1(N__15617),
            .in2(N__16815),
            .in3(N__17560),
            .lcout(\Lab_UT.didp.did_alarmMatch_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNITLJB1_3_LC_8_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITLJB1_3_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNITLJB1_3_LC_8_5_4 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNITLJB1_3_LC_8_5_4  (
            .in0(N__17535),
            .in1(N__15986),
            .in2(N__17263),
            .in3(N__15338),
            .lcout(),
            .ltout(\Lab_UT.didp.did_alarmMatch_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce3.q_RNI08DN5_1_LC_8_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_RNI08DN5_1_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce3.q_RNI08DN5_1_LC_8_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_RNI08DN5_1_LC_8_5_5  (
            .in0(N__15312),
            .in1(N__15306),
            .in2(N__15300),
            .in3(N__15297),
            .lcout(\Lab_UT.did_alarmMatch_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce2.q_2_LC_8_5_7 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \Lab_UT.didp.countrce2.q_2_LC_8_5_7  (
            .in0(N__15594),
            .in1(N__15287),
            .in2(N__15261),
            .in3(N__15618),
            .lcout(\Lab_UT.didp.di_Stens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21651),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_8_6_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_8_6_0 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_1_i_LC_8_6_0  (
            .in0(N__17825),
            .in1(N__19288),
            .in2(_gnd_net_),
            .in3(N__17756),
            .lcout(G_184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_RNIUNGG1_1_LC_8_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIUNGG1_1_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_RNIUNGG1_1_LC_8_6_1 .LUT_INIT=16'b1000001001000001;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_RNIUNGG1_1_LC_8_6_1  (
            .in0(N__17284),
            .in1(N__17308),
            .in2(N__17956),
            .in3(N__16030),
            .lcout(),
            .ltout(\Lab_UT.didp.did_alarmMatch_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIO6DH5_0_LC_8_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIO6DH5_0_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIO6DH5_0_LC_8_6_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIO6DH5_0_LC_8_6_2  (
            .in0(N__17142),
            .in1(N__15690),
            .in2(N__15678),
            .in3(N__15675),
            .lcout(\Lab_UT.did_alarmMatch_13 ),
            .ltout(\Lab_UT.did_alarmMatch_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_8_6_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_LC_8_6_3 .LUT_INIT=16'b0010101010101010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_0__m3_LC_8_6_3  (
            .in0(N__17700),
            .in1(N__17824),
            .in2(N__15669),
            .in3(N__15653),
            .lcout(),
            .ltout(\Lab_UT.dictrl.alarmstate_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_8_6_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_0_LC_8_6_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_0_LC_8_6_4  (
            .in0(N__15512),
            .in1(N__17826),
            .in2(N__15666),
            .in3(N__15493),
            .lcout(G_183),
            .ltout(G_183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_8_6_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_8_6_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_sqmuxa_LC_8_6_5  (
            .in0(N__17757),
            .in1(N__15663),
            .in2(N__15657),
            .in3(N__15654),
            .lcout(\Lab_UT.dictrl.alarmstate_1_sqmuxaZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_8_6_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce2.q_RNO_0_2_LC_8_6_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce2.q_RNO_0_2_LC_8_6_7  (
            .in0(N__20739),
            .in1(N__15642),
            .in2(N__15902),
            .in3(N__15627),
            .lcout(\Lab_UT.didp.countrce2.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_armed_4_LC_8_7_0 .C_ON=1'b0;
    defparam \Lab_UT.un1_armed_4_LC_8_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_armed_4_LC_8_7_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \Lab_UT.un1_armed_4_LC_8_7_0  (
            .in0(N__17813),
            .in1(N__15578),
            .in2(_gnd_net_),
            .in3(N__17736),
            .lcout(\Lab_UT.alarmstate_0_sqmuxa_1 ),
            .ltout(\Lab_UT.alarmstate_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_8_7_1 .C_ON=1'b0;
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_idle_5_0_iclk_LC_8_7_1 .LUT_INIT=16'b1111000111110001;
    LogicCell40 \Lab_UT.un1_idle_5_0_iclk_LC_8_7_1  (
            .in0(N__17738),
            .in1(N__17815),
            .in2(N__15516),
            .in3(_gnd_net_),
            .lcout(\Lab_UT.un1_idle_5_0_iclkZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_8_7_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_latch_1_LC_8_7_2 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_latch_1_LC_8_7_2  (
            .in0(N__17755),
            .in1(N__15513),
            .in2(N__15501),
            .in3(N__17640),
            .lcout(G_185),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_7_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_7_3 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_2_LC_8_7_3  (
            .in0(N__15852),
            .in1(N__20740),
            .in2(N__18002),
            .in3(N__16043),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce1.q_5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_7_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_2_LC_8_7_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \Lab_UT.didp.countrce1.q_2_LC_8_7_4  (
            .in0(N__15801),
            .in1(N__16039),
            .in2(N__15846),
            .in3(N__15832),
            .lcout(\Lab_UT.didp.di_Sones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21637),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_7_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce1.q_1_LC_8_7_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \Lab_UT.didp.countrce1.q_1_LC_8_7_5  (
            .in0(N__15831),
            .in1(N__17910),
            .in2(N__17960),
            .in3(N__15802),
            .lcout(\Lab_UT.didp.di_Sones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21637),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_8_7_6 .C_ON=1'b0;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.un1_armed_2_0_iso_i_LC_8_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \Lab_UT.un1_armed_2_0_iso_i_LC_8_7_6  (
            .in0(N__17814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17737),
            .lcout(\Lab_UT.un1_armed_2_0_iso_iZ0 ),
            .ltout(\Lab_UT.un1_armed_2_0_iso_iZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.alarmchar_latch_1_LC_8_7_7 .C_ON=1'b0;
    defparam \Lab_UT.alarmchar_latch_1_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.alarmchar_latch_1_LC_8_7_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \Lab_UT.alarmchar_latch_1_LC_8_7_7  (
            .in0(N__15765),
            .in1(N__15751),
            .in2(N__15708),
            .in3(N__15705),
            .lcout(G_192),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_0 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_0 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_LC_8_8_0  (
            .in0(N__21103),
            .in1(N__18186),
            .in2(_gnd_net_),
            .in3(N__17859),
            .lcout(\Lab_UT.dictrl.state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(N__15869),
            .sr(N__19205));
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_8_8_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_8_8_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_RNO_0_LC_8_8_1  (
            .in0(N__19527),
            .in1(N__17877),
            .in2(_gnd_net_),
            .in3(N__19756),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_113_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_8_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_8_8_2 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_5_ess_LC_8_8_2 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \Lab_UT.dictrl.state_ret_5_ess_LC_8_8_2  (
            .in0(N__16305),
            .in1(N__21101),
            .in2(N__15693),
            .in3(N__20893),
            .lcout(\Lab_UT.state_i_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(N__15869),
            .sr(N__19205));
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_2_LC_8_8_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_2_LC_8_8_3  (
            .in0(N__17896),
            .in1(N__16115),
            .in2(N__18177),
            .in3(N__16082),
            .lcout(\Lab_UT.dictrl.stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(N__15869),
            .sr(N__19205));
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_8_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_2_LC_8_8_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_2_LC_8_8_4  (
            .in0(N__16083),
            .in1(N__18174),
            .in2(N__16119),
            .in3(N__17897),
            .lcout(\Lab_UT.dictrl.state_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(N__15869),
            .sr(N__19205));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_8_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_LC_8_8_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_LC_8_8_5  (
            .in0(N__17895),
            .in1(N__16114),
            .in2(N__18176),
            .in3(N__16081),
            .lcout(\Lab_UT.dictrl.state_2_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21627),
            .ce(N__15869),
            .sr(N__19205));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIAD6S_LC_8_8_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIAD6S_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNIAD6S_LC_8_8_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNIAD6S_LC_8_8_6  (
            .in0(N__21197),
            .in1(N__18253),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(\Lab_UT.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_8_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_8_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNI28771_3_LC_8_8_7  (
            .in0(N__16034),
            .in1(N__17949),
            .in2(N__18068),
            .in3(N__15998),
            .lcout(\Lab_UT.didp.un18_ce ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_8_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_8_9_1 .SEQ_MODE=4'b1001;
    defparam \Lab_UT.dictrl.state_ret_8_ess_LC_8_9_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_8_ess_LC_8_9_1  (
            .in0(N__16177),
            .in1(N__18297),
            .in2(_gnd_net_),
            .in3(N__21083),
            .lcout(\Lab_UT.LdSones_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21621),
            .ce(N__15870),
            .sr(N__19208));
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_8_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_4_esr_LC_8_9_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_4_esr_LC_8_9_2  (
            .in0(N__21079),
            .in1(N__18287),
            .in2(_gnd_net_),
            .in3(N__16176),
            .lcout(\Lab_UT.LdSones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21621),
            .ce(N__15870),
            .sr(N__19208));
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_0_LC_8_9_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_0_LC_8_9_4  (
            .in0(N__16188),
            .in1(N__18542),
            .in2(N__21102),
            .in3(N__20887),
            .lcout(\Lab_UT.state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21621),
            .ce(N__15870),
            .sr(N__19208));
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_8_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_ret_6_esr_LC_8_9_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_ret_6_esr_LC_8_9_5  (
            .in0(N__16178),
            .in1(N__15917),
            .in2(N__18298),
            .in3(N__21084),
            .lcout(\Lab_UT.LdStens ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21621),
            .ce(N__15870),
            .sr(N__19208));
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_3_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__21078),
            .in2(_gnd_net_),
            .in3(N__18286),
            .lcout(\Lab_UT.state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21621),
            .ce(N__15870),
            .sr(N__19208));
    defparam \Lab_UT.dictrl.m25_0_LC_8_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m25_0_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m25_0_LC_8_10_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \Lab_UT.dictrl.m25_0_LC_8_10_0  (
            .in0(N__16534),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18912),
            .lcout(\Lab_UT.dictrl.m25Z0Z_0 ),
            .ltout(\Lab_UT.dictrl.m25Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m30_LC_8_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m30_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m30_LC_8_10_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.m30_LC_8_10_1  (
            .in0(N__16407),
            .in1(N__16227),
            .in2(N__16206),
            .in3(N__20380),
            .lcout(\Lab_UT.dictrl.N_114_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m59_ns_1_x1_LC_8_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m59_ns_1_x1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m59_ns_1_x1_LC_8_10_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \Lab_UT.dictrl.m59_ns_1_x1_LC_8_10_2  (
            .in0(N__16533),
            .in1(N__18911),
            .in2(N__18605),
            .in3(N__16406),
            .lcout(\Lab_UT.dictrl.m59_ns_1_xZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNILO8G6_LC_8_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNILO8G6_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNILO8G6_LC_8_10_3 .LUT_INIT=16'b0011010100000101;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_RNILO8G6_LC_8_10_3  (
            .in0(N__16160),
            .in1(N__19420),
            .in2(N__18750),
            .in3(N__17586),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_81_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIB544A_2_LC_8_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIB544A_2_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIB544A_2_LC_8_10_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIB544A_2_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__19520),
            .in2(N__16191),
            .in3(N__19794),
            .lcout(\Lab_UT.dictrl.N_113_1 ),
            .ltout(\Lab_UT.dictrl.N_113_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNIC32CN_LC_8_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNIC32CN_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNIC32CN_LC_8_10_5 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNIC32CN_LC_8_10_5  (
            .in0(N__20881),
            .in1(N__21023),
            .in2(N__16182),
            .in3(N__18543),
            .lcout(\Lab_UT.dictrl.next_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITSVD3_LC_8_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITSVD3_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNITSVD3_LC_8_10_6 .LUT_INIT=16'b0001000110101010;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNITSVD3_LC_8_10_6  (
            .in0(N__19421),
            .in1(N__18104),
            .in2(_gnd_net_),
            .in3(N__19793),
            .lcout(\Lab_UT.dictrl.i10_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNII0R67_1_LC_8_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNII0R67_1_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNII0R67_1_LC_8_10_7 .LUT_INIT=16'b0010000001110101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNII0R67_1_LC_8_10_7  (
            .in0(N__19645),
            .in1(N__21196),
            .in2(N__18108),
            .in3(N__16161),
            .lcout(\Lab_UT.dictrl.N_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m40_m2_0_LC_8_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m40_m2_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m40_m2_0_LC_8_11_0 .LUT_INIT=16'b1101110111010101;
    LogicCell40 \Lab_UT.dictrl.m40_m2_0_LC_8_11_0  (
            .in0(N__18789),
            .in1(N__21324),
            .in2(N__20254),
            .in3(N__18846),
            .lcout(\Lab_UT.dictrl.m40_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m73_1_LC_8_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m73_1_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m73_1_LC_8_11_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.m73_1_LC_8_11_1  (
            .in0(N__21325),
            .in1(N__20753),
            .in2(_gnd_net_),
            .in3(N__19912),
            .lcout(\Lab_UT.dictrl.m73Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_11_LC_8_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_11_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_11_LC_8_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_11_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__19407),
            .in2(_gnd_net_),
            .in3(N__18749),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_16_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_7_LC_8_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_7_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_7_LC_8_11_3 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_7_LC_8_11_3  (
            .in0(N__19795),
            .in1(N__16395),
            .in2(N__16389),
            .in3(N__16662),
            .lcout(\Lab_UT.dictrl.N_113_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_23_LC_8_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_23_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_23_LC_8_11_4 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \Lab_UT.dictrl.g0_23_LC_8_11_4  (
            .in0(N__16233),
            .in1(N__18850),
            .in2(N__16751),
            .in3(N__18354),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m40_N_5_mux_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI1N6L5_LC_8_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI1N6L5_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_2_rep1_esr_RNI1N6L5_LC_8_11_5 .LUT_INIT=16'b1001111100000110;
    LogicCell40 \Lab_UT.dictrl.state_0_2_rep1_esr_RNI1N6L5_LC_8_11_5  (
            .in0(N__18748),
            .in1(N__16366),
            .in2(N__16317),
            .in3(N__16551),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI5EFJC_LC_8_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI5EFJC_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI5EFJC_LC_8_11_6 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNI5EFJC_LC_8_11_6  (
            .in0(N__16314),
            .in1(N__16542),
            .in2(N__16308),
            .in3(N__19408),
            .lcout(\Lab_UT.dictrl.i9_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_12_LC_8_11_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_12_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_12_LC_8_11_7 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \Lab_UT.dictrl.g0_12_LC_8_11_7  (
            .in0(N__18353),
            .in1(N__18788),
            .in2(N__18866),
            .in3(N__16745),
            .lcout(\Lab_UT.dictrl.N_77_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_16_LC_8_12_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_16_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_16_LC_8_12_0 .LUT_INIT=16'b0000101100101111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_16_LC_8_12_0  (
            .in0(N__16260),
            .in1(N__18851),
            .in2(N__16752),
            .in3(N__18355),
            .lcout(\Lab_UT.dictrl.g2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_0_1_LC_8_12_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_0_1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_0_1_LC_8_12_1 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Lab_UT.dictrl.g0_0_1_LC_8_12_1  (
            .in0(N__16433),
            .in1(N__16531),
            .in2(N__16485),
            .in3(N__18901),
            .lcout(\Lab_UT.dictrl.g0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_2_4_LC_8_12_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_2_4_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_2_4_LC_8_12_2 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \Lab_UT.dictrl.g0_2_4_LC_8_12_2  (
            .in0(N__18900),
            .in1(_gnd_net_),
            .in2(N__16536),
            .in3(N__18419),
            .lcout(\Lab_UT.dictrl.g0_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_4_2_LC_8_12_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_4_2_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_4_2_LC_8_12_3 .LUT_INIT=16'b0000000000010101;
    LogicCell40 \Lab_UT.dictrl.g0_4_2_LC_8_12_3  (
            .in0(N__16484),
            .in1(N__18940),
            .in2(N__16785),
            .in3(N__16532),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_4Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_22_LC_8_12_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_22_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_22_LC_8_12_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.g0_22_LC_8_12_4  (
            .in0(N__19498),
            .in1(N__16750),
            .in2(N__16554),
            .in3(N__20573),
            .lcout(\Lab_UT.dictrl.N_77_1_0 ),
            .ltout(\Lab_UT.dictrl.N_77_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI11N26_LC_8_12_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI11N26_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_3_rep2_esr_RNI11N26_LC_8_12_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \Lab_UT.dictrl.state_0_3_rep2_esr_RNI11N26_LC_8_12_5  (
            .in0(N__19396),
            .in1(N__16680),
            .in2(N__16545),
            .in3(N__18515),
            .lcout(\Lab_UT.dictrl.N_2353_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m37_LC_8_12_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m37_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m37_LC_8_12_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.dictrl.m37_LC_8_12_6  (
            .in0(N__18899),
            .in1(N__16479),
            .in2(N__16535),
            .in3(N__16432),
            .lcout(\Lab_UT.dictrl.N_103_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTDF1_3_LC_8_12_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTDF1_3_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_fast_esr_RNIQTDF1_3_LC_8_12_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \Lab_UT.dictrl.state_0_fast_esr_RNIQTDF1_3_LC_8_12_7  (
            .in0(N__16480),
            .in1(N__16455),
            .in2(N__18910),
            .in3(N__16779),
            .lcout(\Lab_UT.dictrl.g1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m47_x0_LC_8_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m47_x0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m47_x0_LC_8_13_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \Lab_UT.dictrl.m47_x0_LC_8_13_0  (
            .in0(N__16423),
            .in1(N__20157),
            .in2(N__18628),
            .in3(N__20570),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m47_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m47_ns_LC_8_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m47_ns_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m47_ns_LC_8_13_1 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \Lab_UT.dictrl.m47_ns_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16437),
            .in3(N__16778),
            .lcout(\Lab_UT.dictrl.N_106_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m30_1_LC_8_13_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m30_1_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m30_1_LC_8_13_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.dictrl.m30_1_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(N__16422),
            .in2(_gnd_net_),
            .in3(N__16777),
            .lcout(\Lab_UT.dictrl.m30Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_fast_1_LC_8_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_1_LC_8_13_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_1_LC_8_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_1_LC_8_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20754),
            .lcout(bu_rx_data_fast_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__19314),
            .sr(N__19239));
    defparam \buart.Z_rx.shifter_5_LC_8_13_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_5_LC_8_13_5 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_5_LC_8_13_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_5_LC_8_13_5  (
            .in0(N__20158),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21596),
            .ce(N__19314),
            .sr(N__19239));
    defparam \Lab_UT.dictrl.g1_1_1_LC_8_14_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g1_1_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g1_1_1_LC_8_14_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \Lab_UT.dictrl.g1_1_1_LC_8_14_1  (
            .in0(N__16720),
            .in1(N__18423),
            .in2(_gnd_net_),
            .in3(N__18874),
            .lcout(\Lab_UT.dictrl.g1_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_13_LC_8_14_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_13_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_13_LC_8_14_5 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_13_LC_8_14_5  (
            .in0(N__20003),
            .in1(N__16671),
            .in2(_gnd_net_),
            .in3(N__18570),
            .lcout(\Lab_UT.dictrl.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_2_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_2_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNIAGOP1_3_LC_9_2_3  (
            .in0(N__17049),
            .in1(N__17002),
            .in2(N__16905),
            .in3(N__17087),
            .lcout(\Lab_UT.didp.countrce3.ce_12_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_9_3_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_0_LC_9_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_0_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19956),
            .lcout(\Lab_UT.di_AMtens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21671),
            .ce(N__16605),
            .sr(N__19215));
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_9_3_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_9_3_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce4.q_esr_3_LC_9_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_3_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20508),
            .lcout(\Lab_UT.di_AMtens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21671),
            .ce(N__16605),
            .sr(N__19215));
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_9_4_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.ce_RNI4EIS1_2_LC_9_4_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \Lab_UT.didp.ce_RNI4EIS1_2_LC_9_4_0  (
            .in0(_gnd_net_),
            .in1(N__17231),
            .in2(_gnd_net_),
            .in3(N__16955),
            .lcout(\Lab_UT.didp.un1_dicLdMones_0 ),
            .ltout(\Lab_UT.didp.un1_dicLdMones_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_4_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_1_LC_9_4_1 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \Lab_UT.didp.countrce3.q_1_LC_9_4_1  (
            .in0(N__16991),
            .in1(N__17127),
            .in2(N__16575),
            .in3(N__16572),
            .lcout(\Lab_UT.didp.di_Mones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21664),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_4_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_0_LC_9_4_2 .LUT_INIT=16'b0000110000001001;
    LogicCell40 \Lab_UT.didp.countrce3.q_0_LC_9_4_2  (
            .in0(N__17232),
            .in1(N__17217),
            .in2(N__17130),
            .in3(N__16956),
            .lcout(\Lab_UT.didp.di_Mones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21664),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_4_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_2_LC_9_4_3 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_2_LC_9_4_3  (
            .in0(N__16900),
            .in1(N__17128),
            .in2(N__16857),
            .in3(N__17096),
            .lcout(\Lab_UT.didp.di_Mones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21664),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_9_4_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_9_4_4 .LUT_INIT=16'b1000010000100001;
    LogicCell40 \Lab_UT.didp.regrce4.q_esr_RNIPTIE1_0_LC_9_4_4  (
            .in0(N__17027),
            .in1(N__17197),
            .in2(N__17503),
            .in3(N__17158),
            .lcout(\Lab_UT.didp.regrce4.did_alarmMatch_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.countrce3.q_3_LC_9_4_5 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \Lab_UT.didp.countrce3.q_3_LC_9_4_5  (
            .in0(N__17083),
            .in1(N__17129),
            .in2(N__17106),
            .in3(N__17097),
            .lcout(\Lab_UT.didp.di_Mones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21664),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_4_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_4_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_1_2_LC_9_4_6  (
            .in0(N__17028),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16990),
            .lcout(),
            .ltout(\Lab_UT.didp.countrce3.un13_qPone_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_4_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_4_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_4_7 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \Lab_UT.didp.countrce3.q_RNO_0_2_LC_9_4_7  (
            .in0(N__16954),
            .in1(N__20741),
            .in2(N__16908),
            .in3(N__16899),
            .lcout(\Lab_UT.didp.countrce3.q_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce2.q_0_LC_9_5_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_0_LC_9_5_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.didp.regrce2.q_0_LC_9_5_0  (
            .in0(N__20925),
            .in1(N__16842),
            .in2(N__17400),
            .in3(N__19950),
            .lcout(\Lab_UT.di_AStens_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce2.q_1_LC_9_5_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_1_LC_9_5_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_1_LC_9_5_1  (
            .in0(N__20296),
            .in1(N__20926),
            .in2(N__16822),
            .in3(N__17387),
            .lcout(\Lab_UT.di_AStens_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce2.q_2_LC_9_5_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_2_LC_9_5_2 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce2.q_2_LC_9_5_2  (
            .in0(N__20927),
            .in1(N__20742),
            .in2(N__17401),
            .in3(N__17566),
            .lcout(\Lab_UT.di_AStens_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce2.q_3_LC_9_5_3 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce2.q_3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce2.q_3_LC_9_5_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce2.q_3_LC_9_5_3  (
            .in0(N__20496),
            .in1(N__20928),
            .in2(N__17542),
            .in3(N__17391),
            .lcout(\Lab_UT.di_AStens_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce3.q_0_LC_9_5_4 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_0_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_0_LC_9_5_4 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \Lab_UT.didp.regrce3.q_0_LC_9_5_4  (
            .in0(N__17630),
            .in1(N__17493),
            .in2(N__17402),
            .in3(N__19951),
            .lcout(\Lab_UT.di_AMones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce3.q_1_LC_9_5_5 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_1_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_1_LC_9_5_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_1_LC_9_5_5  (
            .in0(N__20297),
            .in1(N__17631),
            .in2(N__17464),
            .in3(N__17395),
            .lcout(\Lab_UT.di_AMones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce3.q_2_LC_9_5_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_2_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_2_LC_9_5_6 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \Lab_UT.didp.regrce3.q_2_LC_9_5_6  (
            .in0(N__17632),
            .in1(N__20743),
            .in2(N__17403),
            .in3(N__17428),
            .lcout(\Lab_UT.di_AMones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce3.q_3_LC_9_5_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce3.q_3_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce3.q_3_LC_9_5_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \Lab_UT.didp.regrce3.q_3_LC_9_5_7  (
            .in0(N__20497),
            .in1(N__17633),
            .in2(N__17353),
            .in3(N__17399),
            .lcout(\Lab_UT.di_AMones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21658),
            .ce(),
            .sr(N__19213));
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_9_6_0 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_1_LC_9_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_1_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20295),
            .lcout(\Lab_UT.di_ASones_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21652),
            .ce(N__18662),
            .sr(N__19211));
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_6_1 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_2_LC_9_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_2_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20731),
            .lcout(\Lab_UT.di_ASones_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21652),
            .ce(N__18662),
            .sr(N__19211));
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_9_6_2 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \Lab_UT.didp.regrce1.q_esr_3_LC_9_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_3_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20492),
            .lcout(\Lab_UT.di_ASones_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21652),
            .ce(N__18662),
            .sr(N__19211));
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_9_7_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_3_LC_9_7_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_3_LC_9_7_0  (
            .in0(N__19499),
            .in1(N__20168),
            .in2(N__20609),
            .in3(N__19905),
            .lcout(\Lab_UT.dictrl.alarmstate8Z0Z_3 ),
            .ltout(\Lab_UT.dictrl.alarmstate8Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_0_LC_9_7_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_0_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate_1_0__m3_0_LC_9_7_1 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \Lab_UT.dictrl.alarmstate_1_0__m3_0_LC_9_7_1  (
            .in0(N__17827),
            .in1(N__17767),
            .in2(N__17703),
            .in3(N__18077),
            .lcout(\Lab_UT.dictrl.m3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.justentered_1_sqmuxa_i_LC_9_7_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.justentered_1_sqmuxa_i_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.justentered_1_sqmuxa_i_LC_9_7_3 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \Lab_UT.dictrl.justentered_1_sqmuxa_i_LC_9_7_3  (
            .in0(N__17651),
            .in1(N__17676),
            .in2(N__17670),
            .in3(N__19289),
            .lcout(),
            .ltout(\Lab_UT.dictrl.justentered_1_sqmuxa_iZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.justentered_latch_LC_9_7_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.justentered_latch_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.justentered_latch_LC_9_7_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \Lab_UT.dictrl.justentered_latch_LC_9_7_4  (
            .in0(N__17691),
            .in1(_gnd_net_),
            .in2(N__17694),
            .in3(N__17652),
            .lcout(G_188),
            .ltout(G_188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate22_LC_9_7_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate22_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate22_LC_9_7_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \Lab_UT.dictrl.alarmstate22_LC_9_7_5  (
            .in0(N__17685),
            .in1(_gnd_net_),
            .in2(N__17679),
            .in3(N__18078),
            .lcout(G_187),
            .ltout(G_187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_9_7_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_9_7_6 .LUT_INIT=16'b1111111100001100;
    LogicCell40 \Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_i_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__17669),
            .in2(N__17655),
            .in3(N__17650),
            .lcout(\Lab_UT.dictrl.un1_alarmstate_1_sqmuxa_1_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIA8O21_LC_9_8_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIA8O21_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNIA8O21_LC_9_8_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNIA8O21_LC_9_8_0  (
            .in0(N__21251),
            .in1(N__18493),
            .in2(N__17629),
            .in3(N__19739),
            .lcout(\Lab_UT.LdASones ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_2_2_LC_9_8_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_2_2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_2_2_LC_9_8_2 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \Lab_UT.dictrl.g0_2_2_LC_9_8_2  (
            .in0(N__19503),
            .in1(N__20156),
            .in2(N__18632),
            .in3(N__20602),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_2Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_15_LC_9_8_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_15_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_15_LC_9_8_3 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \Lab_UT.dictrl.g0_15_LC_9_8_3  (
            .in0(N__18854),
            .in1(N__18379),
            .in2(N__17589),
            .in3(N__21333),
            .lcout(\Lab_UT.dictrl.m40_N_5_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.alarmstate8_4_LC_9_8_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.alarmstate8_4_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.alarmstate8_4_LC_9_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \Lab_UT.dictrl.alarmstate8_4_LC_9_8_5  (
            .in0(N__18853),
            .in1(N__20379),
            .in2(N__18384),
            .in3(N__21332),
            .lcout(\Lab_UT.dictrl.alarmstate8Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_6 .C_ON=1'b0;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \Lab_UT.didp.countrce1.q_RNO_0_1_LC_9_8_6  (
            .in0(N__20285),
            .in1(N__18069),
            .in2(N__17994),
            .in3(N__17952),
            .lcout(\Lab_UT.didp.countrce1.q_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_2_LC_9_9_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_LC_9_9_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_LC_9_9_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_2_LC_9_9_0  (
            .in0(N__20428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21628),
            .ce(N__19319),
            .sr(N__19236));
    defparam \Lab_UT.dictrl.g0_17_o3_2_LC_9_9_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_o3_2_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_o3_2_LC_9_9_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \Lab_UT.dictrl.g0_17_o3_2_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__20427),
            .in2(_gnd_net_),
            .in3(N__20671),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIS3A93_1_LC_9_9_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIS3A93_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIS3A93_1_LC_9_9_2 .LUT_INIT=16'b0111111101110101;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIS3A93_1_LC_9_9_2  (
            .in0(N__20879),
            .in1(N__18798),
            .in2(N__17904),
            .in3(N__19676),
            .lcout(\Lab_UT.dictrl.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_9_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_9_9_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_5_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__20426),
            .in2(_gnd_net_),
            .in3(N__20670),
            .lcout(\Lab_UT.dictrl.m51_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_9_9_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_9_9_6 .LUT_INIT=16'b0001101110111011;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_0_LC_9_9_6  (
            .in0(N__20880),
            .in1(N__18450),
            .in2(N__17876),
            .in3(N__19755),
            .lcout(\Lab_UT.dictrl.next_state_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_LC_9_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_LC_9_9_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_LC_9_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_3_LC_9_9_7  (
            .in0(N__20057),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21628),
            .ce(N__19319),
            .sr(N__19236));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_5_LC_9_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_5_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_5_LC_9_10_0 .LUT_INIT=16'b1000110101010101;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_5_LC_9_10_0  (
            .in0(N__19655),
            .in1(N__18264),
            .in2(N__18144),
            .in3(N__20038),
            .lcout(\Lab_UT.dictrl.P8_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIUI6O8_0_LC_9_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUI6O8_0_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIUI6O8_0_LC_9_10_1 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIUI6O8_0_LC_9_10_1  (
            .in0(N__20878),
            .in1(N__18219),
            .in2(N__18213),
            .in3(N__18135),
            .lcout(\Lab_UT.dictrl.next_state_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_12_LC_9_10_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_12_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_12_LC_9_10_2 .LUT_INIT=16'b0001000011110111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_12_LC_9_10_2  (
            .in0(N__20264),
            .in1(N__20698),
            .in2(N__19809),
            .in3(N__20472),
            .lcout(\Lab_UT.dictrl.P6_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI0C4D4_LC_9_10_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI0C4D4_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNI0C4D4_LC_9_10_3 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNI0C4D4_LC_9_10_3  (
            .in0(N__18257),
            .in1(N__19419),
            .in2(N__18231),
            .in3(N__19654),
            .lcout(\Lab_UT.dictrl.N_69 ),
            .ltout(\Lab_UT.dictrl.N_69_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_4_LC_9_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_4_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_4_LC_9_10_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_4_LC_9_10_4  (
            .in0(N__18134),
            .in1(N__18212),
            .in2(N__18201),
            .in3(N__20877),
            .lcout(\Lab_UT.dictrl.next_state_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_10_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_1_LC_9_10_5  (
            .in0(N__19781),
            .in1(N__18090),
            .in2(N__19677),
            .in3(N__20775),
            .lcout(\Lab_UT.dictrl.state_ret_1_ess_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNIIOLT_LC_9_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNIIOLT_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNIIOLT_LC_9_10_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNIIOLT_LC_9_10_6  (
            .in0(N__21096),
            .in1(N__21176),
            .in2(_gnd_net_),
            .in3(N__19780),
            .lcout(\Lab_UT.dictrl.g0_17_a6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_11_LC_9_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_11_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_11_LC_9_10_7 .LUT_INIT=16'b0101000101110101;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_11_LC_9_10_7  (
            .in0(N__20471),
            .in1(N__20697),
            .in2(N__21216),
            .in3(N__20263),
            .lcout(\Lab_UT.dictrl.P6_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNI00K56_3_LC_9_11_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNI00K56_3_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNI00K56_3_LC_9_11_0 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNI00K56_3_LC_9_11_0  (
            .in0(N__18133),
            .in1(N__18089),
            .in2(N__21238),
            .in3(N__18103),
            .lcout(\Lab_UT.dictrl.m77_ns_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m55_0_LC_9_11_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m55_0_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m55_0_LC_9_11_1 .LUT_INIT=16'b0000000001001100;
    LogicCell40 \Lab_UT.dictrl.m55_0_LC_9_11_1  (
            .in0(N__20250),
            .in1(N__18790),
            .in2(N__20764),
            .in3(N__21326),
            .lcout(\Lab_UT.dictrl.N_77 ),
            .ltout(\Lab_UT.dictrl.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIRLAN5_3_LC_9_11_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIRLAN5_3_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIRLAN5_3_LC_9_11_2 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIRLAN5_3_LC_9_11_2  (
            .in0(N__18522),
            .in1(N__21211),
            .in2(N__18564),
            .in3(N__18561),
            .lcout(),
            .ltout(\Lab_UT.dictrl.state_0_esr_RNIRLAN5Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_0_esr_RNIASHNC_1_LC_9_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_esr_RNIASHNC_1_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_esr_RNIASHNC_1_LC_9_11_3 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \Lab_UT.dictrl.state_0_esr_RNIASHNC_1_LC_9_11_3  (
            .in0(N__18552),
            .in1(N__19672),
            .in2(N__18546),
            .in3(N__19778),
            .lcout(\Lab_UT.dictrl.i9_mux_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_4_LC_9_11_4  (
            .in0(N__18521),
            .in1(N__18504),
            .in2(N__21239),
            .in3(N__19927),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_118_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_9_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_9_11_5 .LUT_INIT=16'b0101010111000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_2_LC_9_11_5  (
            .in0(N__21212),
            .in1(N__18495),
            .in2(N__18453),
            .in3(N__19779),
            .lcout(\Lab_UT.dictrl.next_state_latmux_3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.g0_17_a6_3_7_LC_9_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.g0_17_a6_3_7_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.g0_17_a6_3_7_LC_9_11_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \Lab_UT.dictrl.g0_17_a6_3_7_LC_9_11_6  (
            .in0(N__20155),
            .in1(N__20604),
            .in2(N__20052),
            .in3(N__19926),
            .lcout(\Lab_UT.dictrl.g0_17_a6_3Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_1_LC_9_12_0 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_LC_9_12_0 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_LC_9_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_LC_9_12_0  (
            .in0(N__20732),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_fast_0_LC_9_12_1 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_0_LC_9_12_1 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_0_LC_9_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_0_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20246),
            .lcout(buart__rx_shifter_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_12_2 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_12_2 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_1_rep1_LC_9_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_1_rep1_LC_9_12_2  (
            .in0(N__20733),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_1_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_12_3 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_2_rep1_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_2_rep1_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20488),
            .lcout(bu_rx_data_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_fast_2_LC_9_12_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_2_LC_9_12_4 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_2_LC_9_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_fast_2_LC_9_12_4  (
            .in0(N__20489),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_fast_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_3_rep2_LC_9_12_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_LC_9_12_6 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_3_rep2_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20048),
            .lcout(bu_rx_data_3_rep2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \buart.Z_rx.shifter_fast_5_LC_9_12_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_fast_5_LC_9_12_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_fast_5_LC_9_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_fast_5_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20160),
            .lcout(buart__rx_shifter_fast_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21609),
            .ce(N__19317),
            .sr(N__19240));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNID53P_LC_9_13_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNID53P_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_RNID53P_LC_9_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_RNID53P_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__19402),
            .in2(_gnd_net_),
            .in3(N__18751),
            .lcout(N_16_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_8_LC_9_13_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_8_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_8_LC_9_13_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_8_LC_9_13_1  (
            .in0(N__21328),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18852),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_11_RNO_5_LC_9_13_2 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_5_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_11_RNO_5_LC_9_13_2 .LUT_INIT=16'b0111111101110101;
    LogicCell40 \Lab_UT.dictrl.state_ret_11_RNO_5_LC_9_13_2  (
            .in0(N__20935),
            .in1(N__18791),
            .in2(N__18756),
            .in3(N__18752),
            .lcout(\Lab_UT.dictrl.N_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_3_rep2_RNIT8A31_LC_9_13_4 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_3_rep2_RNIT8A31_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_3_rep2_RNIT8A31_LC_9_13_4 .LUT_INIT=16'b0000010011011111;
    LogicCell40 \buart.Z_rx.shifter_3_rep2_RNIT8A31_LC_9_13_4  (
            .in0(N__20223),
            .in1(N__19403),
            .in2(N__20755),
            .in3(N__21327),
            .lcout(\buart.Z_rx.P7_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_13_7 .C_ON=1'b0;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_13_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \Lab_UT.didp.regrce1.q_esr_ctle_3_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__18672),
            .in2(_gnd_net_),
            .in3(N__19285),
            .lcout(\Lab_UT.didp.regrce1.LdASones_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_7_rep1_RNIG7Q01_LC_9_14_5 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_7_rep1_RNIG7Q01_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_7_rep1_RNIG7Q01_LC_9_14_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \buart.Z_rx.shifter_7_rep1_RNIG7Q01_LC_9_14_5  (
            .in0(N__18627),
            .in1(N__20159),
            .in2(_gnd_net_),
            .in3(N__20571),
            .lcout(shifter_7_rep1_RNIG7Q01),
            .ltout(shifter_7_rep1_RNIG7Q01_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_RNIUOH63_4_LC_9_14_6 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_RNIUOH63_4_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \buart.Z_rx.shifter_RNIUOH63_4_LC_9_14_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \buart.Z_rx.shifter_RNIUOH63_4_LC_9_14_6  (
            .in0(N__19545),
            .in1(N__19536),
            .in2(N__19530),
            .in3(N__20030),
            .lcout(N_97),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_4_rep1_LC_9_14_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_4_rep1_LC_9_14_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_4_rep1_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \buart.Z_rx.shifter_4_rep1_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20572),
            .lcout(bu_rx_data_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21597),
            .ce(N__19315),
            .sr(N__19241));
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_ctle_LC_11_8_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_ctle_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_0_1_rep1_esr_ctle_LC_11_8_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \Lab_UT.dictrl.state_0_1_rep1_esr_ctle_LC_11_8_4  (
            .in0(N__19017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19283),
            .lcout(bu_rx_data_rdy_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_9_LC_11_9_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_9_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_9_LC_11_9_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_9_LC_11_9_3  (
            .in0(N__19812),
            .in1(N__20169),
            .in2(N__19428),
            .in3(N__19873),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_5_a4_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_3_LC_11_9_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_3_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_3_LC_11_9_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_3_LC_11_9_4  (
            .in0(N__21276),
            .in1(N__20056),
            .in2(N__19338),
            .in3(N__20287),
            .lcout(),
            .ltout(\Lab_UT.dictrl.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_11_9_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_11_9_5 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_0_LC_11_9_5  (
            .in0(N__21236),
            .in1(N__19554),
            .in2(N__19335),
            .in3(N__19671),
            .lcout(\Lab_UT.dictrl.N_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buart.Z_rx.shifter_0_LC_11_9_7 .C_ON=1'b0;
    defparam \buart.Z_rx.shifter_0_LC_11_9_7 .SEQ_MODE=4'b1010;
    defparam \buart.Z_rx.shifter_0_LC_11_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \buart.Z_rx.shifter_0_LC_11_9_7  (
            .in0(N__20288),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(bu_rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21639),
            .ce(N__19320),
            .sr(N__19237));
    defparam \Lab_UT.dictrl.m86_LC_11_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m86_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m86_LC_11_10_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.m86_LC_11_10_0  (
            .in0(N__19010),
            .in1(N__21267),
            .in2(N__18960),
            .in3(N__20388),
            .lcout(N_119_mux),
            .ltout(N_119_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_0_LC_11_10_1 .C_ON=1'b0;
    defparam \resetGen.reset_count_0_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_0_LC_11_10_1 .LUT_INIT=16'b0000110000000011;
    LogicCell40 \resetGen.reset_count_0_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__21398),
            .in2(N__21360),
            .in3(N__21759),
            .lcout(resetGen_reset_count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21631),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_8_LC_11_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_8_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_8_LC_11_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_8_LC_11_10_4  (
            .in0(N__20610),
            .in1(N__20757),
            .in2(N__21357),
            .in3(N__20387),
            .lcout(\Lab_UT.dictrl.g0_5_a4_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m86_0_LC_11_10_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m86_0_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m86_0_LC_11_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \Lab_UT.dictrl.m86_0_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(N__20037),
            .in2(_gnd_net_),
            .in3(N__20284),
            .lcout(),
            .ltout(\Lab_UT.dictrl.m86Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m86_2_LC_11_10_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m86_2_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m86_2_LC_11_10_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \Lab_UT.dictrl.m86_2_LC_11_10_6  (
            .in0(N__20490),
            .in1(N__20756),
            .in2(N__21270),
            .in3(N__19872),
            .lcout(\Lab_UT.dictrl.m86Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_11_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_11_10_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_1_ess_RNO_3_LC_11_10_7  (
            .in0(N__21243),
            .in1(N__21105),
            .in2(_gnd_net_),
            .in3(N__20936),
            .lcout(\Lab_UT.dictrl.next_state_latmux_1_a0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_6_LC_11_11_3 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_6_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_6_LC_11_11_3 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_6_LC_11_11_3  (
            .in0(N__20752),
            .in1(N__20603),
            .in2(N__20506),
            .in3(N__20373),
            .lcout(\Lab_UT.dictrl.g0_5_o4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_7_LC_11_11_5 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_7_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_7_LC_11_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_7_LC_11_11_5  (
            .in0(N__20286),
            .in1(N__20162),
            .in2(N__20058),
            .in3(N__19888),
            .lcout(),
            .ltout(\Lab_UT.dictrl.g0_5_o4_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_2_LC_11_11_6 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_2_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.state_ret_2_ess_RNO_2_LC_11_11_6 .LUT_INIT=16'b0011001000000000;
    LogicCell40 \Lab_UT.dictrl.state_ret_2_ess_RNO_2_LC_11_11_6  (
            .in0(N__19821),
            .in1(N__19811),
            .in2(N__19680),
            .in3(N__19670),
            .lcout(\Lab_UT.dictrl.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m90_LC_12_10_0 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m90_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m90_LC_12_10_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \Lab_UT.dictrl.m90_LC_12_10_0  (
            .in0(N__21417),
            .in1(N__21755),
            .in2(N__21713),
            .in3(N__21729),
            .lcout(N_91_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m93_LC_12_10_1 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m93_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m93_LC_12_10_1 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \Lab_UT.dictrl.m93_LC_12_10_1  (
            .in0(N__21757),
            .in1(N__21419),
            .in2(N__21737),
            .in3(N__21711),
            .lcout(),
            .ltout(N_117_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_3_LC_12_10_2 .C_ON=1'b0;
    defparam \resetGen.reset_count_3_LC_12_10_2 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_3_LC_12_10_2 .LUT_INIT=16'b1011100110101000;
    LogicCell40 \resetGen.reset_count_3_LC_12_10_2  (
            .in0(N__21689),
            .in1(N__21366),
            .in2(N__21762),
            .in3(N__21680),
            .lcout(\resetGen.reset_countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21640),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_1_LC_12_10_3 .C_ON=1'b0;
    defparam \resetGen.reset_count_1_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_1_LC_12_10_3 .LUT_INIT=16'b0011000000010010;
    LogicCell40 \resetGen.reset_count_1_LC_12_10_3  (
            .in0(N__21758),
            .in1(N__21421),
            .in2(N__21738),
            .in3(N__21392),
            .lcout(resetGen_reset_count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21640),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m97_LC_12_10_4 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m97_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m97_LC_12_10_4 .LUT_INIT=16'b0001010001010000;
    LogicCell40 \Lab_UT.dictrl.m97_LC_12_10_4  (
            .in0(N__21418),
            .in1(N__21756),
            .in2(N__21714),
            .in3(N__21730),
            .lcout(),
            .ltout(resetGen_reset_count_2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_2_LC_12_10_5 .C_ON=1'b0;
    defparam \resetGen.reset_count_2_LC_12_10_5 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_2_LC_12_10_5 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \resetGen.reset_count_2_LC_12_10_5  (
            .in0(N__21396),
            .in1(N__21423),
            .in2(N__21717),
            .in3(N__21712),
            .lcout(resetGen_reset_count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21640),
            .ce(),
            .sr(_gnd_net_));
    defparam \resetGen.reset_count_4_LC_12_10_6 .C_ON=1'b0;
    defparam \resetGen.reset_count_4_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \resetGen.reset_count_4_LC_12_10_6 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \resetGen.reset_count_4_LC_12_10_6  (
            .in0(N__21422),
            .in1(N__21397),
            .in2(N__21693),
            .in3(N__21681),
            .lcout(resetGen_reset_count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21640),
            .ce(),
            .sr(_gnd_net_));
    defparam \Lab_UT.dictrl.m87_LC_12_10_7 .C_ON=1'b0;
    defparam \Lab_UT.dictrl.m87_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \Lab_UT.dictrl.m87_LC_12_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \Lab_UT.dictrl.m87_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(N__21420),
            .in2(_gnd_net_),
            .in3(N__21391),
            .lcout(m87),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // latticehx1k
